magic
tech sky130A
magscale 1 2
timestamp 1769196051
<< viali >>
rect 18889 35717 18923 35751
rect 19625 35717 19659 35751
rect 1409 35649 1443 35683
rect 1685 35649 1719 35683
rect 1961 35649 1995 35683
rect 11897 35649 11931 35683
rect 18521 35649 18555 35683
rect 25697 35649 25731 35683
rect 27905 35649 27939 35683
rect 34529 35649 34563 35683
rect 11989 35581 12023 35615
rect 12173 35581 12207 35615
rect 19717 35581 19751 35615
rect 19901 35581 19935 35615
rect 25513 35581 25547 35615
rect 25605 35581 25639 35615
rect 27997 35581 28031 35615
rect 28089 35581 28123 35615
rect 34345 35581 34379 35615
rect 1593 35513 1627 35547
rect 1869 35513 1903 35547
rect 20177 35513 20211 35547
rect 11529 35445 11563 35479
rect 12449 35445 12483 35479
rect 18705 35445 18739 35479
rect 18981 35445 19015 35479
rect 19257 35445 19291 35479
rect 26065 35445 26099 35479
rect 26249 35445 26283 35479
rect 27445 35445 27479 35479
rect 27537 35445 27571 35479
rect 1409 35241 1443 35275
rect 19073 35241 19107 35275
rect 25881 35241 25915 35275
rect 28733 35241 28767 35275
rect 14657 35105 14691 35139
rect 14933 35105 14967 35139
rect 7389 35037 7423 35071
rect 9505 35037 9539 35071
rect 11069 35037 11103 35071
rect 13829 35037 13863 35071
rect 14565 35037 14599 35071
rect 15117 35037 15151 35071
rect 17693 35037 17727 35071
rect 17960 35037 17994 35071
rect 19625 35037 19659 35071
rect 22201 35037 22235 35071
rect 24409 35037 24443 35071
rect 26994 35037 27028 35071
rect 27261 35037 27295 35071
rect 27353 35037 27387 35071
rect 27620 35037 27654 35071
rect 7656 34969 7690 35003
rect 9750 34969 9784 35003
rect 11336 34969 11370 35003
rect 15384 34969 15418 35003
rect 19892 34969 19926 35003
rect 22468 34969 22502 35003
rect 24676 34969 24710 35003
rect 8769 34901 8803 34935
rect 10885 34901 10919 34935
rect 12449 34901 12483 34935
rect 13645 34901 13679 34935
rect 14105 34901 14139 34935
rect 14473 34901 14507 34935
rect 16497 34901 16531 34935
rect 21005 34901 21039 34935
rect 23581 34901 23615 34935
rect 25789 34901 25823 34935
rect 8125 34697 8159 34731
rect 9045 34697 9079 34731
rect 9597 34697 9631 34731
rect 9965 34697 9999 34731
rect 14841 34697 14875 34731
rect 15577 34697 15611 34731
rect 16037 34697 16071 34731
rect 20177 34697 20211 34731
rect 20545 34697 20579 34731
rect 23305 34697 23339 34731
rect 23673 34697 23707 34731
rect 24593 34697 24627 34731
rect 24961 34697 24995 34731
rect 28181 34697 28215 34731
rect 8585 34629 8619 34663
rect 24409 34629 24443 34663
rect 8493 34561 8527 34595
rect 10057 34561 10091 34595
rect 10701 34561 10735 34595
rect 12256 34561 12290 34595
rect 13461 34561 13495 34595
rect 13728 34561 13762 34595
rect 15945 34561 15979 34595
rect 18337 34561 18371 34595
rect 20637 34561 20671 34595
rect 21833 34561 21867 34595
rect 22100 34561 22134 34595
rect 23765 34561 23799 34595
rect 28089 34561 28123 34595
rect 8677 34493 8711 34527
rect 10241 34493 10275 34527
rect 10425 34493 10459 34527
rect 11989 34493 12023 34527
rect 16221 34493 16255 34527
rect 16405 34493 16439 34527
rect 18429 34493 18463 34527
rect 18613 34493 18647 34527
rect 18797 34493 18831 34527
rect 19073 34493 19107 34527
rect 19809 34493 19843 34527
rect 20821 34493 20855 34527
rect 21005 34493 21039 34527
rect 23857 34493 23891 34527
rect 25053 34493 25087 34527
rect 25145 34493 25179 34527
rect 28273 34493 28307 34527
rect 11621 34425 11655 34459
rect 24133 34425 24167 34459
rect 13369 34357 13403 34391
rect 17969 34357 18003 34391
rect 23213 34357 23247 34391
rect 27721 34357 27755 34391
rect 13185 34153 13219 34187
rect 18797 34153 18831 34187
rect 22109 34153 22143 34187
rect 26525 34153 26559 34187
rect 28733 34153 28767 34187
rect 19073 34085 19107 34119
rect 26157 34085 26191 34119
rect 6285 34017 6319 34051
rect 11345 34017 11379 34051
rect 13737 34017 13771 34051
rect 14105 34017 14139 34051
rect 22569 34017 22603 34051
rect 22753 34017 22787 34051
rect 26341 34017 26375 34051
rect 26709 34017 26743 34051
rect 1409 33949 1443 33983
rect 1685 33949 1719 33983
rect 5365 33949 5399 33983
rect 5641 33949 5675 33983
rect 8953 33949 8987 33983
rect 10517 33949 10551 33983
rect 10610 33949 10644 33983
rect 10793 33949 10827 33983
rect 11023 33949 11057 33983
rect 13553 33949 13587 33983
rect 14381 33949 14415 33983
rect 14657 33949 14691 33983
rect 14749 33949 14783 33983
rect 15209 33949 15243 33983
rect 17417 33949 17451 33983
rect 17684 33949 17718 33983
rect 18889 33949 18923 33983
rect 22477 33949 22511 33983
rect 23213 33949 23247 33983
rect 23489 33949 23523 33983
rect 23581 33949 23615 33983
rect 25329 33949 25363 33983
rect 25513 33949 25547 33983
rect 25605 33949 25639 33983
rect 25697 33949 25731 33983
rect 25973 33949 26007 33983
rect 27353 33949 27387 33983
rect 27620 33949 27654 33983
rect 33241 33949 33275 33983
rect 34069 33949 34103 33983
rect 6552 33881 6586 33915
rect 7757 33881 7791 33915
rect 9220 33881 9254 33915
rect 10885 33881 10919 33915
rect 11529 33881 11563 33915
rect 14565 33881 14599 33915
rect 15025 33881 15059 33915
rect 15945 33881 15979 33915
rect 23397 33881 23431 33915
rect 34345 33881 34379 33915
rect 1593 33813 1627 33847
rect 7665 33813 7699 33847
rect 10333 33813 10367 33847
rect 11161 33813 11195 33847
rect 13645 33813 13679 33847
rect 14933 33813 14967 33847
rect 15761 33813 15795 33847
rect 16681 33813 16715 33847
rect 21281 33813 21315 33847
rect 23029 33813 23063 33847
rect 23765 33813 23799 33847
rect 23857 33813 23891 33847
rect 24133 33813 24167 33847
rect 25881 33813 25915 33847
rect 26985 33813 27019 33847
rect 32873 33813 32907 33847
rect 33057 33813 33091 33847
rect 7389 33609 7423 33643
rect 7757 33609 7791 33643
rect 8861 33609 8895 33643
rect 10241 33609 10275 33643
rect 10425 33609 10459 33643
rect 16497 33609 16531 33643
rect 19533 33609 19567 33643
rect 26985 33609 27019 33643
rect 34345 33609 34379 33643
rect 7113 33541 7147 33575
rect 9873 33541 9907 33575
rect 9965 33541 9999 33575
rect 15393 33541 15427 33575
rect 16129 33541 16163 33575
rect 16926 33541 16960 33575
rect 18521 33541 18555 33575
rect 18981 33541 19015 33575
rect 19073 33541 19107 33575
rect 20637 33541 20671 33575
rect 21833 33541 21867 33575
rect 26556 33541 26590 33575
rect 27445 33541 27479 33575
rect 28641 33541 28675 33575
rect 5080 33473 5114 33507
rect 6377 33473 6411 33507
rect 9229 33473 9263 33507
rect 9689 33473 9723 33507
rect 10057 33473 10091 33507
rect 11796 33473 11830 33507
rect 15025 33473 15059 33507
rect 15118 33473 15152 33507
rect 15301 33473 15335 33507
rect 15531 33473 15565 33507
rect 18705 33473 18739 33507
rect 18798 33473 18832 33507
rect 19211 33473 19245 33507
rect 20453 33473 20487 33507
rect 20729 33473 20763 33507
rect 20821 33473 20855 33507
rect 21097 33473 21131 33507
rect 21373 33473 21407 33507
rect 23029 33473 23063 33507
rect 27353 33473 27387 33507
rect 28273 33473 28307 33507
rect 28421 33473 28455 33507
rect 28549 33473 28583 33507
rect 28738 33473 28772 33507
rect 29285 33473 29319 33507
rect 29469 33473 29503 33507
rect 29561 33473 29595 33507
rect 29837 33473 29871 33507
rect 34161 33473 34195 33507
rect 34437 33473 34471 33507
rect 4813 33405 4847 33439
rect 7849 33405 7883 33439
rect 8033 33405 8067 33439
rect 9321 33405 9355 33439
rect 9505 33405 9539 33439
rect 11529 33405 11563 33439
rect 15945 33405 15979 33439
rect 16037 33405 16071 33439
rect 16681 33405 16715 33439
rect 21189 33405 21223 33439
rect 22293 33405 22327 33439
rect 26801 33405 26835 33439
rect 27629 33405 27663 33439
rect 29653 33405 29687 33439
rect 30113 33405 30147 33439
rect 32137 33405 32171 33439
rect 32413 33405 32447 33439
rect 10517 33337 10551 33371
rect 18061 33337 18095 33371
rect 19349 33337 19383 33371
rect 21005 33337 21039 33371
rect 21557 33337 21591 33371
rect 28917 33337 28951 33371
rect 30021 33337 30055 33371
rect 33977 33337 34011 33371
rect 6193 33269 6227 33303
rect 8309 33269 8343 33303
rect 12909 33269 12943 33303
rect 15669 33269 15703 33303
rect 21097 33269 21131 33303
rect 23121 33269 23155 33303
rect 25421 33269 25455 33303
rect 29101 33269 29135 33303
rect 33885 33269 33919 33303
rect 5457 33065 5491 33099
rect 10057 33065 10091 33099
rect 11713 33065 11747 33099
rect 17969 33065 18003 33099
rect 30941 33065 30975 33099
rect 32229 33065 32263 33099
rect 34529 33065 34563 33099
rect 8033 32997 8067 33031
rect 10425 32997 10459 33031
rect 23765 32997 23799 33031
rect 26893 32997 26927 33031
rect 27169 32997 27203 33031
rect 27445 32997 27479 33031
rect 6101 32929 6135 32963
rect 8125 32929 8159 32963
rect 9781 32929 9815 32963
rect 10149 32929 10183 32963
rect 12357 32929 12391 32963
rect 13369 32929 13403 32963
rect 14105 32929 14139 32963
rect 18061 32929 18095 32963
rect 32781 32929 32815 32963
rect 33057 32929 33091 32963
rect 6285 32861 6319 32895
rect 7389 32861 7423 32895
rect 7537 32861 7571 32895
rect 7895 32861 7929 32895
rect 10057 32861 10091 32895
rect 10517 32861 10551 32895
rect 12173 32861 12207 32895
rect 12725 32861 12759 32895
rect 12909 32861 12943 32895
rect 13001 32861 13035 32895
rect 13185 32861 13219 32895
rect 13277 32861 13311 32895
rect 15669 32861 15703 32895
rect 15853 32861 15887 32895
rect 16957 32861 16991 32895
rect 17233 32861 17267 32895
rect 17417 32861 17451 32895
rect 17509 32861 17543 32895
rect 17601 32861 17635 32895
rect 17785 32861 17819 32895
rect 19257 32861 19291 32895
rect 21097 32861 21131 32895
rect 23581 32861 23615 32895
rect 24409 32861 24443 32895
rect 25881 32861 25915 32895
rect 25974 32861 26008 32895
rect 26157 32861 26191 32895
rect 26387 32861 26421 32895
rect 29561 32861 29595 32895
rect 32413 32861 32447 32895
rect 32689 32861 32723 32895
rect 5825 32793 5859 32827
rect 7665 32793 7699 32827
rect 7757 32793 7791 32827
rect 8401 32793 8435 32827
rect 14372 32793 14406 32827
rect 16221 32793 16255 32827
rect 19524 32793 19558 32827
rect 21364 32793 21398 32827
rect 22569 32793 22603 32827
rect 24654 32793 24688 32827
rect 26249 32793 26283 32827
rect 26709 32793 26743 32827
rect 28825 32793 28859 32827
rect 29828 32793 29862 32827
rect 32597 32793 32631 32827
rect 5917 32725 5951 32759
rect 7021 32725 7055 32759
rect 12081 32725 12115 32759
rect 12633 32725 12667 32759
rect 13553 32725 13587 32759
rect 15485 32725 15519 32759
rect 18337 32725 18371 32759
rect 20637 32725 20671 32759
rect 22477 32725 22511 32759
rect 25789 32725 25823 32759
rect 26525 32725 26559 32759
rect 26985 32725 27019 32759
rect 28641 32725 28675 32759
rect 9137 32521 9171 32555
rect 9597 32521 9631 32555
rect 13737 32521 13771 32555
rect 14473 32521 14507 32555
rect 14841 32521 14875 32555
rect 19625 32521 19659 32555
rect 19993 32521 20027 32555
rect 21005 32521 21039 32555
rect 24777 32521 24811 32555
rect 27997 32521 28031 32555
rect 10149 32453 10183 32487
rect 11161 32453 11195 32487
rect 15393 32453 15427 32487
rect 20085 32453 20119 32487
rect 28825 32453 28859 32487
rect 29653 32453 29687 32487
rect 29837 32453 29871 32487
rect 3700 32385 3734 32419
rect 6377 32385 6411 32419
rect 7757 32385 7791 32419
rect 8024 32385 8058 32419
rect 12624 32385 12658 32419
rect 17049 32385 17083 32419
rect 21189 32385 21223 32419
rect 21281 32385 21315 32419
rect 21465 32385 21499 32419
rect 21557 32385 21591 32419
rect 22569 32385 22603 32419
rect 22836 32385 22870 32419
rect 24869 32385 24903 32419
rect 28181 32385 28215 32419
rect 28273 32385 28307 32419
rect 28365 32385 28399 32419
rect 28549 32385 28583 32419
rect 3433 32317 3467 32351
rect 9689 32317 9723 32351
rect 9873 32317 9907 32351
rect 10977 32317 11011 32351
rect 12357 32317 12391 32351
rect 14933 32317 14967 32351
rect 15117 32317 15151 32351
rect 17141 32317 17175 32351
rect 17325 32317 17359 32351
rect 19533 32317 19567 32351
rect 20177 32317 20211 32351
rect 21833 32317 21867 32351
rect 25053 32317 25087 32351
rect 28641 32317 28675 32351
rect 9229 32249 9263 32283
rect 24409 32249 24443 32283
rect 4813 32181 4847 32215
rect 6561 32181 6595 32215
rect 16681 32181 16715 32215
rect 17601 32181 17635 32215
rect 22109 32181 22143 32215
rect 23949 32181 23983 32215
rect 6653 31977 6687 32011
rect 7573 31977 7607 32011
rect 9597 31977 9631 32011
rect 9781 31977 9815 32011
rect 12817 31977 12851 32011
rect 16681 31977 16715 32011
rect 21465 31977 21499 32011
rect 23121 31977 23155 32011
rect 26065 31977 26099 32011
rect 26249 31977 26283 32011
rect 28089 31977 28123 32011
rect 29561 31977 29595 32011
rect 6745 31909 6779 31943
rect 11621 31909 11655 31943
rect 22385 31909 22419 31943
rect 28181 31909 28215 31943
rect 4353 31841 4387 31875
rect 7297 31841 7331 31875
rect 10149 31841 10183 31875
rect 12265 31841 12299 31875
rect 12541 31841 12575 31875
rect 13461 31841 13495 31875
rect 21925 31841 21959 31875
rect 22109 31841 22143 31875
rect 23673 31841 23707 31875
rect 28825 31841 28859 31875
rect 30021 31841 30055 31875
rect 30205 31841 30239 31875
rect 30941 31841 30975 31875
rect 32781 31841 32815 31875
rect 33057 31841 33091 31875
rect 1409 31773 1443 31807
rect 1685 31773 1719 31807
rect 4629 31773 4663 31807
rect 5273 31773 5307 31807
rect 5540 31773 5574 31807
rect 7205 31773 7239 31807
rect 7757 31773 7791 31807
rect 8125 31773 8159 31807
rect 8953 31773 8987 31807
rect 9101 31773 9135 31807
rect 9321 31773 9355 31807
rect 9418 31773 9452 31807
rect 10416 31773 10450 31807
rect 11989 31773 12023 31807
rect 13185 31773 13219 31807
rect 15301 31773 15335 31807
rect 17233 31773 17267 31807
rect 21833 31773 21867 31807
rect 22937 31773 22971 31807
rect 23581 31773 23615 31807
rect 25881 31773 25915 31807
rect 25973 31773 26007 31807
rect 26709 31773 26743 31807
rect 28549 31773 28583 31807
rect 29101 31773 29135 31807
rect 7113 31705 7147 31739
rect 7849 31705 7883 31739
rect 7941 31705 7975 31739
rect 9229 31705 9263 31739
rect 13277 31705 13311 31739
rect 15568 31705 15602 31739
rect 17500 31705 17534 31739
rect 26976 31705 27010 31739
rect 28641 31705 28675 31739
rect 29929 31705 29963 31739
rect 30757 31705 30791 31739
rect 2421 31637 2455 31671
rect 8309 31637 8343 31671
rect 11529 31637 11563 31671
rect 12081 31637 12115 31671
rect 13737 31637 13771 31671
rect 18613 31637 18647 31671
rect 23489 31637 23523 31671
rect 30389 31637 30423 31671
rect 30849 31637 30883 31671
rect 34529 31637 34563 31671
rect 1409 31433 1443 31467
rect 2605 31433 2639 31467
rect 5365 31433 5399 31467
rect 6377 31433 6411 31467
rect 9505 31433 9539 31467
rect 9597 31433 9631 31467
rect 10057 31433 10091 31467
rect 17417 31433 17451 31467
rect 17785 31433 17819 31467
rect 21097 31433 21131 31467
rect 21465 31433 21499 31467
rect 26065 31433 26099 31467
rect 26801 31433 26835 31467
rect 29469 31433 29503 31467
rect 31401 31433 31435 31467
rect 33977 31433 34011 31467
rect 8392 31365 8426 31399
rect 11805 31365 11839 31399
rect 11897 31365 11931 31399
rect 18245 31365 18279 31399
rect 20821 31365 20855 31399
rect 30288 31365 30322 31399
rect 34345 31365 34379 31399
rect 34805 31365 34839 31399
rect 3729 31297 3763 31331
rect 3985 31297 4019 31331
rect 4077 31297 4111 31331
rect 4353 31297 4387 31331
rect 7490 31297 7524 31331
rect 7757 31297 7791 31331
rect 8125 31297 8159 31331
rect 9965 31297 9999 31331
rect 10885 31297 10919 31331
rect 11069 31297 11103 31331
rect 11161 31297 11195 31331
rect 11708 31297 11742 31331
rect 12080 31297 12114 31331
rect 12173 31297 12207 31331
rect 16681 31297 16715 31331
rect 16865 31297 16899 31331
rect 17233 31297 17267 31331
rect 18153 31297 18187 31331
rect 18613 31297 18647 31331
rect 18880 31297 18914 31331
rect 20545 31297 20579 31331
rect 20729 31297 20763 31331
rect 20913 31297 20947 31331
rect 23213 31297 23247 31331
rect 24860 31297 24894 31331
rect 26249 31297 26283 31331
rect 26341 31297 26375 31331
rect 26525 31297 26559 31331
rect 26617 31297 26651 31331
rect 28089 31297 28123 31331
rect 28356 31297 28390 31331
rect 30021 31297 30055 31331
rect 34161 31297 34195 31331
rect 34437 31297 34471 31331
rect 34529 31297 34563 31331
rect 5457 31229 5491 31263
rect 5641 31229 5675 31263
rect 10149 31229 10183 31263
rect 16957 31229 16991 31263
rect 17049 31229 17083 31263
rect 18337 31229 18371 31263
rect 21281 31229 21315 31263
rect 22937 31229 22971 31263
rect 23305 31229 23339 31263
rect 23581 31229 23615 31263
rect 24593 31229 24627 31263
rect 4997 31161 5031 31195
rect 11529 31161 11563 31195
rect 11161 31093 11195 31127
rect 11345 31093 11379 31127
rect 12357 31093 12391 31127
rect 12541 31093 12575 31127
rect 12725 31093 12759 31127
rect 17693 31093 17727 31127
rect 19993 31093 20027 31127
rect 23029 31093 23063 31127
rect 25973 31093 26007 31127
rect 26985 31093 27019 31127
rect 3985 30889 4019 30923
rect 6285 30889 6319 30923
rect 25145 30889 25179 30923
rect 28457 30889 28491 30923
rect 31769 30889 31803 30923
rect 5457 30821 5491 30855
rect 15945 30821 15979 30855
rect 18613 30821 18647 30855
rect 19257 30821 19291 30855
rect 25053 30821 25087 30855
rect 31401 30821 31435 30855
rect 31585 30821 31619 30855
rect 4629 30753 4663 30787
rect 6745 30753 6779 30787
rect 6837 30753 6871 30787
rect 19901 30753 19935 30787
rect 25697 30753 25731 30787
rect 28273 30753 28307 30787
rect 28917 30753 28951 30787
rect 29009 30753 29043 30787
rect 30757 30753 30791 30787
rect 4445 30685 4479 30719
rect 4813 30685 4847 30719
rect 4906 30685 4940 30719
rect 5181 30685 5215 30719
rect 5319 30685 5353 30719
rect 6653 30685 6687 30719
rect 12265 30685 12299 30719
rect 13829 30685 13863 30719
rect 14105 30685 14139 30719
rect 15577 30685 15611 30719
rect 19625 30685 19659 30719
rect 20453 30685 20487 30719
rect 22293 30685 22327 30719
rect 24409 30685 24443 30719
rect 24502 30685 24536 30719
rect 24777 30685 24811 30719
rect 24874 30685 24908 30719
rect 25513 30685 25547 30719
rect 28825 30685 28859 30719
rect 30389 30685 30423 30719
rect 30573 30685 30607 30719
rect 30665 30685 30699 30719
rect 30941 30685 30975 30719
rect 31217 30685 31251 30719
rect 31953 30685 31987 30719
rect 34069 30685 34103 30719
rect 4353 30617 4387 30651
rect 5089 30617 5123 30651
rect 12532 30617 12566 30651
rect 14372 30617 14406 30651
rect 20698 30617 20732 30651
rect 22560 30617 22594 30651
rect 24685 30617 24719 30651
rect 25605 30617 25639 30651
rect 26157 30617 26191 30651
rect 31125 30617 31159 30651
rect 34345 30617 34379 30651
rect 5641 30549 5675 30583
rect 7205 30549 7239 30583
rect 13645 30549 13679 30583
rect 15485 30549 15519 30583
rect 15761 30549 15795 30583
rect 17601 30549 17635 30583
rect 19717 30549 19751 30583
rect 20177 30549 20211 30583
rect 21833 30549 21867 30583
rect 23673 30549 23707 30583
rect 25973 30549 26007 30583
rect 4813 30345 4847 30379
rect 5181 30345 5215 30379
rect 12817 30345 12851 30379
rect 14565 30345 14599 30379
rect 15025 30345 15059 30379
rect 19349 30345 19383 30379
rect 20821 30345 20855 30379
rect 21281 30345 21315 30379
rect 22845 30345 22879 30379
rect 23213 30345 23247 30379
rect 27905 30345 27939 30379
rect 9321 30277 9355 30311
rect 10517 30277 10551 30311
rect 11069 30277 11103 30311
rect 13185 30277 13219 30311
rect 13277 30277 13311 30311
rect 13921 30277 13955 30311
rect 14013 30277 14047 30311
rect 14933 30277 14967 30311
rect 18337 30277 18371 30311
rect 21189 30277 21223 30311
rect 28273 30277 28307 30311
rect 28457 30277 28491 30311
rect 33977 30277 34011 30311
rect 1409 30209 1443 30243
rect 1685 30209 1719 30243
rect 4261 30209 4295 30243
rect 4445 30209 4479 30243
rect 4537 30209 4571 30243
rect 4629 30209 4663 30243
rect 9413 30209 9447 30243
rect 10333 30209 10367 30243
rect 10609 30209 10643 30243
rect 10701 30209 10735 30243
rect 11161 30209 11195 30243
rect 13829 30209 13863 30243
rect 14197 30209 14231 30243
rect 15485 30209 15519 30243
rect 15578 30209 15612 30243
rect 15761 30209 15795 30243
rect 15853 30209 15887 30243
rect 15991 30209 16025 30243
rect 18061 30209 18095 30243
rect 18245 30209 18279 30243
rect 18429 30209 18463 30243
rect 18889 30209 18923 30243
rect 21925 30209 21959 30243
rect 26985 30209 27019 30243
rect 27078 30209 27112 30243
rect 27261 30209 27295 30243
rect 27353 30209 27387 30243
rect 27450 30209 27484 30243
rect 27721 30209 27755 30243
rect 28089 30209 28123 30243
rect 29285 30209 29319 30243
rect 33793 30209 33827 30243
rect 34069 30209 34103 30243
rect 9597 30141 9631 30175
rect 13369 30141 13403 30175
rect 15117 30141 15151 30175
rect 16313 30141 16347 30175
rect 19165 30141 19199 30175
rect 19257 30141 19291 30175
rect 21465 30141 21499 30175
rect 23305 30141 23339 30175
rect 23489 30141 23523 30175
rect 34161 30141 34195 30175
rect 34437 30141 34471 30175
rect 10885 30073 10919 30107
rect 13645 30073 13679 30107
rect 16129 30073 16163 30107
rect 18613 30073 18647 30107
rect 26709 30073 26743 30107
rect 27629 30073 27663 30107
rect 1593 30005 1627 30039
rect 4905 30005 4939 30039
rect 8953 30005 8987 30039
rect 9873 30005 9907 30039
rect 14473 30005 14507 30039
rect 16405 30005 16439 30039
rect 19717 30005 19751 30039
rect 23765 30005 23799 30039
rect 25053 30005 25087 30039
rect 29101 30005 29135 30039
rect 29377 30005 29411 30039
rect 29653 30005 29687 30039
rect 33425 30005 33459 30039
rect 33609 30005 33643 30039
rect 3617 29801 3651 29835
rect 8769 29801 8803 29835
rect 10977 29801 11011 29835
rect 14381 29801 14415 29835
rect 15025 29801 15059 29835
rect 18705 29801 18739 29835
rect 20637 29801 20671 29835
rect 21281 29801 21315 29835
rect 23673 29801 23707 29835
rect 25789 29801 25823 29835
rect 27445 29801 27479 29835
rect 29561 29801 29595 29835
rect 30573 29801 30607 29835
rect 34529 29801 34563 29835
rect 12725 29733 12759 29767
rect 29377 29733 29411 29767
rect 5273 29665 5307 29699
rect 9229 29665 9263 29699
rect 11345 29665 11379 29699
rect 13369 29665 13403 29699
rect 13645 29665 13679 29699
rect 15209 29665 15243 29699
rect 16957 29665 16991 29699
rect 21373 29665 21407 29699
rect 22569 29665 22603 29699
rect 24409 29665 24443 29699
rect 27997 29665 28031 29699
rect 33057 29665 33091 29699
rect 2237 29597 2271 29631
rect 3801 29597 3835 29631
rect 6745 29597 6779 29631
rect 8217 29597 8251 29631
rect 8401 29597 8435 29631
rect 8585 29597 8619 29631
rect 9045 29597 9079 29631
rect 9597 29597 9631 29631
rect 13185 29597 13219 29631
rect 13277 29597 13311 29631
rect 14657 29597 14691 29631
rect 14841 29597 14875 29631
rect 15393 29597 15427 29631
rect 19257 29597 19291 29631
rect 19524 29597 19558 29631
rect 20729 29597 20763 29631
rect 21005 29597 21039 29631
rect 21097 29597 21131 29631
rect 22477 29597 22511 29631
rect 23121 29597 23155 29631
rect 23489 29597 23523 29631
rect 26065 29597 26099 29631
rect 29745 29597 29779 29631
rect 30113 29597 30147 29631
rect 32781 29597 32815 29631
rect 2504 29529 2538 29563
rect 4068 29529 4102 29563
rect 5540 29529 5574 29563
rect 7012 29529 7046 29563
rect 8493 29529 8527 29563
rect 9864 29529 9898 29563
rect 11612 29529 11646 29563
rect 15660 29529 15694 29563
rect 17224 29529 17258 29563
rect 20913 29529 20947 29563
rect 23305 29529 23339 29563
rect 23397 29529 23431 29563
rect 24676 29529 24710 29563
rect 26332 29529 26366 29563
rect 28264 29529 28298 29563
rect 29837 29529 29871 29563
rect 29929 29529 29963 29563
rect 30389 29529 30423 29563
rect 5181 29461 5215 29495
rect 6653 29461 6687 29495
rect 8125 29461 8159 29495
rect 12817 29461 12851 29495
rect 16773 29461 16807 29495
rect 18337 29461 18371 29495
rect 22017 29461 22051 29495
rect 22385 29461 22419 29495
rect 30205 29461 30239 29495
rect 3065 29257 3099 29291
rect 3433 29257 3467 29291
rect 4261 29257 4295 29291
rect 4629 29257 4663 29291
rect 4721 29257 4755 29291
rect 6745 29257 6779 29291
rect 6837 29257 6871 29291
rect 7389 29257 7423 29291
rect 7757 29257 7791 29291
rect 9781 29257 9815 29291
rect 10149 29257 10183 29291
rect 10517 29257 10551 29291
rect 14473 29257 14507 29291
rect 14933 29257 14967 29291
rect 15761 29257 15795 29291
rect 16129 29257 16163 29291
rect 17417 29257 17451 29291
rect 17785 29257 17819 29291
rect 23213 29257 23247 29291
rect 24685 29257 24719 29291
rect 25053 29257 25087 29291
rect 25145 29257 25179 29291
rect 26985 29257 27019 29291
rect 27445 29257 27479 29291
rect 28549 29257 28583 29291
rect 28917 29257 28951 29291
rect 30849 29257 30883 29291
rect 3525 29189 3559 29223
rect 5273 29189 5307 29223
rect 7849 29189 7883 29223
rect 13268 29189 13302 29223
rect 16221 29189 16255 29223
rect 18245 29189 18279 29223
rect 22100 29189 22134 29223
rect 23765 29189 23799 29223
rect 8401 29121 8435 29155
rect 8668 29121 8702 29155
rect 10609 29121 10643 29155
rect 14841 29121 14875 29155
rect 19717 29121 19751 29155
rect 19984 29121 20018 29155
rect 21833 29121 21867 29155
rect 23673 29121 23707 29155
rect 27353 29121 27387 29155
rect 29009 29121 29043 29155
rect 29469 29121 29503 29155
rect 29736 29121 29770 29155
rect 3709 29053 3743 29087
rect 4905 29053 4939 29087
rect 6009 29053 6043 29087
rect 6929 29053 6963 29087
rect 8033 29053 8067 29087
rect 10701 29053 10735 29087
rect 10977 29053 11011 29087
rect 13001 29053 13035 29087
rect 15025 29053 15059 29087
rect 15301 29053 15335 29087
rect 16313 29053 16347 29087
rect 16681 29053 16715 29087
rect 17877 29053 17911 29087
rect 18061 29053 18095 29087
rect 23857 29053 23891 29087
rect 24593 29053 24627 29087
rect 25329 29053 25363 29087
rect 27537 29053 27571 29087
rect 27813 29053 27847 29087
rect 29101 29053 29135 29087
rect 3985 28985 4019 29019
rect 6377 28985 6411 29019
rect 8309 28985 8343 29019
rect 14381 28985 14415 29019
rect 21097 28985 21131 29019
rect 23305 28917 23339 28951
rect 6377 28713 6411 28747
rect 20269 28713 20303 28747
rect 24133 28713 24167 28747
rect 29745 28713 29779 28747
rect 6469 28645 6503 28679
rect 20729 28577 20763 28611
rect 20821 28577 20855 28611
rect 27169 28577 27203 28611
rect 30297 28577 30331 28611
rect 5549 28509 5583 28543
rect 14381 28509 14415 28543
rect 14657 28509 14691 28543
rect 17417 28509 17451 28543
rect 20637 28509 20671 28543
rect 22753 28509 22787 28543
rect 23020 28509 23054 28543
rect 30113 28509 30147 28543
rect 27436 28441 27470 28475
rect 29653 28441 29687 28475
rect 30205 28441 30239 28475
rect 3433 28373 3467 28407
rect 17233 28373 17267 28407
rect 28549 28373 28583 28407
rect 29377 28373 29411 28407
rect 1593 28169 1627 28203
rect 7941 28169 7975 28203
rect 14197 28169 14231 28203
rect 16037 28169 16071 28203
rect 23121 28169 23155 28203
rect 26801 28169 26835 28203
rect 27629 28169 27663 28203
rect 27997 28169 28031 28203
rect 3065 28101 3099 28135
rect 4537 28101 4571 28135
rect 4997 28101 5031 28135
rect 7389 28101 7423 28135
rect 14381 28101 14415 28135
rect 15669 28101 15703 28135
rect 15853 28101 15887 28135
rect 16313 28101 16347 28135
rect 22753 28101 22787 28135
rect 27169 28101 27203 28135
rect 27261 28101 27295 28135
rect 1409 28033 1443 28067
rect 1685 28033 1719 28067
rect 2789 28033 2823 28067
rect 3249 28033 3283 28067
rect 4169 28033 4203 28067
rect 4261 28033 4295 28067
rect 4445 28033 4479 28067
rect 4629 28033 4663 28067
rect 6009 28033 6043 28067
rect 6745 28033 6779 28067
rect 7205 28033 7239 28067
rect 7481 28033 7515 28067
rect 7573 28033 7607 28067
rect 12642 28033 12676 28067
rect 16681 28033 16715 28067
rect 16937 28033 16971 28067
rect 20085 28033 20119 28067
rect 21649 28033 21683 28067
rect 25320 28033 25354 28067
rect 26985 28033 27019 28067
rect 27353 28033 27387 28067
rect 34529 28033 34563 28067
rect 3893 27965 3927 27999
rect 6837 27965 6871 27999
rect 7021 27965 7055 27999
rect 8125 27965 8159 27999
rect 12909 27965 12943 27999
rect 15117 27965 15151 27999
rect 20177 27965 20211 27999
rect 20361 27965 20395 27999
rect 22017 27965 22051 27999
rect 25053 27965 25087 27999
rect 28089 27965 28123 27999
rect 28181 27965 28215 27999
rect 28457 27965 28491 27999
rect 34805 27965 34839 27999
rect 6193 27897 6227 27931
rect 7757 27897 7791 27931
rect 29377 27897 29411 27931
rect 4813 27829 4847 27863
rect 5181 27829 5215 27863
rect 6377 27829 6411 27863
rect 8861 27829 8895 27863
rect 11529 27829 11563 27863
rect 18061 27829 18095 27863
rect 18153 27829 18187 27863
rect 19717 27829 19751 27863
rect 20637 27829 20671 27863
rect 21465 27829 21499 27863
rect 22845 27829 22879 27863
rect 26433 27829 26467 27863
rect 26525 27829 26559 27863
rect 27537 27829 27571 27863
rect 28733 27829 28767 27863
rect 6101 27625 6135 27659
rect 7573 27625 7607 27659
rect 9505 27625 9539 27659
rect 16773 27625 16807 27659
rect 20637 27625 20671 27659
rect 22293 27625 22327 27659
rect 25605 27625 25639 27659
rect 34529 27625 34563 27659
rect 3617 27557 3651 27591
rect 12173 27557 12207 27591
rect 12633 27557 12667 27591
rect 23949 27557 23983 27591
rect 2237 27489 2271 27523
rect 4445 27489 4479 27523
rect 8493 27489 8527 27523
rect 8585 27489 8619 27523
rect 11621 27489 11655 27523
rect 12817 27489 12851 27523
rect 13369 27489 13403 27523
rect 17325 27489 17359 27523
rect 26157 27489 26191 27523
rect 30113 27489 30147 27523
rect 32781 27489 32815 27523
rect 4721 27421 4755 27455
rect 6193 27421 6227 27455
rect 8953 27421 8987 27455
rect 9045 27421 9079 27455
rect 9229 27421 9263 27455
rect 9321 27421 9355 27455
rect 9597 27421 9631 27455
rect 11805 27421 11839 27455
rect 13461 27421 13495 27455
rect 14565 27421 14599 27455
rect 16037 27421 16071 27455
rect 16221 27421 16255 27455
rect 16405 27421 16439 27455
rect 17141 27421 17175 27455
rect 19073 27421 19107 27455
rect 19257 27421 19291 27455
rect 20913 27421 20947 27455
rect 22385 27421 22419 27455
rect 22661 27421 22695 27455
rect 23305 27421 23339 27455
rect 23489 27421 23523 27455
rect 23581 27421 23615 27455
rect 23673 27421 23707 27455
rect 24133 27421 24167 27455
rect 25973 27421 26007 27455
rect 27169 27421 27203 27455
rect 27445 27421 27479 27455
rect 27905 27421 27939 27455
rect 28917 27421 28951 27455
rect 29009 27421 29043 27455
rect 29193 27421 29227 27455
rect 31585 27421 31619 27455
rect 2504 27353 2538 27387
rect 4261 27353 4295 27387
rect 4988 27353 5022 27387
rect 6460 27353 6494 27387
rect 8401 27353 8435 27387
rect 9864 27353 9898 27387
rect 11713 27353 11747 27387
rect 13553 27353 13587 27387
rect 14832 27353 14866 27387
rect 16313 27353 16347 27387
rect 18828 27353 18862 27387
rect 19524 27353 19558 27387
rect 21180 27353 21214 27387
rect 25421 27353 25455 27387
rect 26065 27353 26099 27387
rect 28641 27353 28675 27387
rect 33057 27353 33091 27387
rect 3893 27285 3927 27319
rect 4353 27285 4387 27319
rect 8033 27285 8067 27319
rect 10977 27285 11011 27319
rect 12357 27285 12391 27319
rect 13921 27285 13955 27319
rect 14105 27285 14139 27319
rect 15945 27285 15979 27319
rect 16589 27285 16623 27319
rect 17233 27285 17267 27319
rect 17693 27285 17727 27319
rect 23857 27285 23891 27319
rect 27261 27285 27295 27319
rect 27629 27285 27663 27319
rect 27721 27285 27755 27319
rect 27997 27285 28031 27319
rect 28733 27285 28767 27319
rect 29377 27285 29411 27319
rect 29561 27285 29595 27319
rect 29929 27285 29963 27319
rect 30021 27285 30055 27319
rect 2605 27081 2639 27115
rect 2973 27081 3007 27115
rect 4813 27081 4847 27115
rect 6837 27081 6871 27115
rect 7205 27081 7239 27115
rect 9321 27081 9355 27115
rect 10149 27081 10183 27115
rect 10517 27081 10551 27115
rect 12357 27081 12391 27115
rect 14749 27081 14783 27115
rect 17049 27081 17083 27115
rect 18613 27081 18647 27115
rect 18981 27081 19015 27115
rect 26617 27081 26651 27115
rect 26985 27081 27019 27115
rect 28549 27081 28583 27115
rect 33793 27081 33827 27115
rect 34161 27081 34195 27115
rect 3700 27013 3734 27047
rect 11805 27013 11839 27047
rect 11897 27013 11931 27047
rect 12817 27013 12851 27047
rect 13277 27013 13311 27047
rect 13636 27013 13670 27047
rect 15945 27013 15979 27047
rect 17509 27013 17543 27047
rect 21833 27013 21867 27047
rect 25513 27013 25547 27047
rect 31769 27013 31803 27047
rect 7297 26945 7331 26979
rect 7941 26945 7975 26979
rect 8197 26945 8231 26979
rect 10057 26945 10091 26979
rect 10609 26945 10643 26979
rect 11713 26945 11747 26979
rect 12081 26945 12115 26979
rect 12587 26945 12621 26979
rect 12725 26945 12759 26979
rect 13000 26945 13034 26979
rect 13093 26945 13127 26979
rect 14841 26945 14875 26979
rect 17141 26945 17175 26979
rect 17289 26945 17323 26979
rect 17417 26945 17451 26979
rect 17606 26945 17640 26979
rect 18153 26945 18187 26979
rect 19993 26945 20027 26979
rect 20177 26945 20211 26979
rect 20545 26945 20579 26979
rect 22017 26945 22051 26979
rect 22560 26945 22594 26979
rect 24041 26945 24075 26979
rect 24308 26945 24342 26979
rect 26709 26945 26743 26979
rect 28098 26945 28132 26979
rect 28365 26945 28399 26979
rect 29662 26945 29696 26979
rect 29929 26945 29963 26979
rect 30941 26945 30975 26979
rect 31033 26945 31067 26979
rect 33977 26945 34011 26979
rect 34253 26945 34287 26979
rect 34529 26945 34563 26979
rect 3065 26877 3099 26911
rect 3249 26877 3283 26911
rect 3433 26877 3467 26911
rect 7481 26877 7515 26911
rect 10701 26877 10735 26911
rect 13369 26877 13403 26911
rect 17969 26877 18003 26911
rect 18337 26877 18371 26911
rect 18521 26877 18555 26911
rect 20269 26877 20303 26911
rect 20361 26877 20395 26911
rect 20913 26877 20947 26911
rect 22293 26877 22327 26911
rect 34805 26877 34839 26911
rect 16037 26809 16071 26843
rect 21097 26809 21131 26843
rect 4997 26741 5031 26775
rect 9689 26741 9723 26775
rect 9873 26741 9907 26775
rect 11069 26741 11103 26775
rect 11529 26741 11563 26775
rect 12449 26741 12483 26775
rect 17785 26741 17819 26775
rect 20729 26741 20763 26775
rect 23673 26741 23707 26775
rect 25421 26741 25455 26775
rect 26341 26741 26375 26775
rect 5365 26537 5399 26571
rect 5733 26537 5767 26571
rect 9781 26537 9815 26571
rect 11529 26537 11563 26571
rect 15117 26537 15151 26571
rect 15945 26537 15979 26571
rect 17693 26537 17727 26571
rect 17877 26537 17911 26571
rect 21465 26537 21499 26571
rect 22293 26537 22327 26571
rect 22845 26537 22879 26571
rect 24593 26537 24627 26571
rect 27353 26537 27387 26571
rect 29377 26537 29411 26571
rect 11713 26469 11747 26503
rect 12081 26469 12115 26503
rect 17417 26469 17451 26503
rect 26341 26469 26375 26503
rect 11345 26401 11379 26435
rect 15669 26401 15703 26435
rect 21925 26401 21959 26435
rect 22017 26401 22051 26435
rect 22753 26401 22787 26435
rect 23397 26401 23431 26435
rect 25237 26401 25271 26435
rect 26709 26401 26743 26435
rect 28917 26401 28951 26435
rect 29009 26401 29043 26435
rect 30113 26401 30147 26435
rect 1501 26333 1535 26367
rect 1961 26333 1995 26367
rect 3525 26333 3559 26367
rect 5549 26333 5583 26367
rect 11529 26333 11563 26367
rect 13461 26333 13495 26367
rect 15485 26333 15519 26367
rect 16773 26333 16807 26367
rect 16866 26333 16900 26367
rect 17049 26333 17083 26367
rect 17141 26333 17175 26367
rect 17279 26333 17313 26367
rect 17509 26333 17543 26367
rect 17601 26333 17635 26367
rect 18061 26333 18095 26367
rect 18245 26333 18279 26367
rect 21833 26333 21867 26367
rect 23213 26333 23247 26367
rect 24961 26333 24995 26367
rect 25421 26333 25455 26367
rect 25514 26333 25548 26367
rect 25789 26333 25823 26367
rect 25886 26333 25920 26367
rect 26249 26333 26283 26367
rect 26893 26333 26927 26367
rect 26985 26333 27019 26367
rect 28641 26333 28675 26367
rect 28825 26333 28859 26367
rect 29193 26333 29227 26367
rect 29653 26333 29687 26367
rect 33977 26333 34011 26367
rect 34253 26333 34287 26367
rect 1685 26265 1719 26299
rect 1869 26265 1903 26299
rect 3801 26265 3835 26299
rect 7481 26265 7515 26299
rect 11253 26265 11287 26299
rect 13194 26265 13228 26299
rect 14933 26265 14967 26299
rect 15577 26265 15611 26299
rect 23305 26265 23339 26299
rect 25697 26265 25731 26299
rect 30380 26265 30414 26299
rect 34161 26265 34195 26299
rect 3341 26197 3375 26231
rect 9045 26197 9079 26231
rect 13645 26197 13679 26231
rect 25053 26197 25087 26231
rect 26065 26197 26099 26231
rect 31493 26197 31527 26231
rect 33793 26197 33827 26231
rect 4537 25993 4571 26027
rect 5457 25993 5491 26027
rect 10609 25993 10643 26027
rect 12541 25993 12575 26027
rect 13001 25993 13035 26027
rect 13369 25993 13403 26027
rect 15669 25993 15703 26027
rect 16129 25993 16163 26027
rect 16405 25993 16439 26027
rect 16681 25993 16715 26027
rect 18797 25993 18831 26027
rect 20269 25993 20303 26027
rect 26525 25993 26559 26027
rect 29837 25993 29871 26027
rect 30297 25993 30331 26027
rect 30665 25993 30699 26027
rect 34989 25993 35023 26027
rect 3985 25925 4019 25959
rect 8033 25925 8067 25959
rect 9229 25925 9263 25959
rect 12909 25925 12943 25959
rect 19901 25925 19935 25959
rect 33517 25925 33551 25959
rect 4813 25857 4847 25891
rect 4906 25857 4940 25891
rect 5089 25857 5123 25891
rect 5181 25857 5215 25891
rect 5319 25857 5353 25891
rect 5733 25857 5767 25891
rect 6837 25857 6871 25891
rect 7941 25857 7975 25891
rect 8493 25857 8527 25891
rect 8585 25857 8619 25891
rect 9321 25857 9355 25891
rect 9965 25857 9999 25891
rect 10058 25857 10092 25891
rect 10241 25857 10275 25891
rect 10333 25857 10367 25891
rect 10471 25857 10505 25891
rect 14105 25857 14139 25891
rect 14372 25857 14406 25891
rect 15853 25857 15887 25891
rect 17794 25857 17828 25891
rect 18705 25857 18739 25891
rect 19625 25857 19659 25891
rect 19718 25857 19752 25891
rect 19993 25857 20027 25891
rect 20131 25857 20165 25891
rect 21925 25857 21959 25891
rect 24317 25857 24351 25891
rect 24584 25857 24618 25891
rect 25973 25857 26007 25891
rect 4077 25789 4111 25823
rect 4169 25789 4203 25823
rect 6561 25789 6595 25823
rect 8125 25789 8159 25823
rect 9413 25789 9447 25823
rect 10701 25789 10735 25823
rect 10977 25789 11011 25823
rect 13185 25789 13219 25823
rect 18061 25789 18095 25823
rect 18889 25789 18923 25823
rect 19165 25789 19199 25823
rect 30757 25789 30791 25823
rect 30849 25789 30883 25823
rect 33241 25789 33275 25823
rect 5917 25721 5951 25755
rect 25789 25721 25823 25755
rect 3617 25653 3651 25687
rect 5549 25653 5583 25687
rect 6101 25653 6135 25687
rect 7573 25653 7607 25687
rect 8769 25653 8803 25687
rect 8861 25653 8895 25687
rect 9781 25653 9815 25687
rect 15485 25653 15519 25687
rect 16037 25653 16071 25687
rect 18337 25653 18371 25687
rect 20453 25653 20487 25687
rect 22109 25653 22143 25687
rect 22293 25653 22327 25687
rect 22477 25653 22511 25687
rect 25697 25653 25731 25687
rect 30113 25653 30147 25687
rect 5273 25449 5307 25483
rect 8217 25449 8251 25483
rect 9505 25449 9539 25483
rect 13001 25449 13035 25483
rect 14657 25449 14691 25483
rect 16037 25449 16071 25483
rect 16313 25449 16347 25483
rect 17141 25449 17175 25483
rect 19073 25449 19107 25483
rect 24869 25449 24903 25483
rect 25881 25449 25915 25483
rect 22385 25381 22419 25415
rect 29377 25381 29411 25415
rect 3893 25313 3927 25347
rect 15301 25313 15335 25347
rect 16589 25313 16623 25347
rect 16681 25313 16715 25347
rect 17693 25313 17727 25347
rect 25421 25313 25455 25347
rect 30021 25313 30055 25347
rect 30205 25313 30239 25347
rect 5365 25245 5399 25279
rect 6837 25245 6871 25279
rect 7104 25245 7138 25279
rect 8953 25245 8987 25279
rect 9229 25245 9263 25279
rect 9321 25245 9355 25279
rect 9689 25245 9723 25279
rect 11621 25245 11655 25279
rect 15485 25245 15519 25279
rect 15761 25245 15795 25279
rect 15853 25245 15887 25279
rect 16773 25245 16807 25279
rect 17960 25245 17994 25279
rect 19349 25245 19383 25279
rect 20913 25245 20947 25279
rect 22569 25245 22603 25279
rect 26341 25245 26375 25279
rect 27997 25245 28031 25279
rect 29929 25245 29963 25279
rect 30389 25245 30423 25279
rect 30482 25245 30516 25279
rect 30757 25245 30791 25279
rect 30895 25245 30929 25279
rect 4160 25177 4194 25211
rect 5632 25177 5666 25211
rect 9137 25177 9171 25211
rect 9956 25177 9990 25211
rect 11888 25177 11922 25211
rect 15025 25177 15059 25211
rect 15669 25177 15703 25211
rect 19616 25177 19650 25211
rect 21180 25177 21214 25211
rect 22836 25177 22870 25211
rect 24041 25177 24075 25211
rect 25237 25177 25271 25211
rect 26608 25177 26642 25211
rect 28264 25177 28298 25211
rect 30665 25177 30699 25211
rect 31125 25177 31159 25211
rect 6745 25109 6779 25143
rect 8585 25109 8619 25143
rect 11069 25109 11103 25143
rect 15117 25109 15151 25143
rect 17325 25109 17359 25143
rect 20729 25109 20763 25143
rect 22293 25109 22327 25143
rect 23949 25109 23983 25143
rect 24685 25109 24719 25143
rect 25329 25109 25363 25143
rect 25697 25109 25731 25143
rect 26249 25109 26283 25143
rect 27721 25109 27755 25143
rect 29561 25109 29595 25143
rect 31033 25109 31067 25143
rect 31309 25109 31343 25143
rect 4261 24905 4295 24939
rect 4537 24905 4571 24939
rect 4905 24905 4939 24939
rect 6377 24905 6411 24939
rect 6745 24905 6779 24939
rect 9689 24905 9723 24939
rect 10149 24905 10183 24939
rect 10517 24905 10551 24939
rect 11069 24905 11103 24939
rect 15117 24905 15151 24939
rect 15577 24905 15611 24939
rect 19717 24905 19751 24939
rect 20085 24905 20119 24939
rect 21833 24905 21867 24939
rect 22201 24905 22235 24939
rect 23121 24905 23155 24939
rect 25237 24905 25271 24939
rect 26985 24905 27019 24939
rect 27353 24905 27387 24939
rect 27813 24905 27847 24939
rect 30113 24905 30147 24939
rect 30389 24905 30423 24939
rect 8576 24837 8610 24871
rect 10609 24837 10643 24871
rect 23489 24837 23523 24871
rect 24225 24837 24259 24871
rect 28641 24837 28675 24871
rect 2881 24769 2915 24803
rect 3148 24769 3182 24803
rect 4997 24769 5031 24803
rect 6837 24769 6871 24803
rect 13645 24769 13679 24803
rect 13737 24769 13771 24803
rect 14004 24769 14038 24803
rect 15669 24769 15703 24803
rect 17049 24769 17083 24803
rect 17141 24769 17175 24803
rect 17509 24769 17543 24803
rect 20177 24769 20211 24803
rect 22293 24769 22327 24803
rect 22937 24769 22971 24803
rect 23949 24769 23983 24803
rect 24042 24769 24076 24803
rect 24317 24769 24351 24803
rect 24414 24769 24448 24803
rect 24685 24769 24719 24803
rect 25053 24769 25087 24803
rect 26065 24769 26099 24803
rect 26433 24769 26467 24803
rect 27445 24769 27479 24803
rect 29009 24769 29043 24803
rect 29285 24769 29319 24803
rect 29929 24769 29963 24803
rect 30481 24769 30515 24803
rect 30665 24769 30699 24803
rect 30849 24769 30883 24803
rect 31217 24769 31251 24803
rect 5181 24701 5215 24735
rect 7021 24701 7055 24735
rect 8309 24701 8343 24735
rect 10793 24701 10827 24735
rect 15761 24701 15795 24735
rect 16037 24701 16071 24735
rect 17233 24701 17267 24735
rect 20361 24701 20395 24735
rect 22385 24701 22419 24735
rect 23581 24701 23615 24735
rect 23765 24701 23799 24735
rect 26525 24701 26559 24735
rect 27537 24701 27571 24735
rect 29101 24701 29135 24735
rect 30941 24701 30975 24735
rect 31033 24701 31067 24735
rect 15209 24633 15243 24667
rect 17693 24633 17727 24667
rect 24593 24633 24627 24667
rect 26801 24633 26835 24667
rect 12357 24565 12391 24599
rect 16681 24565 16715 24599
rect 17785 24565 17819 24599
rect 22753 24565 22787 24599
rect 24869 24565 24903 24599
rect 25421 24565 25455 24599
rect 25605 24565 25639 24599
rect 25881 24565 25915 24599
rect 26249 24565 26283 24599
rect 26433 24565 26467 24599
rect 27997 24565 28031 24599
rect 28181 24565 28215 24599
rect 28365 24565 28399 24599
rect 28825 24565 28859 24599
rect 29745 24565 29779 24599
rect 31401 24565 31435 24599
rect 31493 24565 31527 24599
rect 10057 24361 10091 24395
rect 12173 24361 12207 24395
rect 14197 24361 14231 24395
rect 17325 24361 17359 24395
rect 19809 24361 19843 24395
rect 19901 24361 19935 24395
rect 22753 24361 22787 24395
rect 26709 24361 26743 24395
rect 26893 24361 26927 24395
rect 28549 24361 28583 24395
rect 28733 24361 28767 24395
rect 29929 24361 29963 24395
rect 31769 24361 31803 24395
rect 3985 24293 4019 24327
rect 7021 24293 7055 24327
rect 13093 24293 13127 24327
rect 21741 24293 21775 24327
rect 22661 24293 22695 24327
rect 23213 24293 23247 24327
rect 23857 24293 23891 24327
rect 26433 24293 26467 24327
rect 6745 24225 6779 24259
rect 12817 24225 12851 24259
rect 25421 24225 25455 24259
rect 1409 24157 1443 24191
rect 1685 24157 1719 24191
rect 3801 24157 3835 24191
rect 4721 24157 4755 24191
rect 9137 24157 9171 24191
rect 11621 24157 11655 24191
rect 12541 24157 12575 24191
rect 12633 24157 12667 24191
rect 15945 24157 15979 24191
rect 19257 24157 19291 24191
rect 19625 24157 19659 24191
rect 20085 24157 20119 24191
rect 21925 24157 21959 24191
rect 22109 24157 22143 24191
rect 22385 24157 22419 24191
rect 22477 24157 22511 24191
rect 23305 24157 23339 24191
rect 23489 24157 23523 24191
rect 25237 24157 25271 24191
rect 25789 24157 25823 24191
rect 25937 24157 25971 24191
rect 26065 24157 26099 24191
rect 26254 24157 26288 24191
rect 26525 24157 26559 24191
rect 27072 24157 27106 24191
rect 27261 24157 27295 24191
rect 27389 24157 27423 24191
rect 27537 24157 27571 24191
rect 27629 24157 27663 24191
rect 27997 24157 28031 24191
rect 28365 24157 28399 24191
rect 28917 24157 28951 24191
rect 29653 24157 29687 24191
rect 29745 24157 29779 24191
rect 30389 24157 30423 24191
rect 32781 24157 32815 24191
rect 4261 24089 4295 24123
rect 16212 24089 16246 24123
rect 19441 24089 19475 24123
rect 19533 24089 19567 24123
rect 20177 24089 20211 24123
rect 22293 24089 22327 24123
rect 24409 24089 24443 24123
rect 26157 24089 26191 24123
rect 27169 24089 27203 24123
rect 29009 24089 29043 24123
rect 30021 24089 30055 24123
rect 30656 24089 30690 24123
rect 33057 24089 33091 24123
rect 1593 24021 1627 24055
rect 4905 24021 4939 24055
rect 6101 24021 6135 24055
rect 6469 24021 6503 24055
rect 6561 24021 6595 24055
rect 11437 24021 11471 24055
rect 13737 24021 13771 24055
rect 22937 24021 22971 24055
rect 23673 24021 23707 24055
rect 24041 24021 24075 24055
rect 24685 24021 24719 24055
rect 24869 24021 24903 24055
rect 25329 24021 25363 24055
rect 27813 24021 27847 24055
rect 28181 24021 28215 24055
rect 29193 24021 29227 24055
rect 34529 24021 34563 24055
rect 5365 23817 5399 23851
rect 5825 23817 5859 23851
rect 11529 23817 11563 23851
rect 12449 23817 12483 23851
rect 13277 23817 13311 23851
rect 13553 23817 13587 23851
rect 13829 23817 13863 23851
rect 20361 23817 20395 23851
rect 23949 23817 23983 23851
rect 25973 23817 26007 23851
rect 28457 23817 28491 23851
rect 30021 23817 30055 23851
rect 30665 23817 30699 23851
rect 31033 23817 31067 23851
rect 31125 23817 31159 23851
rect 33977 23817 34011 23851
rect 4160 23749 4194 23783
rect 6469 23749 6503 23783
rect 10232 23749 10266 23783
rect 15669 23749 15703 23783
rect 19248 23749 19282 23783
rect 21833 23749 21867 23783
rect 34345 23749 34379 23783
rect 34805 23749 34839 23783
rect 2421 23681 2455 23715
rect 2688 23681 2722 23715
rect 3893 23681 3927 23715
rect 5733 23681 5767 23715
rect 6653 23681 6687 23715
rect 6920 23681 6954 23715
rect 8309 23681 8343 23715
rect 8493 23681 8527 23715
rect 8760 23681 8794 23715
rect 9965 23681 9999 23715
rect 11897 23681 11931 23715
rect 13461 23681 13495 23715
rect 15485 23681 15519 23715
rect 17417 23681 17451 23715
rect 17684 23681 17718 23715
rect 18981 23681 19015 23715
rect 21281 23681 21315 23715
rect 22569 23681 22603 23715
rect 22836 23681 22870 23715
rect 24501 23681 24535 23715
rect 24685 23681 24719 23715
rect 26525 23681 26559 23715
rect 26985 23681 27019 23715
rect 27252 23681 27286 23715
rect 28908 23681 28942 23715
rect 34161 23681 34195 23715
rect 34437 23681 34471 23715
rect 34529 23681 34563 23715
rect 6009 23613 6043 23647
rect 11989 23613 12023 23647
rect 12173 23613 12207 23647
rect 15853 23613 15887 23647
rect 21097 23613 21131 23647
rect 21189 23613 21223 23647
rect 28641 23613 28675 23647
rect 31217 23613 31251 23647
rect 31493 23613 31527 23647
rect 8125 23545 8159 23579
rect 11345 23545 11379 23579
rect 3801 23477 3835 23511
rect 5273 23477 5307 23511
rect 8033 23477 8067 23511
rect 9873 23477 9907 23511
rect 15301 23477 15335 23511
rect 18797 23477 18831 23511
rect 21649 23477 21683 23511
rect 26709 23477 26743 23511
rect 28365 23477 28399 23511
rect 5273 23273 5307 23307
rect 10609 23273 10643 23307
rect 10885 23273 10919 23307
rect 11805 23273 11839 23307
rect 11989 23273 12023 23307
rect 17969 23273 18003 23307
rect 23029 23273 23063 23307
rect 25789 23273 25823 23307
rect 26433 23273 26467 23307
rect 26525 23273 26559 23307
rect 27169 23273 27203 23307
rect 29561 23273 29595 23307
rect 6837 23205 6871 23239
rect 7205 23205 7239 23239
rect 8677 23205 8711 23239
rect 16773 23205 16807 23239
rect 17141 23205 17175 23239
rect 26985 23205 27019 23239
rect 4261 23137 4295 23171
rect 7665 23137 7699 23171
rect 7757 23137 7791 23171
rect 9781 23137 9815 23171
rect 18981 23137 19015 23171
rect 23489 23137 23523 23171
rect 23581 23137 23615 23171
rect 23857 23137 23891 23171
rect 27721 23137 27755 23171
rect 30113 23137 30147 23171
rect 30389 23137 30423 23171
rect 5089 23069 5123 23103
rect 5457 23069 5491 23103
rect 5724 23069 5758 23103
rect 7573 23069 7607 23103
rect 8033 23069 8067 23103
rect 8126 23069 8160 23103
rect 8401 23069 8435 23103
rect 8539 23069 8573 23103
rect 8953 23069 8987 23103
rect 10149 23069 10183 23103
rect 10241 23069 10275 23103
rect 10425 23069 10459 23103
rect 10517 23069 10551 23103
rect 11069 23069 11103 23103
rect 11253 23069 11287 23103
rect 11345 23069 11379 23103
rect 11437 23069 11471 23103
rect 12173 23069 12207 23103
rect 14289 23069 14323 23103
rect 15761 23069 15795 23103
rect 15854 23069 15888 23103
rect 16226 23069 16260 23103
rect 16589 23069 16623 23103
rect 16957 23069 16991 23103
rect 18153 23069 18187 23103
rect 19257 23069 19291 23103
rect 21465 23069 21499 23103
rect 21732 23069 21766 23103
rect 23397 23069 23431 23103
rect 24409 23069 24443 23103
rect 27537 23069 27571 23103
rect 29377 23069 29411 23103
rect 29929 23069 29963 23103
rect 8309 23001 8343 23035
rect 12440 23001 12474 23035
rect 14556 23001 14590 23035
rect 16037 23001 16071 23035
rect 16129 23001 16163 23035
rect 24676 23001 24710 23035
rect 27629 23001 27663 23035
rect 29009 23001 29043 23035
rect 30021 23001 30055 23035
rect 9965 22933 9999 22967
rect 11621 22933 11655 22967
rect 13553 22933 13587 22967
rect 15669 22933 15703 22967
rect 16405 22933 16439 22967
rect 22845 22933 22879 22967
rect 24041 22933 24075 22967
rect 26709 22933 26743 22967
rect 29193 22933 29227 22967
rect 3801 22729 3835 22763
rect 4261 22729 4295 22763
rect 5457 22729 5491 22763
rect 8585 22729 8619 22763
rect 8861 22729 8895 22763
rect 9045 22729 9079 22763
rect 9413 22729 9447 22763
rect 12725 22729 12759 22763
rect 14105 22729 14139 22763
rect 14841 22729 14875 22763
rect 15209 22729 15243 22763
rect 17509 22729 17543 22763
rect 17969 22729 18003 22763
rect 18337 22729 18371 22763
rect 18429 22729 18463 22763
rect 19349 22729 19383 22763
rect 19717 22729 19751 22763
rect 26341 22729 26375 22763
rect 27813 22729 27847 22763
rect 29101 22729 29135 22763
rect 4997 22661 5031 22695
rect 5089 22661 5123 22695
rect 7941 22661 7975 22695
rect 13737 22661 13771 22695
rect 14197 22661 14231 22695
rect 19809 22661 19843 22695
rect 21005 22661 21039 22695
rect 34345 22661 34379 22695
rect 1501 22593 1535 22627
rect 1961 22593 1995 22627
rect 4169 22593 4203 22627
rect 4813 22593 4847 22627
rect 5181 22593 5215 22627
rect 8217 22593 8251 22627
rect 9505 22593 9539 22627
rect 9873 22593 9907 22627
rect 10140 22593 10174 22627
rect 13093 22593 13127 22627
rect 13553 22593 13587 22627
rect 13829 22593 13863 22627
rect 13921 22593 13955 22627
rect 14381 22593 14415 22627
rect 16497 22593 16531 22627
rect 16681 22593 16715 22627
rect 16865 22593 16899 22627
rect 17233 22593 17267 22627
rect 20637 22593 20671 22627
rect 21833 22593 21867 22627
rect 24777 22593 24811 22627
rect 24961 22593 24995 22627
rect 25228 22593 25262 22627
rect 27077 22593 27111 22627
rect 27997 22593 28031 22627
rect 28273 22593 28307 22627
rect 28917 22593 28951 22627
rect 30582 22593 30616 22627
rect 30849 22593 30883 22627
rect 31401 22593 31435 22627
rect 34161 22593 34195 22627
rect 34437 22593 34471 22627
rect 34529 22593 34563 22627
rect 4353 22525 4387 22559
rect 8033 22525 8067 22559
rect 9597 22525 9631 22559
rect 13185 22525 13219 22559
rect 13277 22525 13311 22559
rect 15301 22525 15335 22559
rect 15485 22525 15519 22559
rect 16221 22525 16255 22559
rect 16957 22525 16991 22559
rect 17049 22525 17083 22559
rect 17693 22525 17727 22559
rect 18613 22525 18647 22559
rect 19901 22525 19935 22559
rect 22201 22525 22235 22559
rect 34805 22525 34839 22559
rect 1685 22457 1719 22491
rect 1869 22457 1903 22491
rect 5365 22457 5399 22491
rect 8401 22457 8435 22491
rect 20177 22457 20211 22491
rect 4721 22389 4755 22423
rect 5733 22389 5767 22423
rect 7941 22389 7975 22423
rect 8769 22389 8803 22423
rect 11253 22389 11287 22423
rect 17417 22389 17451 22423
rect 19165 22389 19199 22423
rect 20453 22389 20487 22423
rect 20729 22389 20763 22423
rect 22017 22389 22051 22423
rect 29285 22389 29319 22423
rect 29469 22389 29503 22423
rect 33977 22389 34011 22423
rect 13645 22185 13679 22219
rect 25513 22185 25547 22219
rect 26433 22185 26467 22219
rect 29193 22185 29227 22219
rect 30573 22185 30607 22219
rect 33044 22185 33078 22219
rect 34529 22185 34563 22219
rect 15669 22117 15703 22151
rect 17509 22117 17543 22151
rect 22201 22117 22235 22151
rect 23765 22117 23799 22151
rect 28457 22117 28491 22151
rect 4353 22049 4387 22083
rect 11069 22049 11103 22083
rect 11345 22049 11379 22083
rect 15393 22049 15427 22083
rect 19533 22049 19567 22083
rect 20821 22049 20855 22083
rect 22845 22049 22879 22083
rect 25973 22049 26007 22083
rect 26157 22049 26191 22083
rect 26525 22049 26559 22083
rect 31125 22049 31159 22083
rect 32781 22049 32815 22083
rect 4629 21981 4663 22015
rect 4813 21981 4847 22015
rect 4905 21981 4939 22015
rect 4997 21981 5031 22015
rect 5273 21981 5307 22015
rect 10793 21981 10827 22015
rect 12173 21981 12207 22015
rect 16129 21981 16163 22015
rect 18337 21981 18371 22015
rect 18613 21981 18647 22015
rect 19257 21981 19291 22015
rect 20177 21981 20211 22015
rect 20637 21981 20671 22015
rect 22661 21981 22695 22015
rect 24225 21981 24259 22015
rect 24501 21981 24535 22015
rect 27077 21981 27111 22015
rect 28549 21981 28583 22015
rect 28733 21981 28767 22015
rect 28825 21981 28859 22015
rect 28963 21981 28997 22015
rect 29377 21981 29411 22015
rect 29561 21981 29595 22015
rect 30941 21981 30975 22015
rect 9873 21913 9907 21947
rect 10885 21913 10919 21947
rect 12440 21913 12474 21947
rect 15301 21913 15335 21947
rect 16396 21913 16430 21947
rect 18245 21913 18279 21947
rect 21088 21913 21122 21947
rect 22753 21913 22787 21947
rect 25237 21913 25271 21947
rect 25881 21913 25915 21947
rect 27344 21913 27378 21947
rect 30297 21913 30331 21947
rect 3801 21845 3835 21879
rect 4169 21845 4203 21879
rect 4261 21845 4295 21879
rect 5181 21845 5215 21879
rect 10425 21845 10459 21879
rect 13553 21845 13587 21879
rect 14841 21845 14875 21879
rect 15209 21845 15243 21879
rect 15853 21845 15887 21879
rect 18521 21845 18555 21879
rect 18797 21845 18831 21879
rect 18981 21845 19015 21879
rect 20361 21845 20395 21879
rect 22293 21845 22327 21879
rect 23121 21845 23155 21879
rect 24041 21845 24075 21879
rect 29101 21845 29135 21879
rect 31033 21845 31067 21879
rect 31401 21845 31435 21879
rect 1869 21641 1903 21675
rect 4721 21641 4755 21675
rect 7941 21641 7975 21675
rect 8401 21641 8435 21675
rect 9873 21641 9907 21675
rect 10885 21641 10919 21675
rect 12817 21641 12851 21675
rect 13185 21641 13219 21675
rect 15669 21641 15703 21675
rect 16681 21641 16715 21675
rect 17049 21641 17083 21675
rect 17141 21641 17175 21675
rect 18981 21641 19015 21675
rect 21189 21641 21223 21675
rect 22109 21641 22143 21675
rect 23029 21641 23063 21675
rect 24777 21641 24811 21675
rect 25237 21641 25271 21675
rect 26065 21641 26099 21675
rect 27537 21641 27571 21675
rect 27629 21641 27663 21675
rect 27997 21641 28031 21675
rect 29469 21641 29503 21675
rect 29745 21641 29779 21675
rect 29929 21641 29963 21675
rect 3004 21573 3038 21607
rect 7604 21573 7638 21607
rect 13277 21573 13311 21607
rect 14556 21573 14590 21607
rect 15761 21573 15795 21607
rect 20729 21573 20763 21607
rect 22661 21573 22695 21607
rect 23121 21573 23155 21607
rect 23572 21573 23606 21607
rect 26157 21573 26191 21607
rect 28733 21573 28767 21607
rect 29285 21573 29319 21607
rect 3249 21505 3283 21539
rect 3341 21505 3375 21539
rect 3608 21505 3642 21539
rect 5080 21505 5114 21539
rect 7849 21505 7883 21539
rect 8309 21505 8343 21539
rect 10241 21505 10275 21539
rect 16129 21505 16163 21539
rect 17601 21505 17635 21539
rect 17868 21505 17902 21539
rect 19073 21505 19107 21539
rect 19340 21505 19374 21539
rect 20545 21505 20579 21539
rect 20821 21505 20855 21539
rect 20913 21505 20947 21539
rect 22293 21505 22327 21539
rect 22385 21505 22419 21539
rect 22478 21505 22512 21539
rect 22753 21505 22787 21539
rect 22891 21505 22925 21539
rect 25145 21505 25179 21539
rect 25605 21505 25639 21539
rect 28636 21505 28670 21539
rect 28825 21505 28859 21539
rect 28953 21505 28987 21539
rect 29101 21505 29135 21539
rect 30297 21505 30331 21539
rect 4813 21437 4847 21471
rect 8585 21437 8619 21471
rect 13369 21437 13403 21471
rect 13645 21437 13679 21471
rect 14289 21437 14323 21471
rect 17325 21437 17359 21471
rect 23305 21437 23339 21471
rect 25421 21437 25455 21471
rect 28089 21437 28123 21471
rect 28181 21437 28215 21471
rect 30389 21437 30423 21471
rect 30481 21437 30515 21471
rect 21097 21369 21131 21403
rect 24685 21369 24719 21403
rect 28457 21369 28491 21403
rect 30941 21369 30975 21403
rect 6193 21301 6227 21335
rect 6469 21301 6503 21335
rect 8861 21301 8895 21335
rect 10425 21301 10459 21335
rect 10609 21301 10643 21335
rect 16497 21301 16531 21335
rect 20453 21301 20487 21335
rect 21833 21301 21867 21335
rect 25789 21301 25823 21335
rect 26341 21301 26375 21335
rect 30757 21301 30791 21335
rect 4169 21097 4203 21131
rect 5825 21097 5859 21131
rect 7757 21097 7791 21131
rect 7941 21097 7975 21131
rect 8125 21097 8159 21131
rect 14289 21097 14323 21131
rect 16497 21097 16531 21131
rect 18153 21097 18187 21131
rect 19625 21097 19659 21131
rect 20453 21097 20487 21131
rect 27445 21097 27479 21131
rect 29285 21097 29319 21131
rect 31033 21097 31067 21131
rect 31217 21097 31251 21131
rect 31677 21097 31711 21131
rect 18981 21029 19015 21063
rect 24409 21029 24443 21063
rect 4813 20961 4847 20995
rect 4997 20961 5031 20995
rect 6377 20961 6411 20995
rect 9597 20961 9631 20995
rect 9781 20961 9815 20995
rect 18613 20961 18647 20995
rect 18705 20961 18739 20995
rect 20177 20961 20211 20995
rect 23213 20961 23247 20995
rect 27537 20961 27571 20995
rect 29653 20961 29687 20995
rect 4537 20893 4571 20927
rect 6193 20893 6227 20927
rect 7205 20893 7239 20927
rect 7481 20893 7515 20927
rect 7573 20893 7607 20927
rect 11621 20893 11655 20927
rect 15393 20893 15427 20927
rect 19993 20893 20027 20927
rect 23857 20893 23891 20927
rect 23949 20893 23983 20927
rect 24225 20893 24259 20927
rect 24593 20893 24627 20927
rect 26065 20893 26099 20927
rect 29101 20893 29135 20927
rect 29920 20893 29954 20927
rect 31401 20893 31435 20927
rect 34529 20893 34563 20927
rect 4629 20825 4663 20859
rect 6285 20825 6319 20859
rect 7389 20825 7423 20859
rect 10048 20825 10082 20859
rect 11888 20825 11922 20859
rect 14565 20825 14599 20859
rect 15485 20825 15519 20859
rect 17601 20825 17635 20859
rect 22946 20825 22980 20859
rect 24041 20825 24075 20859
rect 24860 20825 24894 20859
rect 26332 20825 26366 20859
rect 27804 20825 27838 20859
rect 31493 20825 31527 20859
rect 34253 20825 34287 20859
rect 6653 20757 6687 20791
rect 8953 20757 8987 20791
rect 9321 20757 9355 20791
rect 9413 20757 9447 20791
rect 11161 20757 11195 20791
rect 13001 20757 13035 20791
rect 18521 20757 18555 20791
rect 19441 20757 19475 20791
rect 20085 20757 20119 20791
rect 21833 20757 21867 20791
rect 23673 20757 23707 20791
rect 25973 20757 26007 20791
rect 28917 20757 28951 20791
rect 9505 20553 9539 20587
rect 10333 20553 10367 20587
rect 10701 20553 10735 20587
rect 19993 20553 20027 20587
rect 20269 20553 20303 20587
rect 20821 20553 20855 20587
rect 22661 20553 22695 20587
rect 23029 20553 23063 20587
rect 24501 20553 24535 20587
rect 25329 20553 25363 20587
rect 25881 20553 25915 20587
rect 26433 20553 26467 20587
rect 26985 20553 27019 20587
rect 27353 20553 27387 20587
rect 27813 20553 27847 20587
rect 28181 20553 28215 20587
rect 29377 20553 29411 20587
rect 29469 20553 29503 20587
rect 8392 20485 8426 20519
rect 9965 20485 9999 20519
rect 20729 20485 20763 20519
rect 25421 20485 25455 20519
rect 28273 20485 28307 20519
rect 1409 20417 1443 20451
rect 1685 20417 1719 20451
rect 8125 20417 8159 20451
rect 9689 20417 9723 20451
rect 9873 20417 9907 20451
rect 10057 20417 10091 20451
rect 10793 20417 10827 20451
rect 12081 20417 12115 20451
rect 12817 20417 12851 20451
rect 13553 20417 13587 20451
rect 13820 20417 13854 20451
rect 17049 20417 17083 20451
rect 20177 20417 20211 20451
rect 22569 20417 22603 20451
rect 24041 20417 24075 20451
rect 24317 20417 24351 20451
rect 29653 20417 29687 20451
rect 29837 20417 29871 20451
rect 30205 20417 30239 20451
rect 30757 20417 30791 20451
rect 33241 20417 33275 20451
rect 10977 20349 11011 20383
rect 12357 20349 12391 20383
rect 12909 20349 12943 20383
rect 13093 20349 13127 20383
rect 13277 20349 13311 20383
rect 17141 20349 17175 20383
rect 17233 20349 17267 20383
rect 17509 20349 17543 20383
rect 22201 20349 22235 20383
rect 22477 20349 22511 20383
rect 24133 20349 24167 20383
rect 25605 20349 25639 20383
rect 27445 20349 27479 20383
rect 27537 20349 27571 20383
rect 28365 20349 28399 20383
rect 29929 20349 29963 20383
rect 30021 20349 30055 20383
rect 33517 20349 33551 20383
rect 12449 20281 12483 20315
rect 20545 20281 20579 20315
rect 26617 20281 26651 20315
rect 30573 20281 30607 20315
rect 30849 20281 30883 20315
rect 31033 20281 31067 20315
rect 1593 20213 1627 20247
rect 10241 20213 10275 20247
rect 11253 20213 11287 20247
rect 14933 20213 14967 20247
rect 16681 20213 16715 20247
rect 24041 20213 24075 20247
rect 24685 20213 24719 20247
rect 24961 20213 24995 20247
rect 30389 20213 30423 20247
rect 31309 20213 31343 20247
rect 34989 20213 35023 20247
rect 3985 20009 4019 20043
rect 17141 20009 17175 20043
rect 21925 20009 21959 20043
rect 24501 20009 24535 20043
rect 24869 20009 24903 20043
rect 31861 20009 31895 20043
rect 33977 20009 34011 20043
rect 3617 19941 3651 19975
rect 22109 19941 22143 19975
rect 4813 19873 4847 19907
rect 10517 19873 10551 19907
rect 14749 19873 14783 19907
rect 15025 19873 15059 19907
rect 22293 19873 22327 19907
rect 22845 19873 22879 19907
rect 23029 19873 23063 19907
rect 34713 19873 34747 19907
rect 3433 19805 3467 19839
rect 3801 19805 3835 19839
rect 4721 19805 4755 19839
rect 14473 19805 14507 19839
rect 15761 19805 15795 19839
rect 17693 19805 17727 19839
rect 19257 19805 19291 19839
rect 19441 19805 19475 19839
rect 19625 19805 19659 19839
rect 19901 19805 19935 19839
rect 21373 19805 21407 19839
rect 21465 19805 21499 19839
rect 21649 19805 21683 19839
rect 21741 19805 21775 19839
rect 24685 19805 24719 19839
rect 30757 19805 30791 19839
rect 34161 19805 34195 19839
rect 34437 19805 34471 19839
rect 5080 19737 5114 19771
rect 6285 19737 6319 19771
rect 10425 19737 10459 19771
rect 16028 19737 16062 19771
rect 17960 19737 17994 19771
rect 19533 19737 19567 19771
rect 20168 19737 20202 19771
rect 23857 19737 23891 19771
rect 32045 19737 32079 19771
rect 32229 19737 32263 19771
rect 34345 19737 34379 19771
rect 34897 19737 34931 19771
rect 6193 19669 6227 19703
rect 7205 19669 7239 19703
rect 12909 19669 12943 19703
rect 14105 19669 14139 19703
rect 14565 19669 14599 19703
rect 15209 19669 15243 19703
rect 19073 19669 19107 19703
rect 19809 19669 19843 19703
rect 21281 19669 21315 19703
rect 22385 19669 22419 19703
rect 22753 19669 22787 19703
rect 23213 19669 23247 19703
rect 23765 19669 23799 19703
rect 24041 19669 24075 19703
rect 27721 19669 27755 19703
rect 30573 19669 30607 19703
rect 3801 19465 3835 19499
rect 5181 19465 5215 19499
rect 5365 19465 5399 19499
rect 5825 19465 5859 19499
rect 10517 19465 10551 19499
rect 12909 19465 12943 19499
rect 14105 19465 14139 19499
rect 15117 19465 15151 19499
rect 17509 19465 17543 19499
rect 20821 19465 20855 19499
rect 21281 19465 21315 19499
rect 23213 19465 23247 19499
rect 24041 19465 24075 19499
rect 24409 19465 24443 19499
rect 25053 19465 25087 19499
rect 25973 19465 26007 19499
rect 26341 19465 26375 19499
rect 29101 19465 29135 19499
rect 29377 19465 29411 19499
rect 32321 19465 32355 19499
rect 4169 19397 4203 19431
rect 5733 19397 5767 19431
rect 6653 19397 6687 19431
rect 6745 19397 6779 19431
rect 10057 19397 10091 19431
rect 10609 19397 10643 19431
rect 13185 19397 13219 19431
rect 13277 19397 13311 19431
rect 14749 19397 14783 19431
rect 14841 19397 14875 19431
rect 15945 19397 15979 19431
rect 16957 19397 16991 19431
rect 17049 19397 17083 19431
rect 20269 19397 20303 19431
rect 22100 19397 22134 19431
rect 23673 19397 23707 19431
rect 25513 19397 25547 19431
rect 26065 19397 26099 19431
rect 29009 19397 29043 19431
rect 2329 19329 2363 19363
rect 2596 19329 2630 19363
rect 4629 19329 4663 19363
rect 4813 19329 4847 19363
rect 4905 19329 4939 19363
rect 4997 19329 5031 19363
rect 6377 19329 6411 19363
rect 6470 19329 6504 19363
rect 6883 19329 6917 19363
rect 7656 19329 7690 19363
rect 8861 19329 8895 19363
rect 9045 19329 9079 19363
rect 9137 19329 9171 19363
rect 9229 19329 9263 19363
rect 10333 19329 10367 19363
rect 10793 19329 10827 19363
rect 10885 19329 10919 19363
rect 11069 19329 11103 19363
rect 11161 19329 11195 19363
rect 11529 19329 11563 19363
rect 12449 19329 12483 19363
rect 12541 19329 12575 19363
rect 13093 19329 13127 19363
rect 13461 19329 13495 19363
rect 14013 19329 14047 19363
rect 14565 19329 14599 19363
rect 14933 19329 14967 19363
rect 15853 19329 15887 19363
rect 16681 19329 16715 19363
rect 16774 19329 16808 19363
rect 17187 19329 17221 19363
rect 18153 19329 18187 19363
rect 20361 19329 20395 19363
rect 21189 19329 21223 19363
rect 23489 19329 23523 19363
rect 23765 19329 23799 19363
rect 23857 19329 23891 19363
rect 24961 19329 24995 19363
rect 25697 19329 25731 19363
rect 26182 19329 26216 19363
rect 26591 19329 26625 19363
rect 27537 19329 27571 19363
rect 28365 19329 28399 19363
rect 29653 19329 29687 19363
rect 30021 19329 30055 19363
rect 30757 19329 30791 19363
rect 32137 19329 32171 19363
rect 32413 19329 32447 19363
rect 4261 19261 4295 19295
rect 4445 19261 4479 19295
rect 6009 19261 6043 19295
rect 7389 19261 7423 19295
rect 10149 19261 10183 19295
rect 12725 19261 12759 19295
rect 14289 19261 14323 19295
rect 15301 19261 15335 19295
rect 16037 19261 16071 19295
rect 20177 19261 20211 19295
rect 21465 19261 21499 19295
rect 21833 19261 21867 19295
rect 28733 19261 28767 19295
rect 29218 19261 29252 19295
rect 30113 19261 30147 19295
rect 30481 19261 30515 19295
rect 34529 19261 34563 19295
rect 3709 19193 3743 19227
rect 7021 19193 7055 19227
rect 9413 19193 9447 19227
rect 24225 19193 24259 19227
rect 25513 19193 25547 19227
rect 29469 19193 29503 19227
rect 7297 19125 7331 19159
rect 8769 19125 8803 19159
rect 9505 19125 9539 19159
rect 9781 19125 9815 19159
rect 10057 19125 10091 19159
rect 11253 19125 11287 19159
rect 12081 19125 12115 19159
rect 13645 19125 13679 19159
rect 15485 19125 15519 19159
rect 16313 19125 16347 19159
rect 17325 19125 17359 19159
rect 17601 19125 17635 19159
rect 18061 19125 18095 19159
rect 19625 19125 19659 19159
rect 20729 19125 20763 19159
rect 24777 19125 24811 19159
rect 26433 19125 26467 19159
rect 27353 19125 27387 19159
rect 28181 19125 28215 19159
rect 30389 19125 30423 19159
rect 32597 19125 32631 19159
rect 7021 18921 7055 18955
rect 7941 18921 7975 18955
rect 12909 18921 12943 18955
rect 14289 18921 14323 18955
rect 14473 18921 14507 18955
rect 16313 18921 16347 18955
rect 18245 18921 18279 18955
rect 19257 18921 19291 18955
rect 21005 18921 21039 18955
rect 21373 18921 21407 18955
rect 21833 18921 21867 18955
rect 24041 18921 24075 18955
rect 25421 18921 25455 18955
rect 26249 18921 26283 18955
rect 26341 18921 26375 18955
rect 27445 18921 27479 18955
rect 32505 18921 32539 18955
rect 22385 18853 22419 18887
rect 26985 18853 27019 18887
rect 27261 18853 27295 18887
rect 7573 18785 7607 18819
rect 7757 18785 7791 18819
rect 8585 18785 8619 18819
rect 9413 18785 9447 18819
rect 9597 18785 9631 18819
rect 14933 18785 14967 18819
rect 17233 18785 17267 18819
rect 17325 18785 17359 18819
rect 18705 18785 18739 18819
rect 18889 18785 18923 18819
rect 26433 18785 26467 18819
rect 31033 18785 31067 18819
rect 32689 18785 32723 18819
rect 1409 18717 1443 18751
rect 1869 18717 1903 18751
rect 3801 18717 3835 18751
rect 5641 18717 5675 18751
rect 9781 18717 9815 18751
rect 11529 18717 11563 18751
rect 11796 18717 11830 18751
rect 14105 18717 14139 18751
rect 15200 18717 15234 18751
rect 16957 18717 16991 18751
rect 17141 18717 17175 18751
rect 17509 18717 17543 18751
rect 18613 18717 18647 18751
rect 20381 18717 20415 18751
rect 20637 18717 20671 18751
rect 21097 18717 21131 18751
rect 22201 18717 22235 18751
rect 22661 18717 22695 18751
rect 25605 18717 25639 18751
rect 26709 18717 26743 18751
rect 26893 18717 26927 18751
rect 26985 18717 27019 18751
rect 27169 18717 27203 18751
rect 27445 18717 27479 18751
rect 27813 18717 27847 18751
rect 28089 18717 28123 18751
rect 28181 18717 28215 18751
rect 28273 18717 28307 18751
rect 28549 18717 28583 18751
rect 28825 18717 28859 18751
rect 30389 18717 30423 18751
rect 30757 18717 30791 18751
rect 32781 18717 32815 18751
rect 34161 18717 34195 18751
rect 34437 18717 34471 18751
rect 4046 18649 4080 18683
rect 5908 18649 5942 18683
rect 7481 18649 7515 18683
rect 8309 18649 8343 18683
rect 8401 18649 8435 18683
rect 9321 18649 9355 18683
rect 10048 18649 10082 18683
rect 13829 18649 13863 18683
rect 17693 18649 17727 18683
rect 18061 18649 18095 18683
rect 21741 18649 21775 18683
rect 22928 18649 22962 18683
rect 26065 18649 26099 18683
rect 27905 18649 27939 18683
rect 29034 18649 29068 18683
rect 29653 18649 29687 18683
rect 1593 18581 1627 18615
rect 1777 18581 1811 18615
rect 5181 18581 5215 18615
rect 5365 18581 5399 18615
rect 7113 18581 7147 18615
rect 8953 18581 8987 18615
rect 11161 18581 11195 18615
rect 13645 18581 13679 18615
rect 17785 18581 17819 18615
rect 21557 18581 21591 18615
rect 22569 18581 22603 18615
rect 26157 18581 26191 18615
rect 26801 18581 26835 18615
rect 28457 18581 28491 18615
rect 28917 18581 28951 18615
rect 29193 18581 29227 18615
rect 29745 18581 29779 18615
rect 29837 18581 29871 18615
rect 30205 18581 30239 18615
rect 30481 18581 30515 18615
rect 33149 18581 33183 18615
rect 33977 18581 34011 18615
rect 34345 18581 34379 18615
rect 3801 18377 3835 18411
rect 4169 18377 4203 18411
rect 4261 18377 4295 18411
rect 9137 18377 9171 18411
rect 9781 18377 9815 18411
rect 10333 18377 10367 18411
rect 10701 18377 10735 18411
rect 10793 18377 10827 18411
rect 14473 18377 14507 18411
rect 22017 18377 22051 18411
rect 22661 18377 22695 18411
rect 23213 18377 23247 18411
rect 23305 18377 23339 18411
rect 23673 18377 23707 18411
rect 23765 18377 23799 18411
rect 24777 18377 24811 18411
rect 26341 18377 26375 18411
rect 28917 18377 28951 18411
rect 29193 18377 29227 18411
rect 31493 18377 31527 18411
rect 32229 18377 32263 18411
rect 8024 18309 8058 18343
rect 13360 18309 13394 18343
rect 21925 18309 21959 18343
rect 24593 18309 24627 18343
rect 25789 18309 25823 18343
rect 26458 18309 26492 18343
rect 28733 18309 28767 18343
rect 31185 18309 31219 18343
rect 31401 18309 31435 18343
rect 33701 18309 33735 18343
rect 7757 18241 7791 18275
rect 14565 18241 14599 18275
rect 16681 18241 16715 18275
rect 16948 18241 16982 18275
rect 24685 18241 24719 18275
rect 24961 18241 24995 18275
rect 25237 18241 25271 18275
rect 25973 18241 26007 18275
rect 27629 18241 27663 18275
rect 29009 18231 29043 18265
rect 29285 18241 29319 18275
rect 30389 18241 30423 18275
rect 31677 18241 31711 18275
rect 31953 18241 31987 18275
rect 34529 18241 34563 18275
rect 34805 18241 34839 18275
rect 4445 18173 4479 18207
rect 10885 18173 10919 18207
rect 11161 18173 11195 18207
rect 13093 18173 13127 18207
rect 21557 18173 21591 18207
rect 22753 18173 22787 18207
rect 22937 18173 22971 18207
rect 23857 18173 23891 18207
rect 24133 18173 24167 18207
rect 25053 18173 25087 18207
rect 25329 18173 25363 18207
rect 26249 18173 26283 18207
rect 30113 18173 30147 18207
rect 33977 18173 34011 18207
rect 14749 18105 14783 18139
rect 14933 18105 14967 18139
rect 20085 18105 20119 18139
rect 25789 18105 25823 18139
rect 27445 18105 27479 18139
rect 31033 18105 31067 18139
rect 7665 18037 7699 18071
rect 9321 18037 9355 18071
rect 15209 18037 15243 18071
rect 18061 18037 18095 18071
rect 19165 18037 19199 18071
rect 22293 18037 22327 18071
rect 24409 18037 24443 18071
rect 26617 18037 26651 18071
rect 28733 18037 28767 18071
rect 29469 18037 29503 18071
rect 31217 18037 31251 18071
rect 31769 18037 31803 18071
rect 16865 17833 16899 17867
rect 24869 17833 24903 17867
rect 25697 17833 25731 17867
rect 25789 17833 25823 17867
rect 25973 17833 26007 17867
rect 26433 17833 26467 17867
rect 29929 17833 29963 17867
rect 34529 17833 34563 17867
rect 15577 17765 15611 17799
rect 18337 17765 18371 17799
rect 26065 17765 26099 17799
rect 31309 17765 31343 17799
rect 10425 17697 10459 17731
rect 17325 17697 17359 17731
rect 17509 17697 17543 17731
rect 25028 17697 25062 17731
rect 25145 17697 25179 17731
rect 25513 17697 25547 17731
rect 26801 17697 26835 17731
rect 26893 17697 26927 17731
rect 27077 17697 27111 17731
rect 27353 17697 27387 17731
rect 30021 17697 30055 17731
rect 33057 17697 33091 17731
rect 10793 17629 10827 17663
rect 10886 17629 10920 17663
rect 11299 17629 11333 17663
rect 14105 17629 14139 17663
rect 17233 17629 17267 17663
rect 18521 17629 18555 17663
rect 19349 17629 19383 17663
rect 22293 17629 22327 17663
rect 25973 17629 26007 17663
rect 26249 17629 26283 17663
rect 26617 17629 26651 17663
rect 26709 17629 26743 17663
rect 27997 17629 28031 17663
rect 29101 17629 29135 17663
rect 29285 17629 29319 17663
rect 29745 17629 29779 17663
rect 29929 17629 29963 17663
rect 30205 17629 30239 17663
rect 31033 17629 31067 17663
rect 31125 17629 31159 17663
rect 31401 17629 31435 17663
rect 31585 17629 31619 17663
rect 32781 17629 32815 17663
rect 10241 17561 10275 17595
rect 11069 17561 11103 17595
rect 11161 17561 11195 17595
rect 11805 17561 11839 17595
rect 14372 17561 14406 17595
rect 19616 17561 19650 17595
rect 25605 17561 25639 17595
rect 27445 17561 27479 17595
rect 27562 17561 27596 17595
rect 28917 17561 28951 17595
rect 31309 17561 31343 17595
rect 9873 17493 9907 17527
rect 10333 17493 10367 17527
rect 11437 17493 11471 17527
rect 11621 17493 11655 17527
rect 12449 17493 12483 17527
rect 12633 17493 12667 17527
rect 15485 17493 15519 17527
rect 17693 17493 17727 17527
rect 18705 17493 18739 17527
rect 20729 17493 20763 17527
rect 25237 17493 25271 17527
rect 27721 17493 27755 17527
rect 27813 17493 27847 17527
rect 29561 17493 29595 17527
rect 30389 17493 30423 17527
rect 31493 17493 31527 17527
rect 4905 17289 4939 17323
rect 7757 17289 7791 17323
rect 8309 17289 8343 17323
rect 10701 17289 10735 17323
rect 12909 17289 12943 17323
rect 14289 17289 14323 17323
rect 14657 17289 14691 17323
rect 14933 17289 14967 17323
rect 19165 17289 19199 17323
rect 19901 17289 19935 17323
rect 24777 17289 24811 17323
rect 28273 17289 28307 17323
rect 30113 17289 30147 17323
rect 7481 17221 7515 17255
rect 8033 17221 8067 17255
rect 9588 17221 9622 17255
rect 20269 17221 20303 17255
rect 22109 17221 22143 17255
rect 25605 17221 25639 17255
rect 26709 17221 26743 17255
rect 3792 17153 3826 17187
rect 6745 17153 6779 17187
rect 7205 17153 7239 17187
rect 7389 17153 7423 17187
rect 7573 17153 7607 17187
rect 7849 17153 7883 17187
rect 9321 17153 9355 17187
rect 11796 17153 11830 17187
rect 14749 17153 14783 17187
rect 15384 17153 15418 17187
rect 17509 17153 17543 17187
rect 17776 17153 17810 17187
rect 18981 17153 19015 17187
rect 20361 17153 20395 17187
rect 21833 17153 21867 17187
rect 22017 17153 22051 17187
rect 22201 17153 22235 17187
rect 23397 17153 23431 17187
rect 23857 17153 23891 17187
rect 24685 17153 24719 17187
rect 25145 17153 25179 17187
rect 25881 17153 25915 17187
rect 27169 17153 27203 17187
rect 3525 17085 3559 17119
rect 6837 17085 6871 17119
rect 7021 17085 7055 17119
rect 11529 17085 11563 17119
rect 14105 17085 14139 17119
rect 14197 17085 14231 17119
rect 15117 17085 15151 17119
rect 20453 17085 20487 17119
rect 20821 17085 20855 17119
rect 22569 17085 22603 17119
rect 23949 17085 23983 17119
rect 24041 17085 24075 17119
rect 24869 17085 24903 17119
rect 28365 17085 28399 17119
rect 28641 17085 28675 17119
rect 8493 17017 8527 17051
rect 21557 17017 21591 17051
rect 25329 17017 25363 17051
rect 26065 17017 26099 17051
rect 26249 17017 26283 17051
rect 26985 17017 27019 17051
rect 6377 16949 6411 16983
rect 10793 16949 10827 16983
rect 16497 16949 16531 16983
rect 18889 16949 18923 16983
rect 22385 16949 22419 16983
rect 23489 16949 23523 16983
rect 24317 16949 24351 16983
rect 25697 16949 25731 16983
rect 26433 16949 26467 16983
rect 6745 16745 6779 16779
rect 7297 16745 7331 16779
rect 14381 16745 14415 16779
rect 15761 16745 15795 16779
rect 18061 16745 18095 16779
rect 22201 16745 22235 16779
rect 27077 16745 27111 16779
rect 27721 16745 27755 16779
rect 28457 16745 28491 16779
rect 29745 16745 29779 16779
rect 30205 16745 30239 16779
rect 30389 16745 30423 16779
rect 13645 16677 13679 16711
rect 14289 16677 14323 16711
rect 15301 16677 15335 16711
rect 23673 16677 23707 16711
rect 27537 16677 27571 16711
rect 5365 16609 5399 16643
rect 7389 16609 7423 16643
rect 11161 16609 11195 16643
rect 11805 16609 11839 16643
rect 13921 16609 13955 16643
rect 16313 16609 16347 16643
rect 17325 16609 17359 16643
rect 18521 16609 18555 16643
rect 18705 16609 18739 16643
rect 18981 16609 19015 16643
rect 20821 16609 20855 16643
rect 23857 16609 23891 16643
rect 24409 16609 24443 16643
rect 26617 16609 26651 16643
rect 29653 16609 29687 16643
rect 30573 16609 30607 16643
rect 31033 16609 31067 16643
rect 1409 16541 1443 16575
rect 1685 16541 1719 16575
rect 5632 16541 5666 16575
rect 10425 16541 10459 16575
rect 11437 16541 11471 16575
rect 13553 16541 13587 16575
rect 14105 16541 14139 16575
rect 14565 16541 14599 16575
rect 14841 16541 14875 16575
rect 14933 16541 14967 16575
rect 15485 16541 15519 16575
rect 16129 16541 16163 16575
rect 16589 16541 16623 16575
rect 17233 16541 17267 16575
rect 18429 16541 18463 16575
rect 21088 16541 21122 16575
rect 22293 16541 22327 16575
rect 22560 16541 22594 16575
rect 24685 16541 24719 16575
rect 25329 16541 25363 16575
rect 25513 16541 25547 16575
rect 25697 16541 25731 16575
rect 26985 16541 27019 16575
rect 27261 16541 27295 16575
rect 28641 16541 28675 16575
rect 28917 16541 28951 16575
rect 29561 16541 29595 16575
rect 30021 16541 30055 16575
rect 30757 16541 30791 16575
rect 32781 16541 32815 16575
rect 34069 16541 34103 16575
rect 3157 16473 3191 16507
rect 4077 16473 4111 16507
rect 4905 16473 4939 16507
rect 7656 16473 7690 16507
rect 14749 16473 14783 16507
rect 23949 16473 23983 16507
rect 25605 16473 25639 16507
rect 34345 16473 34379 16507
rect 1593 16405 1627 16439
rect 5089 16405 5123 16439
rect 8769 16405 8803 16439
rect 15117 16405 15151 16439
rect 16221 16405 16255 16439
rect 16773 16405 16807 16439
rect 16957 16405 16991 16439
rect 19533 16405 19567 16439
rect 25881 16405 25915 16439
rect 26065 16405 26099 16439
rect 26433 16405 26467 16439
rect 26525 16405 26559 16439
rect 27445 16405 27479 16439
rect 28825 16405 28859 16439
rect 29101 16405 29135 16439
rect 29285 16405 29319 16439
rect 29929 16405 29963 16439
rect 32505 16405 32539 16439
rect 32597 16405 32631 16439
rect 32965 16405 32999 16439
rect 3617 16201 3651 16235
rect 4077 16201 4111 16235
rect 4445 16201 4479 16235
rect 8033 16201 8067 16235
rect 8493 16201 8527 16235
rect 11805 16201 11839 16235
rect 12265 16201 12299 16235
rect 12725 16201 12759 16235
rect 14565 16201 14599 16235
rect 15393 16201 15427 16235
rect 16313 16201 16347 16235
rect 17601 16201 17635 16235
rect 23029 16201 23063 16235
rect 27629 16201 27663 16235
rect 8401 16133 8435 16167
rect 12173 16133 12207 16167
rect 13360 16133 13394 16167
rect 15853 16133 15887 16167
rect 15945 16133 15979 16167
rect 18889 16133 18923 16167
rect 24869 16133 24903 16167
rect 24961 16133 24995 16167
rect 27261 16133 27295 16167
rect 29285 16133 29319 16167
rect 3433 16065 3467 16099
rect 3709 16065 3743 16099
rect 6377 16065 6411 16099
rect 6644 16065 6678 16099
rect 8861 16065 8895 16099
rect 8954 16065 8988 16099
rect 9137 16065 9171 16099
rect 9229 16065 9263 16099
rect 9367 16065 9401 16099
rect 9781 16065 9815 16099
rect 10885 16065 10919 16099
rect 11161 16065 11195 16099
rect 13093 16065 13127 16099
rect 14933 16065 14967 16099
rect 15577 16065 15611 16099
rect 15670 16065 15704 16099
rect 16042 16065 16076 16099
rect 16681 16065 16715 16099
rect 17325 16065 17359 16099
rect 18613 16065 18647 16099
rect 18761 16065 18795 16099
rect 18981 16065 19015 16099
rect 19119 16065 19153 16099
rect 19800 16065 19834 16099
rect 21833 16065 21867 16099
rect 21925 16065 21959 16099
rect 22109 16065 22143 16099
rect 22201 16065 22235 16099
rect 22477 16065 22511 16099
rect 22661 16065 22695 16099
rect 23305 16065 23339 16099
rect 23572 16065 23606 16099
rect 26525 16065 26559 16099
rect 26985 16065 27019 16099
rect 27078 16065 27112 16099
rect 27353 16065 27387 16099
rect 27450 16065 27484 16099
rect 28080 16065 28114 16099
rect 30941 16065 30975 16099
rect 31033 16065 31067 16099
rect 31401 16065 31435 16099
rect 31617 16065 31651 16099
rect 4537 15997 4571 16031
rect 4721 15997 4755 16031
rect 8677 15997 8711 16031
rect 12449 15997 12483 16031
rect 15025 15997 15059 16031
rect 15117 15997 15151 16031
rect 19533 15997 19567 16031
rect 27813 15997 27847 16031
rect 30113 15997 30147 16031
rect 30481 15997 30515 16031
rect 31125 15997 31159 16031
rect 32413 15997 32447 16031
rect 32689 15997 32723 16031
rect 9505 15929 9539 15963
rect 14473 15929 14507 15963
rect 19257 15929 19291 15963
rect 22385 15929 22419 15963
rect 24685 15929 24719 15963
rect 3893 15861 3927 15895
rect 7757 15861 7791 15895
rect 9689 15861 9723 15895
rect 11713 15861 11747 15895
rect 16221 15861 16255 15895
rect 19349 15861 19383 15895
rect 20913 15861 20947 15895
rect 22937 15861 22971 15895
rect 29193 15861 29227 15895
rect 30573 15861 30607 15895
rect 31493 15861 31527 15895
rect 31861 15861 31895 15895
rect 32137 15861 32171 15895
rect 34161 15861 34195 15895
rect 6837 15657 6871 15691
rect 7573 15657 7607 15691
rect 7665 15657 7699 15691
rect 18889 15657 18923 15691
rect 20085 15657 20119 15691
rect 22661 15657 22695 15691
rect 23857 15657 23891 15691
rect 24409 15657 24443 15691
rect 24685 15657 24719 15691
rect 26801 15657 26835 15691
rect 28457 15657 28491 15691
rect 30205 15657 30239 15691
rect 31769 15657 31803 15691
rect 5825 15589 5859 15623
rect 15393 15589 15427 15623
rect 19441 15589 19475 15623
rect 19625 15589 19659 15623
rect 22845 15589 22879 15623
rect 27813 15589 27847 15623
rect 27997 15589 28031 15623
rect 6285 15521 6319 15555
rect 7205 15521 7239 15555
rect 8585 15521 8619 15555
rect 9137 15521 9171 15555
rect 9413 15521 9447 15555
rect 13093 15521 13127 15555
rect 15945 15521 15979 15555
rect 16037 15521 16071 15555
rect 17325 15521 17359 15555
rect 17509 15521 17543 15555
rect 20545 15521 20579 15555
rect 20729 15521 20763 15555
rect 23949 15521 23983 15555
rect 26893 15521 26927 15555
rect 27169 15521 27203 15555
rect 28917 15521 28951 15555
rect 29101 15521 29135 15555
rect 2237 15453 2271 15487
rect 3801 15453 3835 15487
rect 5273 15453 5307 15487
rect 5549 15453 5583 15487
rect 5641 15453 5675 15487
rect 6469 15453 6503 15487
rect 7389 15453 7423 15487
rect 10885 15453 10919 15487
rect 10978 15453 11012 15487
rect 11161 15453 11195 15487
rect 11391 15453 11425 15487
rect 15669 15453 15703 15487
rect 15853 15453 15887 15487
rect 16221 15453 16255 15487
rect 19257 15453 19291 15487
rect 21281 15453 21315 15487
rect 25421 15453 25455 15487
rect 29561 15453 29595 15487
rect 30389 15453 30423 15487
rect 30656 15453 30690 15487
rect 33425 15453 33459 15487
rect 34529 15453 34563 15487
rect 2504 15385 2538 15419
rect 4068 15385 4102 15419
rect 5457 15385 5491 15419
rect 5917 15385 5951 15419
rect 6377 15385 6411 15419
rect 8309 15385 8343 15419
rect 9680 15385 9714 15419
rect 11253 15385 11287 15419
rect 12826 15385 12860 15419
rect 15485 15385 15519 15419
rect 16497 15385 16531 15419
rect 17776 15385 17810 15419
rect 20453 15385 20487 15419
rect 21548 15385 21582 15419
rect 24869 15385 24903 15419
rect 25688 15385 25722 15419
rect 28825 15385 28859 15419
rect 31953 15385 31987 15419
rect 32321 15385 32355 15419
rect 33057 15385 33091 15419
rect 34253 15385 34287 15419
rect 3617 15317 3651 15351
rect 5181 15317 5215 15351
rect 7021 15317 7055 15351
rect 7941 15317 7975 15351
rect 8401 15317 8435 15351
rect 9045 15317 9079 15351
rect 10793 15317 10827 15351
rect 11529 15317 11563 15351
rect 11713 15317 11747 15351
rect 13185 15317 13219 15351
rect 16405 15317 16439 15351
rect 19901 15317 19935 15351
rect 21005 15317 21039 15351
rect 24225 15317 24259 15351
rect 29285 15317 29319 15351
rect 32137 15317 32171 15351
rect 2881 15113 2915 15147
rect 3249 15113 3283 15147
rect 3709 15113 3743 15147
rect 4169 15113 4203 15147
rect 4629 15113 4663 15147
rect 8769 15113 8803 15147
rect 9965 15113 9999 15147
rect 10333 15113 10367 15147
rect 12173 15113 12207 15147
rect 13093 15113 13127 15147
rect 15485 15113 15519 15147
rect 17049 15113 17083 15147
rect 17969 15113 18003 15147
rect 18337 15113 18371 15147
rect 20453 15113 20487 15147
rect 21465 15113 21499 15147
rect 21833 15113 21867 15147
rect 22201 15113 22235 15147
rect 23581 15113 23615 15147
rect 23949 15113 23983 15147
rect 24317 15113 24351 15147
rect 26065 15113 26099 15147
rect 29745 15113 29779 15147
rect 30021 15113 30055 15147
rect 30573 15113 30607 15147
rect 32689 15113 32723 15147
rect 3341 15045 3375 15079
rect 4537 15045 4571 15079
rect 10425 15045 10459 15079
rect 11529 15045 11563 15079
rect 18429 15045 18463 15079
rect 20361 15045 20395 15079
rect 21189 15045 21223 15079
rect 29929 15045 29963 15079
rect 30481 15045 30515 15079
rect 31677 15045 31711 15079
rect 32321 15045 32355 15079
rect 32413 15045 32447 15079
rect 1409 14977 1443 15011
rect 1869 14977 1903 15011
rect 7389 14977 7423 15011
rect 7656 14977 7690 15011
rect 11805 14977 11839 15011
rect 12541 14977 12575 15011
rect 14372 14977 14406 15011
rect 16313 14977 16347 15011
rect 20821 14977 20855 15011
rect 20914 14977 20948 15011
rect 21097 14977 21131 15011
rect 21327 14977 21361 15011
rect 22293 14977 22327 15011
rect 23397 14977 23431 15011
rect 23765 14977 23799 15011
rect 24225 14977 24259 15011
rect 24685 14977 24719 15011
rect 24952 14977 24986 15011
rect 26157 14977 26191 15011
rect 26801 14977 26835 15011
rect 27241 14977 27275 15011
rect 28457 14977 28491 15011
rect 29101 14977 29135 15011
rect 29194 14977 29228 15011
rect 29377 14977 29411 15011
rect 29469 14977 29503 15011
rect 29607 14977 29641 15011
rect 30941 14977 30975 15011
rect 31217 14977 31251 15011
rect 31401 14977 31435 15011
rect 32137 14977 32171 15011
rect 32505 14977 32539 15011
rect 3525 14909 3559 14943
rect 4813 14909 4847 14943
rect 10517 14909 10551 14943
rect 10793 14909 10827 14943
rect 11621 14909 11655 14943
rect 12633 14909 12667 14943
rect 12817 14909 12851 14943
rect 14105 14909 14139 14943
rect 17141 14909 17175 14943
rect 17325 14909 17359 14943
rect 18613 14909 18647 14943
rect 20545 14909 20579 14943
rect 22477 14909 22511 14943
rect 26985 14909 27019 14943
rect 33241 14909 33275 14943
rect 33517 14909 33551 14943
rect 1593 14841 1627 14875
rect 1777 14841 1811 14875
rect 11989 14841 12023 14875
rect 17877 14841 17911 14875
rect 28641 14841 28675 14875
rect 30757 14841 30791 14875
rect 5089 14773 5123 14807
rect 6009 14773 6043 14807
rect 11253 14773 11287 14807
rect 11529 14773 11563 14807
rect 16497 14773 16531 14807
rect 16681 14773 16715 14807
rect 17601 14773 17635 14807
rect 19993 14773 20027 14807
rect 21557 14773 21591 14807
rect 22753 14773 22787 14807
rect 26341 14773 26375 14807
rect 26525 14773 26559 14807
rect 28365 14773 28399 14807
rect 28825 14773 28859 14807
rect 31033 14773 31067 14807
rect 31769 14773 31803 14807
rect 32781 14773 32815 14807
rect 34989 14773 35023 14807
rect 14657 14569 14691 14603
rect 15669 14569 15703 14603
rect 20821 14569 20855 14603
rect 21649 14569 21683 14603
rect 25237 14569 25271 14603
rect 26249 14569 26283 14603
rect 26985 14569 27019 14603
rect 27905 14569 27939 14603
rect 29193 14569 29227 14603
rect 29745 14569 29779 14603
rect 30941 14569 30975 14603
rect 33793 14569 33827 14603
rect 33977 14569 34011 14603
rect 24225 14501 24259 14535
rect 28549 14501 28583 14535
rect 29561 14501 29595 14535
rect 10425 14433 10459 14467
rect 12357 14433 12391 14467
rect 12541 14433 12575 14467
rect 15117 14433 15151 14467
rect 15301 14433 15335 14467
rect 17049 14433 17083 14467
rect 24961 14433 24995 14467
rect 25697 14433 25731 14467
rect 25881 14433 25915 14467
rect 27445 14433 27479 14467
rect 27629 14433 27663 14467
rect 30481 14433 30515 14467
rect 30573 14433 30607 14467
rect 31033 14433 31067 14467
rect 5365 14365 5399 14399
rect 10793 14365 10827 14399
rect 10886 14365 10920 14399
rect 11299 14365 11333 14399
rect 12081 14365 12115 14399
rect 15025 14365 15059 14399
rect 16782 14365 16816 14399
rect 19441 14365 19475 14399
rect 19708 14365 19742 14399
rect 22845 14365 22879 14399
rect 24777 14365 24811 14399
rect 25605 14365 25639 14399
rect 27353 14365 27387 14399
rect 27997 14365 28031 14399
rect 28365 14365 28399 14399
rect 28647 14365 28681 14399
rect 29009 14365 29043 14399
rect 30389 14365 30423 14399
rect 34161 14365 34195 14399
rect 34437 14365 34471 14399
rect 5632 14297 5666 14331
rect 10241 14297 10275 14331
rect 11069 14297 11103 14331
rect 11161 14297 11195 14331
rect 12817 14297 12851 14331
rect 15577 14297 15611 14331
rect 23112 14297 23146 14331
rect 28181 14297 28215 14331
rect 28273 14297 28307 14331
rect 34345 14297 34379 14331
rect 6745 14229 6779 14263
rect 9873 14229 9907 14263
rect 10333 14229 10367 14263
rect 11437 14229 11471 14263
rect 12725 14229 12759 14263
rect 21741 14229 21775 14263
rect 24409 14229 24443 14263
rect 24869 14229 24903 14263
rect 26157 14229 26191 14263
rect 28825 14229 28859 14263
rect 30021 14229 30055 14263
rect 4905 14025 4939 14059
rect 6377 14025 6411 14059
rect 6745 14025 6779 14059
rect 7757 14025 7791 14059
rect 8125 14025 8159 14059
rect 10701 14025 10735 14059
rect 11989 14025 12023 14059
rect 14473 14025 14507 14059
rect 21281 14025 21315 14059
rect 23857 14025 23891 14059
rect 25237 14025 25271 14059
rect 27077 14025 27111 14059
rect 27997 14025 28031 14059
rect 29561 14025 29595 14059
rect 31125 14025 31159 14059
rect 4537 13957 4571 13991
rect 5089 13957 5123 13991
rect 7481 13957 7515 13991
rect 7849 13957 7883 13991
rect 9588 13957 9622 13991
rect 10793 13957 10827 13991
rect 22652 13957 22686 13991
rect 24225 13957 24259 13991
rect 24961 13957 24995 13991
rect 25973 13957 26007 13991
rect 26341 13957 26375 13991
rect 28448 13957 28482 13991
rect 3433 13889 3467 13923
rect 4353 13889 4387 13923
rect 4629 13889 4663 13923
rect 4721 13889 4755 13923
rect 7205 13889 7239 13923
rect 7389 13889 7423 13923
rect 7573 13889 7607 13923
rect 9321 13889 9355 13923
rect 11897 13889 11931 13923
rect 12357 13889 12391 13923
rect 12624 13889 12658 13923
rect 13829 13889 13863 13923
rect 13922 13889 13956 13923
rect 14105 13889 14139 13923
rect 14197 13889 14231 13923
rect 14335 13889 14369 13923
rect 16773 13889 16807 13923
rect 17040 13889 17074 13923
rect 18337 13889 18371 13923
rect 18604 13889 18638 13923
rect 21465 13889 21499 13923
rect 22109 13889 22143 13923
rect 24685 13889 24719 13923
rect 24869 13889 24903 13923
rect 25053 13889 25087 13923
rect 25605 13889 25639 13923
rect 28181 13889 28215 13923
rect 30012 13889 30046 13923
rect 6837 13821 6871 13855
rect 7021 13821 7055 13855
rect 12173 13821 12207 13855
rect 14657 13821 14691 13855
rect 14841 13821 14875 13855
rect 22385 13821 22419 13855
rect 24317 13821 24351 13855
rect 24409 13821 24443 13855
rect 26433 13821 26467 13855
rect 26617 13821 26651 13855
rect 29745 13821 29779 13855
rect 21649 13753 21683 13787
rect 23765 13753 23799 13787
rect 25421 13753 25455 13787
rect 3617 13685 3651 13719
rect 11529 13685 11563 13719
rect 13737 13685 13771 13719
rect 18153 13685 18187 13719
rect 19717 13685 19751 13719
rect 21925 13685 21959 13719
rect 22201 13685 22235 13719
rect 25697 13685 25731 13719
rect 3617 13481 3651 13515
rect 6929 13481 6963 13515
rect 7297 13481 7331 13515
rect 11897 13481 11931 13515
rect 12265 13481 12299 13515
rect 12817 13481 12851 13515
rect 14933 13481 14967 13515
rect 17325 13481 17359 13515
rect 19257 13481 19291 13515
rect 23765 13481 23799 13515
rect 24501 13481 24535 13515
rect 27261 13481 27295 13515
rect 27537 13481 27571 13515
rect 28273 13481 28307 13515
rect 28457 13481 28491 13515
rect 29285 13481 29319 13515
rect 13645 13413 13679 13447
rect 18889 13413 18923 13447
rect 21833 13413 21867 13447
rect 5549 13345 5583 13379
rect 9505 13345 9539 13379
rect 9781 13345 9815 13379
rect 12357 13345 12391 13379
rect 13369 13345 13403 13379
rect 14565 13345 14599 13379
rect 14749 13345 14783 13379
rect 15117 13345 15151 13379
rect 17877 13345 17911 13379
rect 18153 13345 18187 13379
rect 19809 13345 19843 13379
rect 20085 13345 20119 13379
rect 22753 13345 22787 13379
rect 24961 13345 24995 13379
rect 27997 13345 28031 13379
rect 28917 13345 28951 13379
rect 29009 13345 29043 13379
rect 2237 13277 2271 13311
rect 3801 13277 3835 13311
rect 7389 13277 7423 13311
rect 10517 13277 10551 13311
rect 10784 13277 10818 13311
rect 12265 13277 12299 13311
rect 13185 13277 13219 13311
rect 16589 13277 16623 13311
rect 17693 13277 17727 13311
rect 20453 13277 20487 13311
rect 26433 13277 26467 13311
rect 26526 13277 26560 13311
rect 26709 13277 26743 13311
rect 26939 13277 26973 13311
rect 27353 13277 27387 13311
rect 27721 13277 27755 13311
rect 28825 13277 28859 13311
rect 2504 13209 2538 13243
rect 4068 13209 4102 13243
rect 5816 13209 5850 13243
rect 7656 13209 7690 13243
rect 9413 13209 9447 13243
rect 13277 13209 13311 13243
rect 15384 13209 15418 13243
rect 20720 13209 20754 13243
rect 21925 13209 21959 13243
rect 25228 13209 25262 13243
rect 26801 13209 26835 13243
rect 5181 13141 5215 13175
rect 8769 13141 8803 13175
rect 8953 13141 8987 13175
rect 9321 13141 9355 13175
rect 12633 13141 12667 13175
rect 14105 13141 14139 13175
rect 14473 13141 14507 13175
rect 16497 13141 16531 13175
rect 16773 13141 16807 13175
rect 17785 13141 17819 13175
rect 19625 13141 19659 13175
rect 19717 13141 19751 13175
rect 22937 13141 22971 13175
rect 23949 13141 23983 13175
rect 26341 13141 26375 13175
rect 27077 13141 27111 13175
rect 1593 12937 1627 12971
rect 2973 12937 3007 12971
rect 3985 12937 4019 12971
rect 4353 12937 4387 12971
rect 6377 12937 6411 12971
rect 6745 12937 6779 12971
rect 9229 12937 9263 12971
rect 15117 12937 15151 12971
rect 15669 12937 15703 12971
rect 16037 12937 16071 12971
rect 16129 12937 16163 12971
rect 17785 12937 17819 12971
rect 25513 12937 25547 12971
rect 25881 12937 25915 12971
rect 26617 12937 26651 12971
rect 28365 12937 28399 12971
rect 3433 12869 3467 12903
rect 9413 12869 9447 12903
rect 9597 12869 9631 12903
rect 14004 12869 14038 12903
rect 17049 12869 17083 12903
rect 21281 12869 21315 12903
rect 21373 12869 21407 12903
rect 25145 12869 25179 12903
rect 28457 12869 28491 12903
rect 28825 12869 28859 12903
rect 1409 12801 1443 12835
rect 1685 12801 1719 12835
rect 3341 12801 3375 12835
rect 4445 12801 4479 12835
rect 6837 12801 6871 12835
rect 8677 12801 8711 12835
rect 8769 12801 8803 12835
rect 8953 12801 8987 12835
rect 9045 12801 9079 12835
rect 16865 12801 16899 12835
rect 17141 12801 17175 12835
rect 17233 12801 17267 12835
rect 17509 12801 17543 12835
rect 18061 12801 18095 12835
rect 18154 12801 18188 12835
rect 18337 12801 18371 12835
rect 18429 12801 18463 12835
rect 18526 12801 18560 12835
rect 18797 12801 18831 12835
rect 18981 12801 19015 12835
rect 19073 12801 19107 12835
rect 19165 12801 19199 12835
rect 19349 12801 19383 12835
rect 20913 12801 20947 12835
rect 21097 12801 21131 12835
rect 21465 12801 21499 12835
rect 21925 12801 21959 12835
rect 23213 12801 23247 12835
rect 23306 12801 23340 12835
rect 23489 12801 23523 12835
rect 23581 12801 23615 12835
rect 23678 12801 23712 12835
rect 24501 12801 24535 12835
rect 26525 12801 26559 12835
rect 26985 12801 27019 12835
rect 27252 12801 27286 12835
rect 32137 12801 32171 12835
rect 34529 12801 34563 12835
rect 3617 12733 3651 12767
rect 4629 12733 4663 12767
rect 7021 12733 7055 12767
rect 7205 12733 7239 12767
rect 13737 12733 13771 12767
rect 16313 12733 16347 12767
rect 19625 12733 19659 12767
rect 22201 12733 22235 12767
rect 24777 12733 24811 12767
rect 25973 12733 26007 12767
rect 26157 12733 26191 12767
rect 32413 12733 32447 12767
rect 34805 12733 34839 12767
rect 7389 12665 7423 12699
rect 16773 12665 16807 12699
rect 17417 12665 17451 12699
rect 18705 12665 18739 12699
rect 19809 12665 19843 12699
rect 21649 12665 21683 12699
rect 23029 12665 23063 12699
rect 23857 12665 23891 12699
rect 26341 12665 26375 12699
rect 3893 12597 3927 12631
rect 19533 12597 19567 12631
rect 19993 12597 20027 12631
rect 22845 12597 22879 12631
rect 24869 12597 24903 12631
rect 28641 12597 28675 12631
rect 33885 12597 33919 12631
rect 13001 12393 13035 12427
rect 13369 12393 13403 12427
rect 21189 12393 21223 12427
rect 21833 12393 21867 12427
rect 24225 12393 24259 12427
rect 25145 12393 25179 12427
rect 25789 12393 25823 12427
rect 26617 12393 26651 12427
rect 26801 12393 26835 12427
rect 27261 12393 27295 12427
rect 32229 12393 32263 12427
rect 33241 12393 33275 12427
rect 18705 12325 18739 12359
rect 19533 12325 19567 12359
rect 21465 12325 21499 12359
rect 22661 12325 22695 12359
rect 24501 12325 24535 12359
rect 26893 12325 26927 12359
rect 32873 12325 32907 12359
rect 7665 12257 7699 12291
rect 8677 12257 8711 12291
rect 13185 12257 13219 12291
rect 19349 12257 19383 12291
rect 19809 12257 19843 12291
rect 22385 12257 22419 12291
rect 26525 12257 26559 12291
rect 27813 12257 27847 12291
rect 28089 12257 28123 12291
rect 29837 12257 29871 12291
rect 8033 12189 8067 12223
rect 8217 12189 8251 12223
rect 8401 12189 8435 12223
rect 8953 12189 8987 12223
rect 12449 12189 12483 12223
rect 12633 12189 12667 12223
rect 12817 12189 12851 12223
rect 18889 12189 18923 12223
rect 21649 12189 21683 12223
rect 22201 12189 22235 12223
rect 22845 12189 22879 12223
rect 24685 12189 24719 12223
rect 25053 12189 25087 12223
rect 26433 12189 26467 12223
rect 27629 12189 27663 12223
rect 31677 12189 31711 12223
rect 31953 12189 31987 12223
rect 32045 12189 32079 12223
rect 6009 12121 6043 12155
rect 6745 12121 6779 12155
rect 8309 12121 8343 12155
rect 12725 12121 12759 12155
rect 20076 12121 20110 12155
rect 23112 12121 23146 12155
rect 25421 12121 25455 12155
rect 30104 12121 30138 12155
rect 31861 12121 31895 12155
rect 33149 12121 33183 12155
rect 7021 12053 7055 12087
rect 7389 12053 7423 12087
rect 7481 12053 7515 12087
rect 7941 12053 7975 12087
rect 8585 12053 8619 12087
rect 22293 12053 22327 12087
rect 24869 12053 24903 12087
rect 25513 12053 25547 12087
rect 25881 12053 25915 12087
rect 27721 12053 27755 12087
rect 28273 12053 28307 12087
rect 31217 12053 31251 12087
rect 11345 11849 11379 11883
rect 13185 11849 13219 11883
rect 14105 11849 14139 11883
rect 17049 11849 17083 11883
rect 18981 11849 19015 11883
rect 20361 11849 20395 11883
rect 20729 11849 20763 11883
rect 20821 11849 20855 11883
rect 23489 11849 23523 11883
rect 23857 11849 23891 11883
rect 25605 11849 25639 11883
rect 26617 11849 26651 11883
rect 27261 11849 27295 11883
rect 30113 11849 30147 11883
rect 31401 11849 31435 11883
rect 31493 11849 31527 11883
rect 15301 11781 15335 11815
rect 26157 11781 26191 11815
rect 27629 11781 27663 11815
rect 29561 11781 29595 11815
rect 2881 11713 2915 11747
rect 3148 11713 3182 11747
rect 4353 11713 4387 11747
rect 4620 11713 4654 11747
rect 6561 11713 6595 11747
rect 7021 11713 7055 11747
rect 7288 11713 7322 11747
rect 8493 11713 8527 11747
rect 8760 11713 8794 11747
rect 9965 11713 9999 11747
rect 10232 11713 10266 11747
rect 12072 11713 12106 11747
rect 14657 11713 14691 11747
rect 14749 11713 14783 11747
rect 14933 11713 14967 11747
rect 15025 11713 15059 11747
rect 16129 11713 16163 11747
rect 17141 11713 17175 11747
rect 17601 11713 17635 11747
rect 17868 11713 17902 11747
rect 22100 11713 22134 11747
rect 24317 11713 24351 11747
rect 25053 11713 25087 11747
rect 25421 11713 25455 11747
rect 25973 11713 26007 11747
rect 26249 11713 26283 11747
rect 26341 11713 26375 11747
rect 27077 11713 27111 11747
rect 27721 11713 27755 11747
rect 29110 11713 29144 11747
rect 30481 11713 30515 11747
rect 30573 11713 30607 11747
rect 30941 11713 30975 11747
rect 31033 11713 31067 11747
rect 31217 11713 31251 11747
rect 34529 11713 34563 11747
rect 11805 11645 11839 11679
rect 17233 11645 17267 11679
rect 20269 11645 20303 11679
rect 21005 11645 21039 11679
rect 21833 11645 21867 11679
rect 23949 11645 23983 11679
rect 24041 11645 24075 11679
rect 25789 11645 25823 11679
rect 27353 11645 27387 11679
rect 29377 11645 29411 11679
rect 30665 11645 30699 11679
rect 34805 11645 34839 11679
rect 15945 11577 15979 11611
rect 23213 11577 23247 11611
rect 24501 11577 24535 11611
rect 24685 11577 24719 11611
rect 24869 11577 24903 11611
rect 27997 11577 28031 11611
rect 4261 11509 4295 11543
rect 5733 11509 5767 11543
rect 8401 11509 8435 11543
rect 9873 11509 9907 11543
rect 15209 11509 15243 11543
rect 16681 11509 16715 11543
rect 25237 11509 25271 11543
rect 26525 11509 26559 11543
rect 29653 11509 29687 11543
rect 29837 11509 29871 11543
rect 3801 11305 3835 11339
rect 4905 11305 4939 11339
rect 7481 11305 7515 11339
rect 7665 11305 7699 11339
rect 9413 11305 9447 11339
rect 10977 11305 11011 11339
rect 12357 11305 12391 11339
rect 13921 11305 13955 11339
rect 14473 11305 14507 11339
rect 17325 11305 17359 11339
rect 17601 11305 17635 11339
rect 18061 11305 18095 11339
rect 18981 11305 19015 11339
rect 21189 11305 21223 11339
rect 21465 11305 21499 11339
rect 22201 11305 22235 11339
rect 25789 11305 25823 11339
rect 26341 11305 26375 11339
rect 26709 11305 26743 11339
rect 26801 11305 26835 11339
rect 29101 11305 29135 11339
rect 30573 11305 30607 11339
rect 6009 11237 6043 11271
rect 26617 11237 26651 11271
rect 27445 11237 27479 11271
rect 29193 11237 29227 11271
rect 2973 11169 3007 11203
rect 3341 11169 3375 11203
rect 3617 11169 3651 11203
rect 4261 11169 4295 11203
rect 4445 11169 4479 11203
rect 5549 11169 5583 11203
rect 5733 11169 5767 11203
rect 8125 11169 8159 11203
rect 8217 11169 8251 11203
rect 8493 11169 8527 11203
rect 9873 11169 9907 11203
rect 10057 11169 10091 11203
rect 11621 11169 11655 11203
rect 11897 11169 11931 11203
rect 13001 11169 13035 11203
rect 13277 11169 13311 11203
rect 18521 11169 18555 11203
rect 18705 11169 18739 11203
rect 22753 11169 22787 11203
rect 24409 11169 24443 11203
rect 26249 11169 26283 11203
rect 27813 11169 27847 11203
rect 28549 11169 28583 11203
rect 30665 11169 30699 11203
rect 1409 11101 1443 11135
rect 1685 11101 1719 11135
rect 4169 11101 4203 11135
rect 4813 11101 4847 11135
rect 5273 11101 5307 11135
rect 6101 11101 6135 11135
rect 8033 11101 8067 11135
rect 9781 11101 9815 11135
rect 10241 11101 10275 11135
rect 10425 11101 10459 11135
rect 10517 11101 10551 11135
rect 10701 11101 10735 11135
rect 10793 11101 10827 11135
rect 11345 11101 11379 11135
rect 12725 11101 12759 11135
rect 13369 11101 13403 11135
rect 13553 11101 13587 11135
rect 13737 11101 13771 11135
rect 14197 11101 14231 11135
rect 15853 11101 15887 11135
rect 15945 11101 15979 11135
rect 16212 11101 16246 11135
rect 18429 11101 18463 11135
rect 19809 11101 19843 11135
rect 21373 11101 21407 11135
rect 22569 11101 22603 11135
rect 27077 11101 27111 11135
rect 27261 11101 27295 11135
rect 27905 11101 27939 11135
rect 28733 11101 28767 11135
rect 29561 11101 29595 11135
rect 29837 11101 29871 11135
rect 34161 11101 34195 11135
rect 34437 11101 34471 11135
rect 3157 11033 3191 11067
rect 5365 11033 5399 11067
rect 6368 11033 6402 11067
rect 11437 11033 11471 11067
rect 12817 11033 12851 11067
rect 13645 11033 13679 11067
rect 15608 11033 15642 11067
rect 19625 11033 19659 11067
rect 22109 11033 22143 11067
rect 22661 11033 22695 11067
rect 24676 11033 24710 11067
rect 27629 11033 27663 11067
rect 28641 11033 28675 11067
rect 34345 11033 34379 11067
rect 1593 10965 1627 10999
rect 19993 10965 20027 10999
rect 25881 10965 25915 10999
rect 26985 10965 27019 10999
rect 28089 10965 28123 10999
rect 33977 10965 34011 10999
rect 3341 10761 3375 10795
rect 3801 10761 3835 10795
rect 4721 10761 4755 10795
rect 5733 10761 5767 10795
rect 10241 10761 10275 10795
rect 10885 10761 10919 10795
rect 11161 10761 11195 10795
rect 13829 10761 13863 10795
rect 14013 10761 14047 10795
rect 15761 10761 15795 10795
rect 16129 10761 16163 10795
rect 18797 10761 18831 10795
rect 20637 10761 20671 10795
rect 22477 10761 22511 10795
rect 24961 10761 24995 10795
rect 25421 10761 25455 10795
rect 26985 10761 27019 10795
rect 29929 10761 29963 10795
rect 30389 10761 30423 10795
rect 34989 10761 35023 10795
rect 3004 10693 3038 10727
rect 4445 10693 4479 10727
rect 5273 10693 5307 10727
rect 14657 10693 14691 10727
rect 14749 10693 14783 10727
rect 15485 10693 15519 10727
rect 17141 10693 17175 10727
rect 21465 10693 21499 10727
rect 25329 10693 25363 10727
rect 29570 10693 29604 10727
rect 33517 10693 33551 10727
rect 3249 10625 3283 10659
rect 3709 10625 3743 10659
rect 4169 10625 4203 10659
rect 4353 10625 4387 10659
rect 4537 10625 4571 10659
rect 4905 10625 4939 10659
rect 4998 10625 5032 10659
rect 5181 10625 5215 10659
rect 5411 10625 5445 10659
rect 12633 10625 12667 10659
rect 14197 10625 14231 10659
rect 17049 10625 17083 10659
rect 17785 10625 17819 10659
rect 18153 10625 18187 10659
rect 19921 10625 19955 10659
rect 20177 10625 20211 10659
rect 21281 10625 21315 10659
rect 21373 10625 21407 10659
rect 21649 10625 21683 10659
rect 21833 10625 21867 10659
rect 22201 10625 22235 10659
rect 22661 10625 22695 10659
rect 28098 10625 28132 10659
rect 28365 10625 28399 10659
rect 30297 10625 30331 10659
rect 3985 10557 4019 10591
rect 12909 10557 12943 10591
rect 16221 10557 16255 10591
rect 16405 10557 16439 10591
rect 17233 10557 17267 10591
rect 17877 10557 17911 10591
rect 18245 10557 18279 10591
rect 20729 10557 20763 10591
rect 20913 10557 20947 10591
rect 25513 10557 25547 10591
rect 25789 10557 25823 10591
rect 29837 10557 29871 10591
rect 30481 10557 30515 10591
rect 33241 10557 33275 10591
rect 14473 10489 14507 10523
rect 17601 10489 17635 10523
rect 20269 10489 20303 10523
rect 1869 10421 1903 10455
rect 5549 10421 5583 10455
rect 5917 10421 5951 10455
rect 11253 10421 11287 10455
rect 12817 10421 12851 10455
rect 16681 10421 16715 10455
rect 21097 10421 21131 10455
rect 22017 10421 22051 10455
rect 28457 10421 28491 10455
rect 3249 10217 3283 10251
rect 3617 10217 3651 10251
rect 4905 10217 4939 10251
rect 6745 10217 6779 10251
rect 8677 10217 8711 10251
rect 9873 10217 9907 10251
rect 11621 10217 11655 10251
rect 13921 10217 13955 10251
rect 17141 10217 17175 10251
rect 22937 10217 22971 10251
rect 23489 10217 23523 10251
rect 24593 10217 24627 10251
rect 27445 10217 27479 10251
rect 27721 10217 27755 10251
rect 27905 10217 27939 10251
rect 28089 10217 28123 10251
rect 28365 10217 28399 10251
rect 4721 10149 4755 10183
rect 5273 10149 5307 10183
rect 8309 10149 8343 10183
rect 17877 10149 17911 10183
rect 18797 10149 18831 10183
rect 4445 10081 4479 10115
rect 10885 10081 10919 10115
rect 11345 10081 11379 10115
rect 12173 10081 12207 10115
rect 12265 10081 12299 10115
rect 12541 10081 12575 10115
rect 14565 10081 14599 10115
rect 14749 10081 14783 10115
rect 15761 10081 15795 10115
rect 18889 10081 18923 10115
rect 20361 10081 20395 10115
rect 23121 10081 23155 10115
rect 26801 10081 26835 10115
rect 30113 10081 30147 10115
rect 4169 10013 4203 10047
rect 5089 10013 5123 10047
rect 5365 10013 5399 10047
rect 6101 10013 6135 10047
rect 6469 10013 6503 10047
rect 7665 10013 7699 10047
rect 7813 10013 7847 10047
rect 8171 10013 8205 10047
rect 9321 10013 9355 10047
rect 10236 10013 10270 10047
rect 10425 10013 10459 10047
rect 10553 10013 10587 10047
rect 10701 10013 10735 10047
rect 11161 10013 11195 10047
rect 14473 10013 14507 10047
rect 16028 10013 16062 10047
rect 17233 10013 17267 10047
rect 17417 10013 17451 10047
rect 17601 10013 17635 10047
rect 18429 10013 18463 10047
rect 22753 10013 22787 10047
rect 22937 10013 22971 10047
rect 23029 10013 23063 10047
rect 23213 10013 23247 10047
rect 23305 10013 23339 10047
rect 23489 10013 23523 10047
rect 23581 10013 23615 10047
rect 23765 10013 23799 10047
rect 24409 10013 24443 10047
rect 24593 10013 24627 10047
rect 27077 10013 27111 10047
rect 27629 10013 27663 10047
rect 28820 10013 28854 10047
rect 29009 10013 29043 10047
rect 29192 10013 29226 10047
rect 29285 10013 29319 10047
rect 29653 10013 29687 10047
rect 31033 10013 31067 10047
rect 6285 9945 6319 9979
rect 6377 9945 6411 9979
rect 7941 9945 7975 9979
rect 8033 9945 8067 9979
rect 8493 9945 8527 9979
rect 10313 9945 10347 9979
rect 12081 9945 12115 9979
rect 12808 9945 12842 9979
rect 17505 9945 17539 9979
rect 20628 9945 20662 9979
rect 28917 9945 28951 9979
rect 30297 9945 30331 9979
rect 31217 9945 31251 9979
rect 32045 9945 32079 9979
rect 3801 9877 3835 9911
rect 4261 9877 4295 9911
rect 5549 9877 5583 9911
rect 6653 9877 6687 9911
rect 9505 9877 9539 9911
rect 10057 9877 10091 9911
rect 11713 9877 11747 9911
rect 14105 9877 14139 9911
rect 17785 9877 17819 9911
rect 18245 9877 18279 9911
rect 18521 9877 18555 9911
rect 21741 9877 21775 9911
rect 23673 9877 23707 9911
rect 26985 9877 27019 9911
rect 28457 9877 28491 9911
rect 28641 9877 28675 9911
rect 29745 9877 29779 9911
rect 30481 9877 30515 9911
rect 4353 9673 4387 9707
rect 8217 9673 8251 9707
rect 9781 9673 9815 9707
rect 13001 9673 13035 9707
rect 14013 9673 14047 9707
rect 20637 9673 20671 9707
rect 21005 9673 21039 9707
rect 25697 9673 25731 9707
rect 26709 9673 26743 9707
rect 28457 9673 28491 9707
rect 31125 9673 31159 9707
rect 3648 9605 3682 9639
rect 4905 9605 4939 9639
rect 5825 9605 5859 9639
rect 11866 9605 11900 9639
rect 24225 9605 24259 9639
rect 25237 9605 25271 9639
rect 25513 9605 25547 9639
rect 30297 9605 30331 9639
rect 4169 9537 4203 9571
rect 6653 9537 6687 9571
rect 6837 9537 6871 9571
rect 7104 9537 7138 9571
rect 8668 9537 8702 9571
rect 11078 9537 11112 9571
rect 14841 9537 14875 9571
rect 17417 9537 17451 9571
rect 17684 9537 17718 9571
rect 20085 9537 20119 9571
rect 20453 9537 20487 9571
rect 22937 9537 22971 9571
rect 23213 9537 23247 9571
rect 24041 9537 24075 9571
rect 24133 9537 24167 9571
rect 24317 9537 24351 9571
rect 24409 9537 24443 9571
rect 24593 9537 24627 9571
rect 24869 9537 24903 9571
rect 25053 9537 25087 9571
rect 25145 9537 25179 9571
rect 25329 9537 25363 9571
rect 25421 9537 25455 9571
rect 25605 9537 25639 9571
rect 26525 9537 26559 9571
rect 27077 9537 27111 9571
rect 27537 9537 27571 9571
rect 28181 9537 28215 9571
rect 29581 9537 29615 9571
rect 29837 9537 29871 9571
rect 34069 9537 34103 9571
rect 34253 9537 34287 9571
rect 34345 9537 34379 9571
rect 3893 9469 3927 9503
rect 4997 9469 5031 9503
rect 5089 9469 5123 9503
rect 5917 9469 5951 9503
rect 6101 9469 6135 9503
rect 8401 9469 8435 9503
rect 11345 9469 11379 9503
rect 11621 9469 11655 9503
rect 14933 9469 14967 9503
rect 16773 9469 16807 9503
rect 21097 9469 21131 9503
rect 21281 9469 21315 9503
rect 21833 9469 21867 9503
rect 28365 9469 28399 9503
rect 30389 9469 30423 9503
rect 30481 9469 30515 9503
rect 30757 9469 30791 9503
rect 4537 9401 4571 9435
rect 6469 9401 6503 9435
rect 18797 9401 18831 9435
rect 23213 9401 23247 9435
rect 24685 9401 24719 9435
rect 24869 9401 24903 9435
rect 26341 9401 26375 9435
rect 27721 9401 27755 9435
rect 29929 9401 29963 9435
rect 2513 9333 2547 9367
rect 3985 9333 4019 9367
rect 5457 9333 5491 9367
rect 9965 9333 9999 9367
rect 14933 9333 14967 9367
rect 15209 9333 15243 9367
rect 21465 9333 21499 9367
rect 23489 9333 23523 9367
rect 23857 9333 23891 9367
rect 27169 9333 27203 9367
rect 27997 9333 28031 9367
rect 33885 9333 33919 9367
rect 1593 9129 1627 9163
rect 5181 9129 5215 9163
rect 6653 9129 6687 9163
rect 7389 9129 7423 9163
rect 8953 9129 8987 9163
rect 10057 9129 10091 9163
rect 10333 9129 10367 9163
rect 11161 9129 11195 9163
rect 13645 9129 13679 9163
rect 14933 9129 14967 9163
rect 17785 9129 17819 9163
rect 23029 9129 23063 9163
rect 25237 9129 25271 9163
rect 28549 9129 28583 9163
rect 34529 9129 34563 9163
rect 8309 9061 8343 9095
rect 20637 9061 20671 9095
rect 24409 9061 24443 9095
rect 27077 9061 27111 9095
rect 28825 9061 28859 9095
rect 29561 9061 29595 9095
rect 8033 8993 8067 9027
rect 9597 8993 9631 9027
rect 10517 8993 10551 9027
rect 13461 8993 13495 9027
rect 18337 8993 18371 9027
rect 18613 8993 18647 9027
rect 21189 8993 21223 9027
rect 21281 8993 21315 9027
rect 21833 8993 21867 9027
rect 21925 8993 21959 9027
rect 22569 8993 22603 9027
rect 25697 8993 25731 9027
rect 27629 8993 27663 9027
rect 27813 8993 27847 9027
rect 33057 8993 33091 9027
rect 1409 8925 1443 8959
rect 1685 8925 1719 8959
rect 3801 8925 3835 8959
rect 4068 8925 4102 8959
rect 5273 8925 5307 8959
rect 5540 8925 5574 8959
rect 6837 8925 6871 8959
rect 7757 8925 7791 8959
rect 9321 8925 9355 8959
rect 9965 8925 9999 8959
rect 10057 8925 10091 8959
rect 10793 8925 10827 8959
rect 12725 8925 12759 8959
rect 13001 8925 13035 8959
rect 13093 8925 13127 8959
rect 14289 8925 14323 8959
rect 14437 8925 14471 8959
rect 14657 8925 14691 8959
rect 14793 8925 14827 8959
rect 15117 8925 15151 8959
rect 18245 8925 18279 8959
rect 19257 8925 19291 8959
rect 21097 8925 21131 8959
rect 21557 8925 21591 8959
rect 21741 8925 21775 8959
rect 22109 8925 22143 8959
rect 22844 8925 22878 8959
rect 22937 8925 22971 8959
rect 24623 8925 24657 8959
rect 24770 8925 24804 8959
rect 27537 8925 27571 8959
rect 27997 8925 28031 8959
rect 28365 8925 28399 8959
rect 28641 8925 28675 8959
rect 32781 8925 32815 8959
rect 10701 8857 10735 8891
rect 12909 8857 12943 8891
rect 14565 8857 14599 8891
rect 15301 8857 15335 8891
rect 19524 8857 19558 8891
rect 24869 8857 24903 8891
rect 25053 8857 25087 8891
rect 25964 8857 25998 8891
rect 28181 8857 28215 8891
rect 28273 8857 28307 8891
rect 29009 8857 29043 8891
rect 29193 8857 29227 8891
rect 7849 8789 7883 8823
rect 9413 8789 9447 8823
rect 9873 8789 9907 8823
rect 11253 8789 11287 8823
rect 13277 8789 13311 8823
rect 18153 8789 18187 8823
rect 20729 8789 20763 8823
rect 22293 8789 22327 8823
rect 22477 8789 22511 8823
rect 27169 8789 27203 8823
rect 4445 8585 4479 8619
rect 4629 8585 4663 8619
rect 10425 8585 10459 8619
rect 10793 8585 10827 8619
rect 15025 8585 15059 8619
rect 16497 8585 16531 8619
rect 17141 8585 17175 8619
rect 17785 8585 17819 8619
rect 18981 8585 19015 8619
rect 21097 8585 21131 8619
rect 21925 8585 21959 8619
rect 22753 8585 22787 8619
rect 22845 8585 22879 8619
rect 23121 8585 23155 8619
rect 28457 8585 28491 8619
rect 6469 8517 6503 8551
rect 7481 8517 7515 8551
rect 10057 8517 10091 8551
rect 10517 8517 10551 8551
rect 18797 8517 18831 8551
rect 19993 8517 20027 8551
rect 20821 8517 20855 8551
rect 21373 8517 21407 8551
rect 27252 8517 27286 8551
rect 28641 8517 28675 8551
rect 34805 8517 34839 8551
rect 7205 8449 7239 8483
rect 9873 8449 9907 8483
rect 10149 8449 10183 8483
rect 10241 8449 10275 8483
rect 12072 8449 12106 8483
rect 13912 8449 13946 8483
rect 15117 8449 15151 8483
rect 15384 8449 15418 8483
rect 17049 8449 17083 8483
rect 17877 8449 17911 8483
rect 18061 8449 18095 8483
rect 18153 8449 18187 8483
rect 18245 8449 18279 8483
rect 18429 8449 18463 8483
rect 20453 8449 20487 8483
rect 20601 8449 20635 8483
rect 20729 8449 20763 8483
rect 20959 8449 20993 8483
rect 23029 8449 23063 8483
rect 23213 8449 23247 8483
rect 23489 8449 23523 8483
rect 26985 8449 27019 8483
rect 30665 8449 30699 8483
rect 34529 8449 34563 8483
rect 11805 8381 11839 8415
rect 13645 8381 13679 8415
rect 17233 8381 17267 8415
rect 17509 8381 17543 8415
rect 21649 8381 21683 8415
rect 22477 8381 22511 8415
rect 30757 8381 30791 8415
rect 32137 8381 32171 8415
rect 32413 8381 32447 8415
rect 33885 8381 33919 8415
rect 16681 8313 16715 8347
rect 18613 8313 18647 8347
rect 22109 8313 22143 8347
rect 28365 8313 28399 8347
rect 13185 8245 13219 8279
rect 20085 8245 20119 8279
rect 21189 8245 21223 8279
rect 23305 8245 23339 8279
rect 30297 8245 30331 8279
rect 9873 8041 9907 8075
rect 17969 8041 18003 8075
rect 19993 8041 20027 8075
rect 20269 8041 20303 8075
rect 22201 8041 22235 8075
rect 23489 8041 23523 8075
rect 27077 8041 27111 8075
rect 27997 8041 28031 8075
rect 31309 8041 31343 8075
rect 32597 8041 32631 8075
rect 12357 7973 12391 8007
rect 21925 7973 21959 8007
rect 23029 7973 23063 8007
rect 23949 7973 23983 8007
rect 7757 7905 7791 7939
rect 7941 7905 7975 7939
rect 9597 7905 9631 7939
rect 12817 7905 12851 7939
rect 13001 7905 13035 7939
rect 17141 7905 17175 7939
rect 18061 7905 18095 7939
rect 20637 7905 20671 7939
rect 21281 7905 21315 7939
rect 21373 7905 21407 7939
rect 27721 7905 27755 7939
rect 29561 7905 29595 7939
rect 31953 7905 31987 7939
rect 6929 7837 6963 7871
rect 7665 7837 7699 7871
rect 9321 7837 9355 7871
rect 13737 7837 13771 7871
rect 14105 7837 14139 7871
rect 16865 7837 16899 7871
rect 17325 7837 17359 7871
rect 17418 7837 17452 7871
rect 17831 7837 17865 7871
rect 18245 7837 18279 7871
rect 20177 7837 20211 7871
rect 21189 7837 21223 7871
rect 22017 7837 22051 7871
rect 22845 7837 22879 7871
rect 23029 7837 23063 7871
rect 23121 7837 23155 7871
rect 23489 7837 23523 7871
rect 23857 7837 23891 7871
rect 27445 7837 27479 7871
rect 27537 7837 27571 7871
rect 32229 7837 32263 7871
rect 34529 7837 34563 7871
rect 8217 7769 8251 7803
rect 14933 7769 14967 7803
rect 17601 7769 17635 7803
rect 17693 7769 17727 7803
rect 21741 7769 21775 7803
rect 29837 7769 29871 7803
rect 32873 7769 32907 7803
rect 34253 7769 34287 7803
rect 7297 7701 7331 7735
rect 8953 7701 8987 7735
rect 9413 7701 9447 7735
rect 12725 7701 12759 7735
rect 16497 7701 16531 7735
rect 16957 7701 16991 7735
rect 20453 7701 20487 7735
rect 20821 7701 20855 7735
rect 23305 7701 23339 7735
rect 32137 7701 32171 7735
rect 32689 7701 32723 7735
rect 33241 7701 33275 7735
rect 7849 7497 7883 7531
rect 9321 7497 9355 7531
rect 10793 7497 10827 7531
rect 12909 7497 12943 7531
rect 13277 7497 13311 7531
rect 14013 7497 14047 7531
rect 14197 7497 14231 7531
rect 14565 7497 14599 7531
rect 15117 7497 15151 7531
rect 18797 7497 18831 7531
rect 20361 7497 20395 7531
rect 20821 7497 20855 7531
rect 21833 7497 21867 7531
rect 22017 7497 22051 7531
rect 22477 7497 22511 7531
rect 23121 7497 23155 7531
rect 23581 7497 23615 7531
rect 23765 7497 23799 7531
rect 31585 7497 31619 7531
rect 31953 7497 31987 7531
rect 32321 7497 32355 7531
rect 32689 7497 32723 7531
rect 14657 7429 14691 7463
rect 19156 7429 19190 7463
rect 24133 7429 24167 7463
rect 28825 7429 28859 7463
rect 29101 7429 29135 7463
rect 1501 7361 1535 7395
rect 1961 7361 1995 7395
rect 6469 7361 6503 7395
rect 6736 7361 6770 7395
rect 7941 7361 7975 7395
rect 8208 7361 8242 7395
rect 9413 7361 9447 7395
rect 9680 7361 9714 7395
rect 11529 7361 11563 7395
rect 11785 7361 11819 7395
rect 17684 7361 17718 7395
rect 18889 7361 18923 7395
rect 20729 7361 20763 7395
rect 22385 7361 22419 7395
rect 22753 7361 22787 7395
rect 22845 7361 22879 7395
rect 22937 7361 22971 7395
rect 23213 7361 23247 7395
rect 23306 7361 23340 7395
rect 23924 7361 23958 7395
rect 24501 7361 24535 7395
rect 24777 7361 24811 7395
rect 25053 7361 25087 7395
rect 25329 7361 25363 7395
rect 25421 7361 25455 7395
rect 25513 7361 25547 7395
rect 25697 7361 25731 7395
rect 26065 7361 26099 7395
rect 26157 7361 26191 7395
rect 26341 7361 26375 7395
rect 28733 7361 28767 7395
rect 28917 7361 28951 7395
rect 29285 7361 29319 7395
rect 31217 7361 31251 7395
rect 32229 7361 32263 7395
rect 32597 7361 32631 7395
rect 33057 7361 33091 7395
rect 14841 7293 14875 7327
rect 17417 7293 17451 7327
rect 20913 7293 20947 7327
rect 24041 7293 24075 7327
rect 24409 7293 24443 7327
rect 25145 7293 25179 7327
rect 31309 7293 31343 7327
rect 33241 7293 33275 7327
rect 33517 7293 33551 7327
rect 1685 7225 1719 7259
rect 1777 7225 1811 7259
rect 20269 7225 20303 7259
rect 21557 7157 21591 7191
rect 26433 7157 26467 7191
rect 29377 7157 29411 7191
rect 32965 7157 32999 7191
rect 34989 7157 35023 7191
rect 10057 6953 10091 6987
rect 11529 6953 11563 6987
rect 17325 6953 17359 6987
rect 17877 6953 17911 6987
rect 20269 6953 20303 6987
rect 21741 6953 21775 6987
rect 24041 6953 24075 6987
rect 24869 6953 24903 6987
rect 26065 6953 26099 6987
rect 27549 6953 27583 6987
rect 32229 6953 32263 6987
rect 33885 6953 33919 6987
rect 32965 6885 32999 6919
rect 10517 6817 10551 6851
rect 10701 6817 10735 6851
rect 11437 6817 11471 6851
rect 11989 6817 12023 6851
rect 12173 6817 12207 6851
rect 12449 6817 12483 6851
rect 15945 6817 15979 6851
rect 18521 6817 18555 6851
rect 20361 6817 20395 6851
rect 24567 6817 24601 6851
rect 28641 6817 28675 6851
rect 29101 6817 29135 6851
rect 30849 6817 30883 6851
rect 10425 6749 10459 6783
rect 11897 6749 11931 6783
rect 14105 6749 14139 6783
rect 16212 6749 16246 6783
rect 18245 6749 18279 6783
rect 18797 6749 18831 6783
rect 21925 6749 21959 6783
rect 22753 6749 22787 6783
rect 23397 6749 23431 6783
rect 23673 6749 23707 6783
rect 23765 6749 23799 6783
rect 24409 6749 24443 6783
rect 24777 6749 24811 6783
rect 25053 6749 25087 6783
rect 25421 6749 25455 6783
rect 25513 6749 25547 6783
rect 27813 6749 27847 6783
rect 29009 6749 29043 6783
rect 29929 6749 29963 6783
rect 31033 6749 31067 6783
rect 31309 6749 31343 6783
rect 31493 6749 31527 6783
rect 31677 6749 31711 6783
rect 31861 6749 31895 6783
rect 31953 6749 31987 6783
rect 32505 6749 32539 6783
rect 32597 6749 32631 6783
rect 32781 6749 32815 6783
rect 33149 6749 33183 6783
rect 33701 6749 33735 6783
rect 34069 6749 34103 6783
rect 34253 6749 34287 6783
rect 34345 6749 34379 6783
rect 10977 6681 11011 6715
rect 14350 6681 14384 6715
rect 18337 6681 18371 6715
rect 20628 6681 20662 6715
rect 25145 6681 25179 6715
rect 32208 6681 32242 6715
rect 32413 6681 32447 6715
rect 33425 6681 33459 6715
rect 33609 6681 33643 6715
rect 15485 6613 15519 6647
rect 23949 6613 23983 6647
rect 25329 6613 25363 6647
rect 25697 6613 25731 6647
rect 31217 6613 31251 6647
rect 32045 6613 32079 6647
rect 14197 6409 14231 6443
rect 14565 6409 14599 6443
rect 14657 6409 14691 6443
rect 15025 6409 15059 6443
rect 21281 6409 21315 6443
rect 25789 6409 25823 6443
rect 28825 6409 28859 6443
rect 31309 6409 31343 6443
rect 32137 6409 32171 6443
rect 32781 6409 32815 6443
rect 33425 6409 33459 6443
rect 29193 6341 29227 6375
rect 31585 6341 31619 6375
rect 33609 6341 33643 6375
rect 21097 6273 21131 6307
rect 21281 6273 21315 6307
rect 21465 6273 21499 6307
rect 22293 6273 22327 6307
rect 23121 6273 23155 6307
rect 23489 6273 23523 6307
rect 23765 6273 23799 6307
rect 24593 6273 24627 6307
rect 24777 6273 24811 6307
rect 24869 6273 24903 6307
rect 25421 6273 25455 6307
rect 28733 6273 28767 6307
rect 30573 6273 30607 6307
rect 31217 6273 31251 6307
rect 31401 6273 31435 6307
rect 31493 6273 31527 6307
rect 31677 6273 31711 6307
rect 32321 6273 32355 6307
rect 32873 6273 32907 6307
rect 33333 6273 33367 6307
rect 14841 6205 14875 6239
rect 23397 6205 23431 6239
rect 25513 6205 25547 6239
rect 28917 6205 28951 6239
rect 29929 6205 29963 6239
rect 30205 6205 30239 6239
rect 30481 6205 30515 6239
rect 32597 6205 32631 6239
rect 33053 6205 33087 6239
rect 31861 6137 31895 6171
rect 33149 6137 33183 6171
rect 21557 6069 21591 6103
rect 24409 6069 24443 6103
rect 25053 6069 25087 6103
rect 28365 6069 28399 6103
rect 32505 6069 32539 6103
rect 33241 6069 33275 6103
rect 22937 5865 22971 5899
rect 28825 5865 28859 5899
rect 29101 5865 29135 5899
rect 31217 5865 31251 5899
rect 33977 5865 34011 5899
rect 30849 5797 30883 5831
rect 33701 5797 33735 5831
rect 34069 5797 34103 5831
rect 21189 5729 21223 5763
rect 23489 5729 23523 5763
rect 23949 5729 23983 5763
rect 24133 5729 24167 5763
rect 27077 5729 27111 5763
rect 31033 5729 31067 5763
rect 33333 5729 33367 5763
rect 33885 5729 33919 5763
rect 23581 5661 23615 5695
rect 23765 5661 23799 5695
rect 29745 5661 29779 5695
rect 29929 5661 29963 5695
rect 30205 5661 30239 5695
rect 30389 5661 30423 5695
rect 30481 5661 30515 5695
rect 30573 5661 30607 5695
rect 30665 5661 30699 5695
rect 30941 5661 30975 5695
rect 31217 5661 31251 5695
rect 33517 5661 33551 5695
rect 33793 5661 33827 5695
rect 34161 5661 34195 5695
rect 34345 5661 34379 5695
rect 34437 5661 34471 5695
rect 21465 5593 21499 5627
rect 23121 5593 23155 5627
rect 23305 5593 23339 5627
rect 27353 5593 27387 5627
rect 29561 5593 29595 5627
rect 29837 5593 29871 5627
rect 30047 5593 30081 5627
rect 33149 5593 33183 5627
rect 29285 5525 29319 5559
rect 31401 5525 31435 5559
rect 26249 5321 26283 5355
rect 30481 5321 30515 5355
rect 33701 5321 33735 5355
rect 1501 5185 1535 5219
rect 1961 5185 1995 5219
rect 23581 5185 23615 5219
rect 24041 5185 24075 5219
rect 24501 5185 24535 5219
rect 30665 5185 30699 5219
rect 33977 5185 34011 5219
rect 34161 5185 34195 5219
rect 34253 5185 34287 5219
rect 34437 5185 34471 5219
rect 34529 5185 34563 5219
rect 23305 5117 23339 5151
rect 23949 5117 23983 5151
rect 24777 5117 24811 5151
rect 30941 5117 30975 5151
rect 34345 5117 34379 5151
rect 34805 5117 34839 5151
rect 24409 5049 24443 5083
rect 1593 4981 1627 5015
rect 1869 4981 1903 5015
rect 30849 4981 30883 5015
rect 34161 4981 34195 5015
rect 31769 4709 31803 4743
rect 32413 4709 32447 4743
rect 22477 4641 22511 4675
rect 30297 4641 30331 4675
rect 30573 4641 30607 4675
rect 31309 4641 31343 4675
rect 31953 4641 31987 4675
rect 30665 4573 30699 4607
rect 31401 4573 31435 4607
rect 32045 4573 32079 4607
rect 32689 4573 32723 4607
rect 22753 4505 22787 4539
rect 32965 4505 32999 4539
rect 24225 4437 24259 4471
rect 34437 4437 34471 4471
rect 22477 4233 22511 4267
rect 32781 4233 32815 4267
rect 33241 4233 33275 4267
rect 32873 4165 32907 4199
rect 22845 4097 22879 4131
rect 28641 4097 28675 4131
rect 29101 4097 29135 4131
rect 30941 4097 30975 4131
rect 31125 4097 31159 4131
rect 22937 4029 22971 4063
rect 28733 4029 28767 4063
rect 29377 4029 29411 4063
rect 32597 4029 32631 4063
rect 29009 3893 29043 3927
rect 30849 3893 30883 3927
rect 29837 3689 29871 3723
rect 30297 3553 30331 3587
rect 30389 3553 30423 3587
rect 1409 3485 1443 3519
rect 1869 3485 1903 3519
rect 30205 3485 30239 3519
rect 34069 3485 34103 3519
rect 1777 3417 1811 3451
rect 34345 3417 34379 3451
rect 1593 3349 1627 3383
<< metal1 >>
rect 1104 35930 35328 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35328 35930
rect 1104 35856 35328 35878
rect 1210 35708 1216 35760
rect 1268 35748 1274 35760
rect 18877 35751 18935 35757
rect 18877 35748 18889 35751
rect 1268 35720 1716 35748
rect 1268 35708 1274 35720
rect 1302 35640 1308 35692
rect 1360 35680 1366 35692
rect 1688 35689 1716 35720
rect 2746 35720 18889 35748
rect 1397 35683 1455 35689
rect 1397 35680 1409 35683
rect 1360 35652 1409 35680
rect 1360 35640 1366 35652
rect 1397 35649 1409 35652
rect 1443 35649 1455 35683
rect 1397 35643 1455 35649
rect 1673 35683 1731 35689
rect 1673 35649 1685 35683
rect 1719 35680 1731 35683
rect 1949 35683 2007 35689
rect 1949 35680 1961 35683
rect 1719 35652 1961 35680
rect 1719 35649 1731 35652
rect 1673 35643 1731 35649
rect 1949 35649 1961 35652
rect 1995 35649 2007 35683
rect 1949 35643 2007 35649
rect 2746 35612 2774 35720
rect 18877 35717 18889 35720
rect 18923 35717 18935 35751
rect 18877 35711 18935 35717
rect 19613 35751 19671 35757
rect 19613 35717 19625 35751
rect 19659 35748 19671 35751
rect 19702 35748 19708 35760
rect 19659 35720 19708 35748
rect 19659 35717 19671 35720
rect 19613 35711 19671 35717
rect 19702 35708 19708 35720
rect 19760 35708 19766 35760
rect 10962 35640 10968 35692
rect 11020 35680 11026 35692
rect 11885 35683 11943 35689
rect 11885 35680 11897 35683
rect 11020 35652 11897 35680
rect 11020 35640 11026 35652
rect 11885 35649 11897 35652
rect 11931 35649 11943 35683
rect 11885 35643 11943 35649
rect 18509 35683 18567 35689
rect 18509 35649 18521 35683
rect 18555 35680 18567 35683
rect 18555 35652 19012 35680
rect 18555 35649 18567 35652
rect 18509 35643 18567 35649
rect 1596 35584 2774 35612
rect 11977 35615 12035 35621
rect 1596 35553 1624 35584
rect 11977 35581 11989 35615
rect 12023 35612 12035 35615
rect 12066 35612 12072 35624
rect 12023 35584 12072 35612
rect 12023 35581 12035 35584
rect 11977 35575 12035 35581
rect 12066 35572 12072 35584
rect 12124 35572 12130 35624
rect 12161 35615 12219 35621
rect 12161 35581 12173 35615
rect 12207 35612 12219 35615
rect 12207 35584 12480 35612
rect 12207 35581 12219 35584
rect 12161 35575 12219 35581
rect 1581 35547 1639 35553
rect 1581 35513 1593 35547
rect 1627 35513 1639 35547
rect 1581 35507 1639 35513
rect 1857 35547 1915 35553
rect 1857 35513 1869 35547
rect 1903 35544 1915 35547
rect 3602 35544 3608 35556
rect 1903 35516 3608 35544
rect 1903 35513 1915 35516
rect 1857 35507 1915 35513
rect 3602 35504 3608 35516
rect 3660 35504 3666 35556
rect 11330 35436 11336 35488
rect 11388 35476 11394 35488
rect 12452 35485 12480 35584
rect 11517 35479 11575 35485
rect 11517 35476 11529 35479
rect 11388 35448 11529 35476
rect 11388 35436 11394 35448
rect 11517 35445 11529 35448
rect 11563 35445 11575 35479
rect 11517 35439 11575 35445
rect 12437 35479 12495 35485
rect 12437 35445 12449 35479
rect 12483 35476 12495 35479
rect 13998 35476 14004 35488
rect 12483 35448 14004 35476
rect 12483 35445 12495 35448
rect 12437 35439 12495 35445
rect 13998 35436 14004 35448
rect 14056 35436 14062 35488
rect 18693 35479 18751 35485
rect 18693 35445 18705 35479
rect 18739 35476 18751 35479
rect 18874 35476 18880 35488
rect 18739 35448 18880 35476
rect 18739 35445 18751 35448
rect 18693 35439 18751 35445
rect 18874 35436 18880 35448
rect 18932 35436 18938 35488
rect 18984 35485 19012 35652
rect 25682 35640 25688 35692
rect 25740 35640 25746 35692
rect 27893 35683 27951 35689
rect 27893 35649 27905 35683
rect 27939 35680 27951 35683
rect 28718 35680 28724 35692
rect 27939 35652 28724 35680
rect 27939 35649 27951 35652
rect 27893 35643 27951 35649
rect 28718 35640 28724 35652
rect 28776 35640 28782 35692
rect 34514 35640 34520 35692
rect 34572 35640 34578 35692
rect 19058 35572 19064 35624
rect 19116 35612 19122 35624
rect 19705 35615 19763 35621
rect 19705 35612 19717 35615
rect 19116 35584 19717 35612
rect 19116 35572 19122 35584
rect 19705 35581 19717 35584
rect 19751 35581 19763 35615
rect 19705 35575 19763 35581
rect 19889 35615 19947 35621
rect 19889 35581 19901 35615
rect 19935 35581 19947 35615
rect 19889 35575 19947 35581
rect 25501 35615 25559 35621
rect 25501 35581 25513 35615
rect 25547 35581 25559 35615
rect 25501 35575 25559 35581
rect 19904 35544 19932 35575
rect 20165 35547 20223 35553
rect 20165 35544 20177 35547
rect 19904 35516 20177 35544
rect 20165 35513 20177 35516
rect 20211 35544 20223 35547
rect 25516 35544 25544 35575
rect 25590 35572 25596 35624
rect 25648 35572 25654 35624
rect 27982 35572 27988 35624
rect 28040 35572 28046 35624
rect 28077 35615 28135 35621
rect 28077 35581 28089 35615
rect 28123 35581 28135 35615
rect 28077 35575 28135 35581
rect 28092 35544 28120 35575
rect 34330 35572 34336 35624
rect 34388 35572 34394 35624
rect 20211 35516 26280 35544
rect 20211 35513 20223 35516
rect 20165 35507 20223 35513
rect 26252 35488 26280 35516
rect 27448 35516 28120 35544
rect 27448 35488 27476 35516
rect 18969 35479 19027 35485
rect 18969 35445 18981 35479
rect 19015 35476 19027 35479
rect 19150 35476 19156 35488
rect 19015 35448 19156 35476
rect 19015 35445 19027 35448
rect 18969 35439 19027 35445
rect 19150 35436 19156 35448
rect 19208 35436 19214 35488
rect 19242 35436 19248 35488
rect 19300 35436 19306 35488
rect 26050 35436 26056 35488
rect 26108 35436 26114 35488
rect 26234 35436 26240 35488
rect 26292 35436 26298 35488
rect 27430 35436 27436 35488
rect 27488 35436 27494 35488
rect 27525 35479 27583 35485
rect 27525 35445 27537 35479
rect 27571 35476 27583 35479
rect 27614 35476 27620 35488
rect 27571 35448 27620 35476
rect 27571 35445 27583 35448
rect 27525 35439 27583 35445
rect 27614 35436 27620 35448
rect 27672 35436 27678 35488
rect 1104 35386 35328 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 35328 35386
rect 1104 35312 35328 35334
rect 1302 35232 1308 35284
rect 1360 35272 1366 35284
rect 1397 35275 1455 35281
rect 1397 35272 1409 35275
rect 1360 35244 1409 35272
rect 1360 35232 1366 35244
rect 1397 35241 1409 35244
rect 1443 35241 1455 35275
rect 1397 35235 1455 35241
rect 9030 35232 9036 35284
rect 9088 35272 9094 35284
rect 17218 35272 17224 35284
rect 9088 35244 17224 35272
rect 9088 35232 9094 35244
rect 17218 35232 17224 35244
rect 17276 35232 17282 35284
rect 19058 35232 19064 35284
rect 19116 35232 19122 35284
rect 19150 35232 19156 35284
rect 19208 35272 19214 35284
rect 19208 35244 25544 35272
rect 19208 35232 19214 35244
rect 25516 35204 25544 35244
rect 25590 35232 25596 35284
rect 25648 35272 25654 35284
rect 25869 35275 25927 35281
rect 25869 35272 25881 35275
rect 25648 35244 25881 35272
rect 25648 35232 25654 35244
rect 25869 35241 25881 35244
rect 25915 35241 25927 35275
rect 27982 35272 27988 35284
rect 25869 35235 25927 35241
rect 26344 35244 27988 35272
rect 26344 35204 26372 35244
rect 27982 35232 27988 35244
rect 28040 35232 28046 35284
rect 28442 35232 28448 35284
rect 28500 35272 28506 35284
rect 28718 35272 28724 35284
rect 28500 35244 28724 35272
rect 28500 35232 28506 35244
rect 28718 35232 28724 35244
rect 28776 35232 28782 35284
rect 25516 35176 26372 35204
rect 13998 35096 14004 35148
rect 14056 35136 14062 35148
rect 14645 35139 14703 35145
rect 14645 35136 14657 35139
rect 14056 35108 14657 35136
rect 14056 35096 14062 35108
rect 14645 35105 14657 35108
rect 14691 35136 14703 35139
rect 14921 35139 14979 35145
rect 14921 35136 14933 35139
rect 14691 35108 14933 35136
rect 14691 35105 14703 35108
rect 14645 35099 14703 35105
rect 14921 35105 14933 35108
rect 14967 35105 14979 35139
rect 14921 35099 14979 35105
rect 7098 35028 7104 35080
rect 7156 35068 7162 35080
rect 7377 35071 7435 35077
rect 7377 35068 7389 35071
rect 7156 35040 7389 35068
rect 7156 35028 7162 35040
rect 7377 35037 7389 35040
rect 7423 35037 7435 35071
rect 7377 35031 7435 35037
rect 9493 35071 9551 35077
rect 9493 35037 9505 35071
rect 9539 35068 9551 35071
rect 11057 35071 11115 35077
rect 11057 35068 11069 35071
rect 9539 35040 11069 35068
rect 9539 35037 9551 35040
rect 9493 35031 9551 35037
rect 11057 35037 11069 35040
rect 11103 35068 11115 35071
rect 11103 35040 11560 35068
rect 11103 35037 11115 35040
rect 11057 35031 11115 35037
rect 11532 35012 11560 35040
rect 11882 35028 11888 35080
rect 11940 35068 11946 35080
rect 13817 35071 13875 35077
rect 13817 35068 13829 35071
rect 11940 35040 13829 35068
rect 11940 35028 11946 35040
rect 13817 35037 13829 35040
rect 13863 35068 13875 35071
rect 14553 35071 14611 35077
rect 14553 35068 14565 35071
rect 13863 35040 14565 35068
rect 13863 35037 13875 35040
rect 13817 35031 13875 35037
rect 14553 35037 14565 35040
rect 14599 35037 14611 35071
rect 14553 35031 14611 35037
rect 15102 35028 15108 35080
rect 15160 35028 15166 35080
rect 17402 35028 17408 35080
rect 17460 35068 17466 35080
rect 17681 35071 17739 35077
rect 17681 35068 17693 35071
rect 17460 35040 17693 35068
rect 17460 35028 17466 35040
rect 17681 35037 17693 35040
rect 17727 35037 17739 35071
rect 17681 35031 17739 35037
rect 17948 35071 18006 35077
rect 17948 35037 17960 35071
rect 17994 35068 18006 35071
rect 19242 35068 19248 35080
rect 17994 35040 19248 35068
rect 17994 35037 18006 35040
rect 17948 35031 18006 35037
rect 19242 35028 19248 35040
rect 19300 35028 19306 35080
rect 19613 35071 19671 35077
rect 19613 35037 19625 35071
rect 19659 35068 19671 35071
rect 22186 35068 22192 35080
rect 19659 35040 22192 35068
rect 19659 35037 19671 35040
rect 19613 35031 19671 35037
rect 22186 35028 22192 35040
rect 22244 35068 22250 35080
rect 24397 35071 24455 35077
rect 24397 35068 24409 35071
rect 22244 35040 24409 35068
rect 22244 35028 22250 35040
rect 24397 35037 24409 35040
rect 24443 35037 24455 35071
rect 24397 35031 24455 35037
rect 26050 35028 26056 35080
rect 26108 35068 26114 35080
rect 26982 35071 27040 35077
rect 26982 35068 26994 35071
rect 26108 35040 26994 35068
rect 26108 35028 26114 35040
rect 26982 35037 26994 35040
rect 27028 35037 27040 35071
rect 26982 35031 27040 35037
rect 27246 35028 27252 35080
rect 27304 35068 27310 35080
rect 27614 35077 27620 35080
rect 27341 35071 27399 35077
rect 27341 35068 27353 35071
rect 27304 35040 27353 35068
rect 27304 35028 27310 35040
rect 27341 35037 27353 35040
rect 27387 35037 27399 35071
rect 27608 35068 27620 35077
rect 27575 35040 27620 35068
rect 27341 35031 27399 35037
rect 27608 35031 27620 35040
rect 27614 35028 27620 35031
rect 27672 35028 27678 35080
rect 7644 35003 7702 35009
rect 7644 34969 7656 35003
rect 7690 35000 7702 35003
rect 8110 35000 8116 35012
rect 7690 34972 8116 35000
rect 7690 34969 7702 34972
rect 7644 34963 7702 34969
rect 8110 34960 8116 34972
rect 8168 34960 8174 35012
rect 9582 34960 9588 35012
rect 9640 35000 9646 35012
rect 11330 35009 11336 35012
rect 9738 35003 9796 35009
rect 9738 35000 9750 35003
rect 9640 34972 9750 35000
rect 9640 34960 9646 34972
rect 9738 34969 9750 34972
rect 9784 34969 9796 35003
rect 11324 35000 11336 35009
rect 11291 34972 11336 35000
rect 9738 34963 9796 34969
rect 11324 34963 11336 34972
rect 11330 34960 11336 34963
rect 11388 34960 11394 35012
rect 11514 34960 11520 35012
rect 11572 34960 11578 35012
rect 15372 35003 15430 35009
rect 15372 34969 15384 35003
rect 15418 35000 15430 35003
rect 15562 35000 15568 35012
rect 15418 34972 15568 35000
rect 15418 34969 15430 34972
rect 15372 34963 15430 34969
rect 15562 34960 15568 34972
rect 15620 34960 15626 35012
rect 19880 35003 19938 35009
rect 19880 34969 19892 35003
rect 19926 35000 19938 35003
rect 20162 35000 20168 35012
rect 19926 34972 20168 35000
rect 19926 34969 19938 34972
rect 19880 34963 19938 34969
rect 20162 34960 20168 34972
rect 20220 34960 20226 35012
rect 22456 35003 22514 35009
rect 22456 34969 22468 35003
rect 22502 35000 22514 35003
rect 23290 35000 23296 35012
rect 22502 34972 23296 35000
rect 22502 34969 22514 34972
rect 22456 34963 22514 34969
rect 23290 34960 23296 34972
rect 23348 34960 23354 35012
rect 24670 35009 24676 35012
rect 24664 34963 24676 35009
rect 24670 34960 24676 34963
rect 24728 34960 24734 35012
rect 8754 34892 8760 34944
rect 8812 34892 8818 34944
rect 10870 34892 10876 34944
rect 10928 34892 10934 34944
rect 10962 34892 10968 34944
rect 11020 34932 11026 34944
rect 12437 34935 12495 34941
rect 12437 34932 12449 34935
rect 11020 34904 12449 34932
rect 11020 34892 11026 34904
rect 12437 34901 12449 34904
rect 12483 34901 12495 34935
rect 12437 34895 12495 34901
rect 13630 34892 13636 34944
rect 13688 34892 13694 34944
rect 13722 34892 13728 34944
rect 13780 34932 13786 34944
rect 14093 34935 14151 34941
rect 14093 34932 14105 34935
rect 13780 34904 14105 34932
rect 13780 34892 13786 34904
rect 14093 34901 14105 34904
rect 14139 34901 14151 34935
rect 14093 34895 14151 34901
rect 14458 34892 14464 34944
rect 14516 34892 14522 34944
rect 16022 34892 16028 34944
rect 16080 34932 16086 34944
rect 16485 34935 16543 34941
rect 16485 34932 16497 34935
rect 16080 34904 16497 34932
rect 16080 34892 16086 34904
rect 16485 34901 16497 34904
rect 16531 34901 16543 34935
rect 16485 34895 16543 34901
rect 20990 34892 20996 34944
rect 21048 34892 21054 34944
rect 23566 34892 23572 34944
rect 23624 34892 23630 34944
rect 25774 34892 25780 34944
rect 25832 34892 25838 34944
rect 1104 34842 35328 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35328 34842
rect 1104 34768 35328 34790
rect 8110 34688 8116 34740
rect 8168 34688 8174 34740
rect 9030 34688 9036 34740
rect 9088 34688 9094 34740
rect 9582 34688 9588 34740
rect 9640 34688 9646 34740
rect 9953 34731 10011 34737
rect 9953 34697 9965 34731
rect 9999 34728 10011 34731
rect 10594 34728 10600 34740
rect 9999 34700 10600 34728
rect 9999 34697 10011 34700
rect 9953 34691 10011 34697
rect 10594 34688 10600 34700
rect 10652 34728 10658 34740
rect 10870 34728 10876 34740
rect 10652 34700 10876 34728
rect 10652 34688 10658 34700
rect 10870 34688 10876 34700
rect 10928 34688 10934 34740
rect 14458 34688 14464 34740
rect 14516 34728 14522 34740
rect 14829 34731 14887 34737
rect 14829 34728 14841 34731
rect 14516 34700 14841 34728
rect 14516 34688 14522 34700
rect 14829 34697 14841 34700
rect 14875 34697 14887 34731
rect 14829 34691 14887 34697
rect 15562 34688 15568 34740
rect 15620 34688 15626 34740
rect 16022 34688 16028 34740
rect 16080 34688 16086 34740
rect 20162 34688 20168 34740
rect 20220 34688 20226 34740
rect 20533 34731 20591 34737
rect 20533 34697 20545 34731
rect 20579 34728 20591 34731
rect 20714 34728 20720 34740
rect 20579 34700 20720 34728
rect 20579 34697 20591 34700
rect 20533 34691 20591 34697
rect 20714 34688 20720 34700
rect 20772 34728 20778 34740
rect 20990 34728 20996 34740
rect 20772 34700 20996 34728
rect 20772 34688 20778 34700
rect 20990 34688 20996 34700
rect 21048 34688 21054 34740
rect 21100 34700 23244 34728
rect 8573 34663 8631 34669
rect 8573 34629 8585 34663
rect 8619 34660 8631 34663
rect 10410 34660 10416 34672
rect 8619 34632 10416 34660
rect 8619 34629 8631 34632
rect 8573 34623 8631 34629
rect 10410 34620 10416 34632
rect 10468 34620 10474 34672
rect 14090 34660 14096 34672
rect 13464 34632 14096 34660
rect 8481 34595 8539 34601
rect 8481 34561 8493 34595
rect 8527 34592 8539 34595
rect 8754 34592 8760 34604
rect 8527 34564 8760 34592
rect 8527 34561 8539 34564
rect 8481 34555 8539 34561
rect 8754 34552 8760 34564
rect 8812 34592 8818 34604
rect 9674 34592 9680 34604
rect 8812 34564 9680 34592
rect 8812 34552 8818 34564
rect 9674 34552 9680 34564
rect 9732 34552 9738 34604
rect 10045 34595 10103 34601
rect 10045 34561 10057 34595
rect 10091 34592 10103 34595
rect 10689 34595 10747 34601
rect 10689 34592 10701 34595
rect 10091 34564 10701 34592
rect 10091 34561 10103 34564
rect 10045 34555 10103 34561
rect 10689 34561 10701 34564
rect 10735 34592 10747 34595
rect 12066 34592 12072 34604
rect 10735 34564 12072 34592
rect 10735 34561 10747 34564
rect 10689 34555 10747 34561
rect 12066 34552 12072 34564
rect 12124 34552 12130 34604
rect 12244 34595 12302 34601
rect 12244 34561 12256 34595
rect 12290 34592 12302 34595
rect 13170 34592 13176 34604
rect 12290 34564 13176 34592
rect 12290 34561 12302 34564
rect 12244 34555 12302 34561
rect 13170 34552 13176 34564
rect 13228 34552 13234 34604
rect 13464 34601 13492 34632
rect 14090 34620 14096 34632
rect 14148 34660 14154 34672
rect 15102 34660 15108 34672
rect 14148 34632 15108 34660
rect 14148 34620 14154 34632
rect 15102 34620 15108 34632
rect 15160 34620 15166 34672
rect 17218 34620 17224 34672
rect 17276 34660 17282 34672
rect 21100 34660 21128 34700
rect 22186 34660 22192 34672
rect 17276 34632 21128 34660
rect 21836 34632 22192 34660
rect 17276 34620 17282 34632
rect 13722 34601 13728 34604
rect 13449 34595 13507 34601
rect 13449 34561 13461 34595
rect 13495 34561 13507 34595
rect 13716 34592 13728 34601
rect 13683 34564 13728 34592
rect 13449 34555 13507 34561
rect 13716 34555 13728 34564
rect 13722 34552 13728 34555
rect 13780 34552 13786 34604
rect 15933 34595 15991 34601
rect 15933 34561 15945 34595
rect 15979 34561 15991 34595
rect 15933 34555 15991 34561
rect 8665 34527 8723 34533
rect 8665 34493 8677 34527
rect 8711 34524 8723 34527
rect 9030 34524 9036 34536
rect 8711 34496 9036 34524
rect 8711 34493 8723 34496
rect 8665 34487 8723 34493
rect 9030 34484 9036 34496
rect 9088 34524 9094 34536
rect 9398 34524 9404 34536
rect 9088 34496 9404 34524
rect 9088 34484 9094 34496
rect 9398 34484 9404 34496
rect 9456 34484 9462 34536
rect 10229 34527 10287 34533
rect 10229 34493 10241 34527
rect 10275 34493 10287 34527
rect 10229 34487 10287 34493
rect 10244 34456 10272 34487
rect 10410 34484 10416 34536
rect 10468 34484 10474 34536
rect 11514 34484 11520 34536
rect 11572 34524 11578 34536
rect 11977 34527 12035 34533
rect 11977 34524 11989 34527
rect 11572 34496 11989 34524
rect 11572 34484 11578 34496
rect 11977 34493 11989 34496
rect 12023 34493 12035 34527
rect 11977 34487 12035 34493
rect 10318 34456 10324 34468
rect 10244 34428 10324 34456
rect 10318 34416 10324 34428
rect 10376 34456 10382 34468
rect 11606 34456 11612 34468
rect 10376 34428 11612 34456
rect 10376 34416 10382 34428
rect 11606 34416 11612 34428
rect 11664 34416 11670 34468
rect 13354 34348 13360 34400
rect 13412 34348 13418 34400
rect 13630 34348 13636 34400
rect 13688 34388 13694 34400
rect 15948 34388 15976 34555
rect 18322 34552 18328 34604
rect 18380 34552 18386 34604
rect 21836 34601 21864 34632
rect 22186 34620 22192 34632
rect 22244 34660 22250 34672
rect 22554 34660 22560 34672
rect 22244 34632 22560 34660
rect 22244 34620 22250 34632
rect 22554 34620 22560 34632
rect 22612 34620 22618 34672
rect 23216 34660 23244 34700
rect 23290 34688 23296 34740
rect 23348 34688 23354 34740
rect 23566 34688 23572 34740
rect 23624 34728 23630 34740
rect 23661 34731 23719 34737
rect 23661 34728 23673 34731
rect 23624 34700 23673 34728
rect 23624 34688 23630 34700
rect 23661 34697 23673 34700
rect 23707 34697 23719 34731
rect 23661 34691 23719 34697
rect 24581 34731 24639 34737
rect 24581 34697 24593 34731
rect 24627 34728 24639 34731
rect 24670 34728 24676 34740
rect 24627 34700 24676 34728
rect 24627 34697 24639 34700
rect 24581 34691 24639 34697
rect 24670 34688 24676 34700
rect 24728 34688 24734 34740
rect 24949 34731 25007 34737
rect 24949 34697 24961 34731
rect 24995 34728 25007 34731
rect 25314 34728 25320 34740
rect 24995 34700 25320 34728
rect 24995 34697 25007 34700
rect 24949 34691 25007 34697
rect 25314 34688 25320 34700
rect 25372 34728 25378 34740
rect 25774 34728 25780 34740
rect 25372 34700 25780 34728
rect 25372 34688 25378 34700
rect 25774 34688 25780 34700
rect 25832 34688 25838 34740
rect 27982 34688 27988 34740
rect 28040 34728 28046 34740
rect 28169 34731 28227 34737
rect 28169 34728 28181 34731
rect 28040 34700 28181 34728
rect 28040 34688 28046 34700
rect 28169 34697 28181 34700
rect 28215 34697 28227 34731
rect 28169 34691 28227 34697
rect 24397 34663 24455 34669
rect 24397 34660 24409 34663
rect 23216 34632 24409 34660
rect 24397 34629 24409 34632
rect 24443 34629 24455 34663
rect 24397 34623 24455 34629
rect 22094 34601 22100 34604
rect 20625 34595 20683 34601
rect 20625 34592 20637 34595
rect 18432 34564 20637 34592
rect 18432 34536 18460 34564
rect 20625 34561 20637 34564
rect 20671 34561 20683 34595
rect 20625 34555 20683 34561
rect 21821 34595 21879 34601
rect 21821 34561 21833 34595
rect 21867 34561 21879 34595
rect 21821 34555 21879 34561
rect 22088 34555 22100 34601
rect 22094 34552 22100 34555
rect 22152 34552 22158 34604
rect 23750 34552 23756 34604
rect 23808 34592 23814 34604
rect 24412 34592 24440 34623
rect 23808 34564 23980 34592
rect 24412 34564 25176 34592
rect 23808 34552 23814 34564
rect 16206 34484 16212 34536
rect 16264 34524 16270 34536
rect 16393 34527 16451 34533
rect 16393 34524 16405 34527
rect 16264 34496 16405 34524
rect 16264 34484 16270 34496
rect 16393 34493 16405 34496
rect 16439 34493 16451 34527
rect 16393 34487 16451 34493
rect 18414 34484 18420 34536
rect 18472 34484 18478 34536
rect 18601 34527 18659 34533
rect 18601 34493 18613 34527
rect 18647 34493 18659 34527
rect 18601 34487 18659 34493
rect 18785 34527 18843 34533
rect 18785 34493 18797 34527
rect 18831 34524 18843 34527
rect 18874 34524 18880 34536
rect 18831 34496 18880 34524
rect 18831 34493 18843 34496
rect 18785 34487 18843 34493
rect 18616 34456 18644 34487
rect 18874 34484 18880 34496
rect 18932 34484 18938 34536
rect 19061 34527 19119 34533
rect 19061 34493 19073 34527
rect 19107 34524 19119 34527
rect 19702 34524 19708 34536
rect 19107 34496 19708 34524
rect 19107 34493 19119 34496
rect 19061 34487 19119 34493
rect 19702 34484 19708 34496
rect 19760 34484 19766 34536
rect 19797 34527 19855 34533
rect 19797 34493 19809 34527
rect 19843 34493 19855 34527
rect 19797 34487 19855 34493
rect 19812 34456 19840 34487
rect 20806 34484 20812 34536
rect 20864 34524 20870 34536
rect 20993 34527 21051 34533
rect 20993 34524 21005 34527
rect 20864 34496 21005 34524
rect 20864 34484 20870 34496
rect 20993 34493 21005 34496
rect 21039 34493 21051 34527
rect 23845 34527 23903 34533
rect 23845 34524 23857 34527
rect 20993 34487 21051 34493
rect 23124 34496 23857 34524
rect 18616 34428 21128 34456
rect 16114 34388 16120 34400
rect 13688 34360 16120 34388
rect 13688 34348 13694 34360
rect 16114 34348 16120 34360
rect 16172 34348 16178 34400
rect 17678 34348 17684 34400
rect 17736 34388 17742 34400
rect 17957 34391 18015 34397
rect 17957 34388 17969 34391
rect 17736 34360 17969 34388
rect 17736 34348 17742 34360
rect 17957 34357 17969 34360
rect 18003 34357 18015 34391
rect 21100 34388 21128 34428
rect 22462 34388 22468 34400
rect 21100 34360 22468 34388
rect 17957 34351 18015 34357
rect 22462 34348 22468 34360
rect 22520 34388 22526 34400
rect 23124 34388 23152 34496
rect 23845 34493 23857 34496
rect 23891 34493 23903 34527
rect 23952 34524 23980 34564
rect 25148 34533 25176 34564
rect 28074 34552 28080 34604
rect 28132 34552 28138 34604
rect 25041 34527 25099 34533
rect 25041 34524 25053 34527
rect 23952 34496 25053 34524
rect 23845 34487 23903 34493
rect 25041 34493 25053 34496
rect 25087 34493 25099 34527
rect 25041 34487 25099 34493
rect 25133 34527 25191 34533
rect 25133 34493 25145 34527
rect 25179 34493 25191 34527
rect 25133 34487 25191 34493
rect 28261 34527 28319 34533
rect 28261 34493 28273 34527
rect 28307 34493 28319 34527
rect 28261 34487 28319 34493
rect 23860 34456 23888 34487
rect 24121 34459 24179 34465
rect 24121 34456 24133 34459
rect 23860 34428 24133 34456
rect 24121 34425 24133 34428
rect 24167 34425 24179 34459
rect 24121 34419 24179 34425
rect 27798 34416 27804 34468
rect 27856 34456 27862 34468
rect 28276 34456 28304 34487
rect 27856 34428 28304 34456
rect 27856 34416 27862 34428
rect 22520 34360 23152 34388
rect 22520 34348 22526 34360
rect 23198 34348 23204 34400
rect 23256 34348 23262 34400
rect 27614 34348 27620 34400
rect 27672 34388 27678 34400
rect 27709 34391 27767 34397
rect 27709 34388 27721 34391
rect 27672 34360 27721 34388
rect 27672 34348 27678 34360
rect 27709 34357 27721 34360
rect 27755 34357 27767 34391
rect 27709 34351 27767 34357
rect 1104 34298 35328 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 35328 34298
rect 1104 34224 35328 34246
rect 13170 34144 13176 34196
rect 13228 34144 13234 34196
rect 13446 34144 13452 34196
rect 13504 34184 13510 34196
rect 14734 34184 14740 34196
rect 13504 34156 14740 34184
rect 13504 34144 13510 34156
rect 14734 34144 14740 34156
rect 14792 34144 14798 34196
rect 18322 34144 18328 34196
rect 18380 34184 18386 34196
rect 18782 34184 18788 34196
rect 18380 34156 18788 34184
rect 18380 34144 18386 34156
rect 18782 34144 18788 34156
rect 18840 34144 18846 34196
rect 22094 34144 22100 34196
rect 22152 34144 22158 34196
rect 25774 34144 25780 34196
rect 25832 34184 25838 34196
rect 26326 34184 26332 34196
rect 25832 34156 26332 34184
rect 25832 34144 25838 34156
rect 26326 34144 26332 34156
rect 26384 34184 26390 34196
rect 26513 34187 26571 34193
rect 26513 34184 26525 34187
rect 26384 34156 26525 34184
rect 26384 34144 26390 34156
rect 26513 34153 26525 34156
rect 26559 34153 26571 34187
rect 26513 34147 26571 34153
rect 28074 34144 28080 34196
rect 28132 34184 28138 34196
rect 28626 34184 28632 34196
rect 28132 34156 28632 34184
rect 28132 34144 28138 34156
rect 28626 34144 28632 34156
rect 28684 34184 28690 34196
rect 28721 34187 28779 34193
rect 28721 34184 28733 34187
rect 28684 34156 28733 34184
rect 28684 34144 28690 34156
rect 28721 34153 28733 34156
rect 28767 34153 28779 34187
rect 28721 34147 28779 34153
rect 16298 34116 16304 34128
rect 13648 34088 16304 34116
rect 4798 34008 4804 34060
rect 4856 34048 4862 34060
rect 6273 34051 6331 34057
rect 6273 34048 6285 34051
rect 4856 34020 6285 34048
rect 4856 34008 4862 34020
rect 6273 34017 6285 34020
rect 6319 34017 6331 34051
rect 11333 34051 11391 34057
rect 11333 34048 11345 34051
rect 6273 34011 6331 34017
rect 10796 34020 11345 34048
rect 1302 33940 1308 33992
rect 1360 33980 1366 33992
rect 1397 33983 1455 33989
rect 1397 33980 1409 33983
rect 1360 33952 1409 33980
rect 1360 33940 1366 33952
rect 1397 33949 1409 33952
rect 1443 33980 1455 33983
rect 1673 33983 1731 33989
rect 1673 33980 1685 33983
rect 1443 33952 1685 33980
rect 1443 33949 1455 33952
rect 1397 33943 1455 33949
rect 1673 33949 1685 33952
rect 1719 33949 1731 33983
rect 1673 33943 1731 33949
rect 3602 33940 3608 33992
rect 3660 33980 3666 33992
rect 5353 33983 5411 33989
rect 5353 33980 5365 33983
rect 3660 33952 5365 33980
rect 3660 33940 3666 33952
rect 5353 33949 5365 33952
rect 5399 33949 5411 33983
rect 5353 33943 5411 33949
rect 5629 33983 5687 33989
rect 5629 33949 5641 33983
rect 5675 33980 5687 33983
rect 5902 33980 5908 33992
rect 5675 33952 5908 33980
rect 5675 33949 5687 33952
rect 5629 33943 5687 33949
rect 5902 33940 5908 33952
rect 5960 33940 5966 33992
rect 6288 33980 6316 34011
rect 7098 33980 7104 33992
rect 6288 33952 7104 33980
rect 7098 33940 7104 33952
rect 7156 33980 7162 33992
rect 8941 33983 8999 33989
rect 8941 33980 8953 33983
rect 7156 33952 8953 33980
rect 7156 33940 7162 33952
rect 8941 33949 8953 33952
rect 8987 33949 8999 33983
rect 8941 33943 8999 33949
rect 10226 33940 10232 33992
rect 10284 33980 10290 33992
rect 10505 33983 10563 33989
rect 10505 33980 10517 33983
rect 10284 33952 10517 33980
rect 10284 33940 10290 33952
rect 10505 33949 10517 33952
rect 10551 33949 10563 33983
rect 10505 33943 10563 33949
rect 10594 33940 10600 33992
rect 10652 33980 10658 33992
rect 10796 33989 10824 34020
rect 11333 34017 11345 34020
rect 11379 34048 11391 34051
rect 13648 34048 13676 34088
rect 16298 34076 16304 34088
rect 16356 34076 16362 34128
rect 18414 34076 18420 34128
rect 18472 34116 18478 34128
rect 19061 34119 19119 34125
rect 19061 34116 19073 34119
rect 18472 34088 19073 34116
rect 18472 34076 18478 34088
rect 19061 34085 19073 34088
rect 19107 34116 19119 34119
rect 19242 34116 19248 34128
rect 19107 34088 19248 34116
rect 19107 34085 19119 34088
rect 19061 34079 19119 34085
rect 19242 34076 19248 34088
rect 19300 34076 19306 34128
rect 23750 34116 23756 34128
rect 22572 34088 23756 34116
rect 11379 34020 13676 34048
rect 11379 34017 11391 34020
rect 11333 34011 11391 34017
rect 13722 34008 13728 34060
rect 13780 34048 13786 34060
rect 14093 34051 14151 34057
rect 14093 34048 14105 34051
rect 13780 34020 14105 34048
rect 13780 34008 13786 34020
rect 14093 34017 14105 34020
rect 14139 34048 14151 34051
rect 17218 34048 17224 34060
rect 14139 34020 17224 34048
rect 14139 34017 14151 34020
rect 14093 34011 14151 34017
rect 17218 34008 17224 34020
rect 17276 34008 17282 34060
rect 22572 34057 22600 34088
rect 23750 34076 23756 34088
rect 23808 34076 23814 34128
rect 26145 34119 26203 34125
rect 26145 34085 26157 34119
rect 26191 34085 26203 34119
rect 26145 34079 26203 34085
rect 22557 34051 22615 34057
rect 22557 34017 22569 34051
rect 22603 34017 22615 34051
rect 22557 34011 22615 34017
rect 22741 34051 22799 34057
rect 22741 34017 22753 34051
rect 22787 34048 22799 34051
rect 23290 34048 23296 34060
rect 22787 34020 23296 34048
rect 22787 34017 22799 34020
rect 22741 34011 22799 34017
rect 23290 34008 23296 34020
rect 23348 34008 23354 34060
rect 26160 34048 26188 34079
rect 26329 34051 26387 34057
rect 26329 34048 26341 34051
rect 23400 34020 26341 34048
rect 10781 33983 10839 33989
rect 10652 33952 10697 33980
rect 10652 33940 10658 33952
rect 10781 33949 10793 33983
rect 10827 33949 10839 33983
rect 10781 33943 10839 33949
rect 11011 33983 11069 33989
rect 11011 33949 11023 33983
rect 11057 33980 11069 33983
rect 11057 33952 11560 33980
rect 11057 33949 11069 33952
rect 11011 33943 11069 33949
rect 6540 33915 6598 33921
rect 6540 33881 6552 33915
rect 6586 33912 6598 33915
rect 7374 33912 7380 33924
rect 6586 33884 7380 33912
rect 6586 33881 6598 33884
rect 6540 33875 6598 33881
rect 7374 33872 7380 33884
rect 7432 33872 7438 33924
rect 7745 33915 7803 33921
rect 7745 33912 7757 33915
rect 7576 33884 7757 33912
rect 1581 33847 1639 33853
rect 1581 33813 1593 33847
rect 1627 33844 1639 33847
rect 4062 33844 4068 33856
rect 1627 33816 4068 33844
rect 1627 33813 1639 33816
rect 1581 33807 1639 33813
rect 4062 33804 4068 33816
rect 4120 33804 4126 33856
rect 6362 33804 6368 33856
rect 6420 33844 6426 33856
rect 7576 33844 7604 33884
rect 7745 33881 7757 33884
rect 7791 33912 7803 33915
rect 9030 33912 9036 33924
rect 7791 33884 9036 33912
rect 7791 33881 7803 33884
rect 7745 33875 7803 33881
rect 9030 33872 9036 33884
rect 9088 33872 9094 33924
rect 9214 33921 9220 33924
rect 9208 33875 9220 33921
rect 9214 33872 9220 33875
rect 9272 33872 9278 33924
rect 10870 33872 10876 33924
rect 10928 33872 10934 33924
rect 11532 33921 11560 33952
rect 13354 33940 13360 33992
rect 13412 33980 13418 33992
rect 13541 33983 13599 33989
rect 13541 33980 13553 33983
rect 13412 33952 13553 33980
rect 13412 33940 13418 33952
rect 13541 33949 13553 33952
rect 13587 33980 13599 33983
rect 14369 33983 14427 33989
rect 14369 33980 14381 33983
rect 13587 33952 14381 33980
rect 13587 33949 13599 33952
rect 13541 33943 13599 33949
rect 14369 33949 14381 33952
rect 14415 33949 14427 33983
rect 14369 33943 14427 33949
rect 14458 33940 14464 33992
rect 14516 33980 14522 33992
rect 14645 33983 14703 33989
rect 14645 33980 14657 33983
rect 14516 33952 14657 33980
rect 14516 33940 14522 33952
rect 14645 33949 14657 33952
rect 14691 33949 14703 33983
rect 14645 33943 14703 33949
rect 14734 33940 14740 33992
rect 14792 33980 14798 33992
rect 15197 33983 15255 33989
rect 15197 33980 15209 33983
rect 14792 33952 15209 33980
rect 14792 33940 14798 33952
rect 15197 33949 15209 33952
rect 15243 33980 15255 33983
rect 15286 33980 15292 33992
rect 15243 33952 15292 33980
rect 15243 33949 15255 33952
rect 15197 33943 15255 33949
rect 15286 33940 15292 33952
rect 15344 33980 15350 33992
rect 16482 33980 16488 33992
rect 15344 33952 16488 33980
rect 15344 33940 15350 33952
rect 16482 33940 16488 33952
rect 16540 33940 16546 33992
rect 16666 33940 16672 33992
rect 16724 33980 16730 33992
rect 17402 33980 17408 33992
rect 16724 33952 17408 33980
rect 16724 33940 16730 33952
rect 17402 33940 17408 33952
rect 17460 33940 17466 33992
rect 17678 33989 17684 33992
rect 17672 33980 17684 33989
rect 17639 33952 17684 33980
rect 17672 33943 17684 33952
rect 17678 33940 17684 33943
rect 17736 33940 17742 33992
rect 18874 33940 18880 33992
rect 18932 33980 18938 33992
rect 20898 33980 20904 33992
rect 18932 33952 20904 33980
rect 18932 33940 18938 33952
rect 20898 33940 20904 33952
rect 20956 33940 20962 33992
rect 22465 33983 22523 33989
rect 22465 33949 22477 33983
rect 22511 33980 22523 33983
rect 23198 33980 23204 33992
rect 22511 33952 23204 33980
rect 22511 33949 22523 33952
rect 22465 33943 22523 33949
rect 23198 33940 23204 33952
rect 23256 33940 23262 33992
rect 23400 33980 23428 34020
rect 23308 33952 23428 33980
rect 11517 33915 11575 33921
rect 11517 33881 11529 33915
rect 11563 33912 11575 33915
rect 13446 33912 13452 33924
rect 11563 33884 13452 33912
rect 11563 33881 11575 33884
rect 11517 33875 11575 33881
rect 13446 33872 13452 33884
rect 13504 33872 13510 33924
rect 14550 33872 14556 33924
rect 14608 33912 14614 33924
rect 15013 33915 15071 33921
rect 15013 33912 15025 33915
rect 14608 33884 15025 33912
rect 14608 33872 14614 33884
rect 15013 33881 15025 33884
rect 15059 33881 15071 33915
rect 15013 33875 15071 33881
rect 15654 33872 15660 33924
rect 15712 33912 15718 33924
rect 15933 33915 15991 33921
rect 15933 33912 15945 33915
rect 15712 33884 15945 33912
rect 15712 33872 15718 33884
rect 15933 33881 15945 33884
rect 15979 33881 15991 33915
rect 15933 33875 15991 33881
rect 16298 33872 16304 33924
rect 16356 33912 16362 33924
rect 16356 33884 17448 33912
rect 16356 33872 16362 33884
rect 6420 33816 7604 33844
rect 6420 33804 6426 33816
rect 7650 33804 7656 33856
rect 7708 33804 7714 33856
rect 9950 33804 9956 33856
rect 10008 33844 10014 33856
rect 10321 33847 10379 33853
rect 10321 33844 10333 33847
rect 10008 33816 10333 33844
rect 10008 33804 10014 33816
rect 10321 33813 10333 33816
rect 10367 33813 10379 33847
rect 10321 33807 10379 33813
rect 11146 33804 11152 33856
rect 11204 33804 11210 33856
rect 13630 33804 13636 33856
rect 13688 33804 13694 33856
rect 14918 33804 14924 33856
rect 14976 33804 14982 33856
rect 15378 33804 15384 33856
rect 15436 33844 15442 33856
rect 15749 33847 15807 33853
rect 15749 33844 15761 33847
rect 15436 33816 15761 33844
rect 15436 33804 15442 33816
rect 15749 33813 15761 33816
rect 15795 33813 15807 33847
rect 15749 33807 15807 33813
rect 16574 33804 16580 33856
rect 16632 33844 16638 33856
rect 16669 33847 16727 33853
rect 16669 33844 16681 33847
rect 16632 33816 16681 33844
rect 16632 33804 16638 33816
rect 16669 33813 16681 33816
rect 16715 33844 16727 33847
rect 17310 33844 17316 33856
rect 16715 33816 17316 33844
rect 16715 33813 16727 33816
rect 16669 33807 16727 33813
rect 17310 33804 17316 33816
rect 17368 33804 17374 33856
rect 17420 33844 17448 33884
rect 17586 33872 17592 33924
rect 17644 33912 17650 33924
rect 23308 33912 23336 33952
rect 23474 33940 23480 33992
rect 23532 33940 23538 33992
rect 23569 33983 23627 33989
rect 23569 33949 23581 33983
rect 23615 33980 23627 33983
rect 23842 33980 23848 33992
rect 23615 33952 23848 33980
rect 23615 33949 23627 33952
rect 23569 33943 23627 33949
rect 23842 33940 23848 33952
rect 23900 33940 23906 33992
rect 25314 33940 25320 33992
rect 25372 33940 25378 33992
rect 25516 33989 25544 34020
rect 26329 34017 26341 34020
rect 26375 34048 26387 34051
rect 26697 34051 26755 34057
rect 26697 34048 26709 34051
rect 26375 34020 26709 34048
rect 26375 34017 26387 34020
rect 26329 34011 26387 34017
rect 26697 34017 26709 34020
rect 26743 34017 26755 34051
rect 26697 34011 26755 34017
rect 25501 33983 25559 33989
rect 25501 33949 25513 33983
rect 25547 33949 25559 33983
rect 25501 33943 25559 33949
rect 25590 33940 25596 33992
rect 25648 33940 25654 33992
rect 25685 33983 25743 33989
rect 25685 33949 25697 33983
rect 25731 33980 25743 33983
rect 25774 33980 25780 33992
rect 25731 33952 25780 33980
rect 25731 33949 25743 33952
rect 25685 33943 25743 33949
rect 25774 33940 25780 33952
rect 25832 33940 25838 33992
rect 25961 33983 26019 33989
rect 25961 33949 25973 33983
rect 26007 33980 26019 33983
rect 26007 33952 26740 33980
rect 26007 33949 26019 33952
rect 25961 33943 26019 33949
rect 17644 33884 23336 33912
rect 23385 33915 23443 33921
rect 17644 33872 17650 33884
rect 23385 33881 23397 33915
rect 23431 33912 23443 33915
rect 23658 33912 23664 33924
rect 23431 33884 23664 33912
rect 23431 33881 23443 33884
rect 23385 33875 23443 33881
rect 23658 33872 23664 33884
rect 23716 33872 23722 33924
rect 26418 33912 26424 33924
rect 23768 33884 26424 33912
rect 20806 33844 20812 33856
rect 17420 33816 20812 33844
rect 20806 33804 20812 33816
rect 20864 33844 20870 33856
rect 21269 33847 21327 33853
rect 21269 33844 21281 33847
rect 20864 33816 21281 33844
rect 20864 33804 20870 33816
rect 21269 33813 21281 33816
rect 21315 33844 21327 33847
rect 22922 33844 22928 33856
rect 21315 33816 22928 33844
rect 21315 33813 21327 33816
rect 21269 33807 21327 33813
rect 22922 33804 22928 33816
rect 22980 33804 22986 33856
rect 23017 33847 23075 33853
rect 23017 33813 23029 33847
rect 23063 33844 23075 33847
rect 23290 33844 23296 33856
rect 23063 33816 23296 33844
rect 23063 33813 23075 33816
rect 23017 33807 23075 33813
rect 23290 33804 23296 33816
rect 23348 33804 23354 33856
rect 23768 33853 23796 33884
rect 26418 33872 26424 33884
rect 26476 33872 26482 33924
rect 26712 33912 26740 33952
rect 26786 33940 26792 33992
rect 26844 33980 26850 33992
rect 27246 33980 27252 33992
rect 26844 33952 27252 33980
rect 26844 33940 26850 33952
rect 27246 33940 27252 33952
rect 27304 33980 27310 33992
rect 27614 33989 27620 33992
rect 27341 33983 27399 33989
rect 27341 33980 27353 33983
rect 27304 33952 27353 33980
rect 27304 33940 27310 33952
rect 27341 33949 27353 33952
rect 27387 33949 27399 33983
rect 27608 33980 27620 33989
rect 27575 33952 27620 33980
rect 27341 33943 27399 33949
rect 27608 33943 27620 33952
rect 27614 33940 27620 33943
rect 27672 33940 27678 33992
rect 33229 33983 33287 33989
rect 33229 33980 33241 33983
rect 32876 33952 33241 33980
rect 26712 33884 27016 33912
rect 23753 33847 23811 33853
rect 23753 33813 23765 33847
rect 23799 33813 23811 33847
rect 23753 33807 23811 33813
rect 23842 33804 23848 33856
rect 23900 33804 23906 33856
rect 24118 33804 24124 33856
rect 24176 33804 24182 33856
rect 25866 33804 25872 33856
rect 25924 33804 25930 33856
rect 26988 33853 27016 33884
rect 32876 33856 32904 33952
rect 33229 33949 33241 33952
rect 33275 33949 33287 33983
rect 33229 33943 33287 33949
rect 34054 33940 34060 33992
rect 34112 33940 34118 33992
rect 34330 33872 34336 33924
rect 34388 33872 34394 33924
rect 26973 33847 27031 33853
rect 26973 33813 26985 33847
rect 27019 33844 27031 33847
rect 29178 33844 29184 33856
rect 27019 33816 29184 33844
rect 27019 33813 27031 33816
rect 26973 33807 27031 33813
rect 29178 33804 29184 33816
rect 29236 33804 29242 33856
rect 32858 33804 32864 33856
rect 32916 33804 32922 33856
rect 33045 33847 33103 33853
rect 33045 33813 33057 33847
rect 33091 33844 33103 33847
rect 34422 33844 34428 33856
rect 33091 33816 34428 33844
rect 33091 33813 33103 33816
rect 33045 33807 33103 33813
rect 34422 33804 34428 33816
rect 34480 33804 34486 33856
rect 1104 33754 35328 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35328 33754
rect 1104 33680 35328 33702
rect 7374 33600 7380 33652
rect 7432 33600 7438 33652
rect 7650 33600 7656 33652
rect 7708 33640 7714 33652
rect 7745 33643 7803 33649
rect 7745 33640 7757 33643
rect 7708 33612 7757 33640
rect 7708 33600 7714 33612
rect 7745 33609 7757 33612
rect 7791 33609 7803 33643
rect 7745 33603 7803 33609
rect 8849 33643 8907 33649
rect 8849 33609 8861 33643
rect 8895 33640 8907 33643
rect 9214 33640 9220 33652
rect 8895 33612 9220 33640
rect 8895 33609 8907 33612
rect 8849 33603 8907 33609
rect 9214 33600 9220 33612
rect 9272 33600 9278 33652
rect 10226 33600 10232 33652
rect 10284 33600 10290 33652
rect 10413 33643 10471 33649
rect 10413 33609 10425 33643
rect 10459 33640 10471 33643
rect 10502 33640 10508 33652
rect 10459 33612 10508 33640
rect 10459 33609 10471 33612
rect 10413 33603 10471 33609
rect 10502 33600 10508 33612
rect 10560 33600 10566 33652
rect 14550 33640 14556 33652
rect 10704 33612 14556 33640
rect 7098 33532 7104 33584
rect 7156 33532 7162 33584
rect 9232 33544 9812 33572
rect 5068 33507 5126 33513
rect 5068 33473 5080 33507
rect 5114 33504 5126 33507
rect 5442 33504 5448 33516
rect 5114 33476 5448 33504
rect 5114 33473 5126 33476
rect 5068 33467 5126 33473
rect 5442 33464 5448 33476
rect 5500 33464 5506 33516
rect 6362 33464 6368 33516
rect 6420 33464 6426 33516
rect 9232 33513 9260 33544
rect 9217 33507 9275 33513
rect 9217 33473 9229 33507
rect 9263 33473 9275 33507
rect 9217 33467 9275 33473
rect 9674 33464 9680 33516
rect 9732 33464 9738 33516
rect 9784 33504 9812 33544
rect 9858 33532 9864 33584
rect 9916 33532 9922 33584
rect 9950 33532 9956 33584
rect 10008 33532 10014 33584
rect 10704 33572 10732 33612
rect 14550 33600 14556 33612
rect 14608 33640 14614 33652
rect 16298 33640 16304 33652
rect 14608 33612 16304 33640
rect 14608 33600 14614 33612
rect 16298 33600 16304 33612
rect 16356 33600 16362 33652
rect 16485 33643 16543 33649
rect 16485 33609 16497 33643
rect 16531 33609 16543 33643
rect 16485 33603 16543 33609
rect 19521 33643 19579 33649
rect 19521 33609 19533 33643
rect 19567 33640 19579 33643
rect 25774 33640 25780 33652
rect 19567 33612 25780 33640
rect 19567 33609 19579 33612
rect 19521 33603 19579 33609
rect 15381 33575 15439 33581
rect 10520 33544 10732 33572
rect 10796 33544 14412 33572
rect 9784 33476 9895 33504
rect 4798 33396 4804 33448
rect 4856 33396 4862 33448
rect 7834 33396 7840 33448
rect 7892 33396 7898 33448
rect 8021 33439 8079 33445
rect 8021 33405 8033 33439
rect 8067 33436 8079 33439
rect 9309 33439 9367 33445
rect 9309 33436 9321 33439
rect 8067 33408 8340 33436
rect 8067 33405 8079 33408
rect 8021 33399 8079 33405
rect 6178 33260 6184 33312
rect 6236 33260 6242 33312
rect 8312 33309 8340 33408
rect 9232 33408 9321 33436
rect 9232 33380 9260 33408
rect 9309 33405 9321 33408
rect 9355 33405 9367 33439
rect 9309 33399 9367 33405
rect 9493 33439 9551 33445
rect 9493 33405 9505 33439
rect 9539 33436 9551 33439
rect 9766 33436 9772 33448
rect 9539 33408 9772 33436
rect 9539 33405 9551 33408
rect 9493 33399 9551 33405
rect 9766 33396 9772 33408
rect 9824 33396 9830 33448
rect 9214 33328 9220 33380
rect 9272 33328 9278 33380
rect 9867 33368 9895 33476
rect 10042 33464 10048 33516
rect 10100 33464 10106 33516
rect 9950 33368 9956 33380
rect 9867 33340 9956 33368
rect 9950 33328 9956 33340
rect 10008 33328 10014 33380
rect 10042 33328 10048 33380
rect 10100 33368 10106 33380
rect 10520 33377 10548 33544
rect 10505 33371 10563 33377
rect 10505 33368 10517 33371
rect 10100 33340 10517 33368
rect 10100 33328 10106 33340
rect 10505 33337 10517 33340
rect 10551 33337 10563 33371
rect 10505 33331 10563 33337
rect 8297 33303 8355 33309
rect 8297 33269 8309 33303
rect 8343 33300 8355 33303
rect 10796 33300 10824 33544
rect 11790 33513 11796 33516
rect 11784 33467 11796 33513
rect 11790 33464 11796 33467
rect 11848 33464 11854 33516
rect 11514 33396 11520 33448
rect 11572 33396 11578 33448
rect 14384 33368 14412 33544
rect 15381 33541 15393 33575
rect 15427 33572 15439 33575
rect 16022 33572 16028 33584
rect 15427 33544 16028 33572
rect 15427 33541 15439 33544
rect 15381 33535 15439 33541
rect 16022 33532 16028 33544
rect 16080 33532 16086 33584
rect 16114 33532 16120 33584
rect 16172 33532 16178 33584
rect 16500 33572 16528 33603
rect 16914 33575 16972 33581
rect 16914 33572 16926 33575
rect 16500 33544 16926 33572
rect 16914 33541 16926 33544
rect 16960 33541 16972 33575
rect 16914 33535 16972 33541
rect 17034 33532 17040 33584
rect 17092 33572 17098 33584
rect 18509 33575 18567 33581
rect 18509 33572 18521 33575
rect 17092 33544 18521 33572
rect 17092 33532 17098 33544
rect 18509 33541 18521 33544
rect 18555 33572 18567 33575
rect 18969 33575 19027 33581
rect 18969 33572 18981 33575
rect 18555 33544 18981 33572
rect 18555 33541 18567 33544
rect 18509 33535 18567 33541
rect 18969 33541 18981 33544
rect 19015 33541 19027 33575
rect 18969 33535 19027 33541
rect 19058 33532 19064 33584
rect 19116 33532 19122 33584
rect 14918 33464 14924 33516
rect 14976 33504 14982 33516
rect 15013 33507 15071 33513
rect 15013 33504 15025 33507
rect 14976 33476 15025 33504
rect 14976 33464 14982 33476
rect 15013 33473 15025 33476
rect 15059 33473 15071 33507
rect 15013 33467 15071 33473
rect 15102 33464 15108 33516
rect 15160 33504 15166 33516
rect 15289 33507 15347 33513
rect 15160 33476 15205 33504
rect 15160 33464 15166 33476
rect 15289 33473 15301 33507
rect 15335 33473 15347 33507
rect 15289 33467 15347 33473
rect 15519 33507 15577 33513
rect 15519 33473 15531 33507
rect 15565 33504 15577 33507
rect 15654 33504 15660 33516
rect 15565 33476 15660 33504
rect 15565 33473 15577 33476
rect 15519 33467 15577 33473
rect 15304 33436 15332 33467
rect 15654 33464 15660 33476
rect 15712 33464 15718 33516
rect 16592 33476 17724 33504
rect 15378 33436 15384 33448
rect 15304 33408 15384 33436
rect 15378 33396 15384 33408
rect 15436 33396 15442 33448
rect 15933 33439 15991 33445
rect 15933 33405 15945 33439
rect 15979 33405 15991 33439
rect 15933 33399 15991 33405
rect 16025 33439 16083 33445
rect 16025 33405 16037 33439
rect 16071 33436 16083 33439
rect 16592 33436 16620 33476
rect 16071 33408 16620 33436
rect 16071 33405 16083 33408
rect 16025 33399 16083 33405
rect 15838 33368 15844 33380
rect 14384 33340 15844 33368
rect 15838 33328 15844 33340
rect 15896 33328 15902 33380
rect 15948 33368 15976 33399
rect 16666 33396 16672 33448
rect 16724 33396 16730 33448
rect 16574 33368 16580 33380
rect 15948 33340 16580 33368
rect 16574 33328 16580 33340
rect 16632 33328 16638 33380
rect 17696 33368 17724 33476
rect 18690 33464 18696 33516
rect 18748 33464 18754 33516
rect 18782 33464 18788 33516
rect 18840 33504 18846 33516
rect 19199 33507 19257 33513
rect 18840 33476 18885 33504
rect 18840 33464 18846 33476
rect 19199 33473 19211 33507
rect 19245 33504 19257 33507
rect 19536 33504 19564 33603
rect 25774 33600 25780 33612
rect 25832 33600 25838 33652
rect 26973 33643 27031 33649
rect 26973 33609 26985 33643
rect 27019 33609 27031 33643
rect 34333 33643 34391 33649
rect 26973 33603 27031 33609
rect 27080 33612 29592 33640
rect 19610 33532 19616 33584
rect 19668 33572 19674 33584
rect 20625 33575 20683 33581
rect 20625 33572 20637 33575
rect 19668 33544 20637 33572
rect 19668 33532 19674 33544
rect 20625 33541 20637 33544
rect 20671 33572 20683 33575
rect 21821 33575 21879 33581
rect 21821 33572 21833 33575
rect 20671 33544 21833 33572
rect 20671 33541 20683 33544
rect 20625 33535 20683 33541
rect 21821 33541 21833 33544
rect 21867 33572 21879 33575
rect 22002 33572 22008 33584
rect 21867 33544 22008 33572
rect 21867 33541 21879 33544
rect 21821 33535 21879 33541
rect 22002 33532 22008 33544
rect 22060 33532 22066 33584
rect 26544 33575 26602 33581
rect 26544 33541 26556 33575
rect 26590 33572 26602 33575
rect 26988 33572 27016 33603
rect 26590 33544 27016 33572
rect 26590 33541 26602 33544
rect 26544 33535 26602 33541
rect 19245 33476 19564 33504
rect 19245 33473 19257 33476
rect 19199 33467 19257 33473
rect 20438 33464 20444 33516
rect 20496 33464 20502 33516
rect 20714 33464 20720 33516
rect 20772 33464 20778 33516
rect 20806 33464 20812 33516
rect 20864 33464 20870 33516
rect 20990 33464 20996 33516
rect 21048 33504 21054 33516
rect 21085 33507 21143 33513
rect 21085 33504 21097 33507
rect 21048 33476 21097 33504
rect 21048 33464 21054 33476
rect 21085 33473 21097 33476
rect 21131 33473 21143 33507
rect 21361 33507 21419 33513
rect 21361 33504 21373 33507
rect 21085 33467 21143 33473
rect 21284 33476 21373 33504
rect 21177 33439 21235 33445
rect 21177 33436 21189 33439
rect 19352 33408 21189 33436
rect 17770 33368 17776 33380
rect 17696 33340 17776 33368
rect 17770 33328 17776 33340
rect 17828 33368 17834 33380
rect 19352 33377 19380 33408
rect 21177 33405 21189 33408
rect 21223 33405 21235 33439
rect 21177 33399 21235 33405
rect 18049 33371 18107 33377
rect 18049 33368 18061 33371
rect 17828 33340 18061 33368
rect 17828 33328 17834 33340
rect 18049 33337 18061 33340
rect 18095 33337 18107 33371
rect 18049 33331 18107 33337
rect 19337 33371 19395 33377
rect 19337 33337 19349 33371
rect 19383 33337 19395 33371
rect 19337 33331 19395 33337
rect 20993 33371 21051 33377
rect 20993 33337 21005 33371
rect 21039 33368 21051 33371
rect 21284 33368 21312 33476
rect 21361 33473 21373 33476
rect 21407 33473 21419 33507
rect 21361 33467 21419 33473
rect 23017 33507 23075 33513
rect 23017 33473 23029 33507
rect 23063 33504 23075 33507
rect 23106 33504 23112 33516
rect 23063 33476 23112 33504
rect 23063 33473 23075 33476
rect 23017 33467 23075 33473
rect 23106 33464 23112 33476
rect 23164 33464 23170 33516
rect 27080 33504 27108 33612
rect 27433 33575 27491 33581
rect 27433 33541 27445 33575
rect 27479 33572 27491 33575
rect 27522 33572 27528 33584
rect 27479 33544 27528 33572
rect 27479 33541 27491 33544
rect 27433 33535 27491 33541
rect 27522 33532 27528 33544
rect 27580 33532 27586 33584
rect 28626 33532 28632 33584
rect 28684 33532 28690 33584
rect 25792 33476 27108 33504
rect 27341 33507 27399 33513
rect 22281 33439 22339 33445
rect 22281 33405 22293 33439
rect 22327 33436 22339 33439
rect 22554 33436 22560 33448
rect 22327 33408 22560 33436
rect 22327 33405 22339 33408
rect 22281 33399 22339 33405
rect 22554 33396 22560 33408
rect 22612 33396 22618 33448
rect 21039 33340 21312 33368
rect 21545 33371 21603 33377
rect 21039 33337 21051 33340
rect 20993 33331 21051 33337
rect 21545 33337 21557 33371
rect 21591 33368 21603 33371
rect 25792 33368 25820 33476
rect 27341 33473 27353 33507
rect 27387 33473 27399 33507
rect 27341 33467 27399 33473
rect 26786 33396 26792 33448
rect 26844 33396 26850 33448
rect 21591 33340 25820 33368
rect 21591 33337 21603 33340
rect 21545 33331 21603 33337
rect 8343 33272 10824 33300
rect 8343 33269 8355 33272
rect 8297 33263 8355 33269
rect 12158 33260 12164 33312
rect 12216 33300 12222 33312
rect 12897 33303 12955 33309
rect 12897 33300 12909 33303
rect 12216 33272 12909 33300
rect 12216 33260 12222 33272
rect 12897 33269 12909 33272
rect 12943 33269 12955 33303
rect 12897 33263 12955 33269
rect 15657 33303 15715 33309
rect 15657 33269 15669 33303
rect 15703 33300 15715 33303
rect 17402 33300 17408 33312
rect 15703 33272 17408 33300
rect 15703 33269 15715 33272
rect 15657 33263 15715 33269
rect 17402 33260 17408 33272
rect 17460 33260 17466 33312
rect 21082 33260 21088 33312
rect 21140 33260 21146 33312
rect 23106 33260 23112 33312
rect 23164 33260 23170 33312
rect 25409 33303 25467 33309
rect 25409 33269 25421 33303
rect 25455 33300 25467 33303
rect 26602 33300 26608 33312
rect 25455 33272 26608 33300
rect 25455 33269 25467 33272
rect 25409 33263 25467 33269
rect 26602 33260 26608 33272
rect 26660 33300 26666 33312
rect 27356 33300 27384 33467
rect 28258 33464 28264 33516
rect 28316 33464 28322 33516
rect 28442 33513 28448 33516
rect 28409 33507 28448 33513
rect 28409 33473 28421 33507
rect 28409 33467 28448 33473
rect 28442 33464 28448 33467
rect 28500 33464 28506 33516
rect 28537 33507 28595 33513
rect 28537 33473 28549 33507
rect 28583 33504 28595 33507
rect 28583 33476 28672 33504
rect 28583 33473 28595 33476
rect 28537 33467 28595 33473
rect 27617 33439 27675 33445
rect 27617 33405 27629 33439
rect 27663 33436 27675 33439
rect 27706 33436 27712 33448
rect 27663 33408 27712 33436
rect 27663 33405 27675 33408
rect 27617 33399 27675 33405
rect 27706 33396 27712 33408
rect 27764 33396 27770 33448
rect 26660 33272 27384 33300
rect 28644 33300 28672 33476
rect 28718 33464 28724 33516
rect 28776 33513 28782 33516
rect 28776 33504 28784 33513
rect 28776 33476 28821 33504
rect 28776 33467 28784 33476
rect 28776 33464 28782 33467
rect 29270 33464 29276 33516
rect 29328 33464 29334 33516
rect 29564 33513 29592 33612
rect 34333 33609 34345 33643
rect 34379 33640 34391 33643
rect 34514 33640 34520 33652
rect 34379 33612 34520 33640
rect 34379 33609 34391 33612
rect 34333 33603 34391 33609
rect 34514 33600 34520 33612
rect 34572 33600 34578 33652
rect 29457 33507 29515 33513
rect 29457 33473 29469 33507
rect 29503 33473 29515 33507
rect 29457 33467 29515 33473
rect 29549 33507 29607 33513
rect 29549 33473 29561 33507
rect 29595 33473 29607 33507
rect 29549 33467 29607 33473
rect 29472 33436 29500 33467
rect 29822 33464 29828 33516
rect 29880 33464 29886 33516
rect 33502 33464 33508 33516
rect 33560 33464 33566 33516
rect 34146 33464 34152 33516
rect 34204 33464 34210 33516
rect 34422 33464 34428 33516
rect 34480 33464 34486 33516
rect 28920 33408 29500 33436
rect 29641 33439 29699 33445
rect 28920 33377 28948 33408
rect 29641 33405 29653 33439
rect 29687 33436 29699 33439
rect 30101 33439 30159 33445
rect 30101 33436 30113 33439
rect 29687 33408 30113 33436
rect 29687 33405 29699 33408
rect 29641 33399 29699 33405
rect 30101 33405 30113 33408
rect 30147 33405 30159 33439
rect 30101 33399 30159 33405
rect 28905 33371 28963 33377
rect 28905 33337 28917 33371
rect 28951 33337 28963 33371
rect 28905 33331 28963 33337
rect 29546 33328 29552 33380
rect 29604 33368 29610 33380
rect 29656 33368 29684 33399
rect 32122 33396 32128 33448
rect 32180 33396 32186 33448
rect 32398 33396 32404 33448
rect 32456 33396 32462 33448
rect 29604 33340 29684 33368
rect 30009 33371 30067 33377
rect 29604 33328 29610 33340
rect 30009 33337 30021 33371
rect 30055 33368 30067 33371
rect 31018 33368 31024 33380
rect 30055 33340 31024 33368
rect 30055 33337 30067 33340
rect 30009 33331 30067 33337
rect 31018 33328 31024 33340
rect 31076 33328 31082 33380
rect 33410 33328 33416 33380
rect 33468 33368 33474 33380
rect 33965 33371 34023 33377
rect 33965 33368 33977 33371
rect 33468 33340 33977 33368
rect 33468 33328 33474 33340
rect 33965 33337 33977 33340
rect 34011 33337 34023 33371
rect 33965 33331 34023 33337
rect 29089 33303 29147 33309
rect 29089 33300 29101 33303
rect 28644 33272 29101 33300
rect 26660 33260 26666 33272
rect 29089 33269 29101 33272
rect 29135 33300 29147 33303
rect 29178 33300 29184 33312
rect 29135 33272 29184 33300
rect 29135 33269 29147 33272
rect 29089 33263 29147 33269
rect 29178 33260 29184 33272
rect 29236 33260 29242 33312
rect 33134 33260 33140 33312
rect 33192 33300 33198 33312
rect 33873 33303 33931 33309
rect 33873 33300 33885 33303
rect 33192 33272 33885 33300
rect 33192 33260 33198 33272
rect 33873 33269 33885 33272
rect 33919 33300 33931 33303
rect 34054 33300 34060 33312
rect 33919 33272 34060 33300
rect 33919 33269 33931 33272
rect 33873 33263 33931 33269
rect 34054 33260 34060 33272
rect 34112 33260 34118 33312
rect 1104 33210 35328 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 35328 33210
rect 1104 33136 35328 33158
rect 5442 33056 5448 33108
rect 5500 33056 5506 33108
rect 9582 33056 9588 33108
rect 9640 33096 9646 33108
rect 10045 33099 10103 33105
rect 10045 33096 10057 33099
rect 9640 33068 10057 33096
rect 9640 33056 9646 33068
rect 10045 33065 10057 33068
rect 10091 33065 10103 33099
rect 10045 33059 10103 33065
rect 11701 33099 11759 33105
rect 11701 33065 11713 33099
rect 11747 33096 11759 33099
rect 11790 33096 11796 33108
rect 11747 33068 11796 33096
rect 11747 33065 11759 33068
rect 11701 33059 11759 33065
rect 11790 33056 11796 33068
rect 11848 33056 11854 33108
rect 14090 33056 14096 33108
rect 14148 33096 14154 33108
rect 17957 33099 18015 33105
rect 14148 33068 15792 33096
rect 14148 33056 14154 33068
rect 8021 33031 8079 33037
rect 8021 32997 8033 33031
rect 8067 33028 8079 33031
rect 10413 33031 10471 33037
rect 8067 33000 10180 33028
rect 8067 32997 8079 33000
rect 8021 32991 8079 32997
rect 6089 32963 6147 32969
rect 6089 32929 6101 32963
rect 6135 32960 6147 32963
rect 7006 32960 7012 32972
rect 6135 32932 7012 32960
rect 6135 32929 6147 32932
rect 6089 32923 6147 32929
rect 7006 32920 7012 32932
rect 7064 32920 7070 32972
rect 7650 32920 7656 32972
rect 7708 32920 7714 32972
rect 7742 32920 7748 32972
rect 7800 32960 7806 32972
rect 8113 32963 8171 32969
rect 8113 32960 8125 32963
rect 7800 32932 8125 32960
rect 7800 32920 7806 32932
rect 8113 32929 8125 32932
rect 8159 32929 8171 32963
rect 8113 32923 8171 32929
rect 9766 32920 9772 32972
rect 9824 32960 9830 32972
rect 9950 32960 9956 32972
rect 9824 32932 9956 32960
rect 9824 32920 9830 32932
rect 9950 32920 9956 32932
rect 10008 32920 10014 32972
rect 10152 32969 10180 33000
rect 10413 32997 10425 33031
rect 10459 33028 10471 33031
rect 10459 33000 14044 33028
rect 10459 32997 10471 33000
rect 10413 32991 10471 32997
rect 10137 32963 10195 32969
rect 10137 32929 10149 32963
rect 10183 32929 10195 32963
rect 10137 32923 10195 32929
rect 12345 32963 12403 32969
rect 12345 32929 12357 32963
rect 12391 32960 12403 32963
rect 13357 32963 13415 32969
rect 13357 32960 13369 32963
rect 12391 32932 12848 32960
rect 12391 32929 12403 32932
rect 12345 32923 12403 32929
rect 4798 32852 4804 32904
rect 4856 32892 4862 32904
rect 6273 32895 6331 32901
rect 6273 32892 6285 32895
rect 4856 32864 6285 32892
rect 4856 32852 4862 32864
rect 6273 32861 6285 32864
rect 6319 32861 6331 32895
rect 6273 32855 6331 32861
rect 7374 32852 7380 32904
rect 7432 32852 7438 32904
rect 7525 32895 7583 32901
rect 7525 32861 7537 32895
rect 7571 32892 7583 32895
rect 7668 32892 7696 32920
rect 7571 32864 7696 32892
rect 7883 32895 7941 32901
rect 7571 32861 7583 32864
rect 7525 32855 7583 32861
rect 7883 32861 7895 32895
rect 7929 32892 7941 32895
rect 10045 32895 10103 32901
rect 7929 32864 8432 32892
rect 7929 32861 7941 32864
rect 7883 32855 7941 32861
rect 5813 32827 5871 32833
rect 5813 32793 5825 32827
rect 5859 32824 5871 32827
rect 6178 32824 6184 32836
rect 5859 32796 6184 32824
rect 5859 32793 5871 32796
rect 5813 32787 5871 32793
rect 6178 32784 6184 32796
rect 6236 32824 6242 32836
rect 6236 32796 7144 32824
rect 6236 32784 6242 32796
rect 5902 32716 5908 32768
rect 5960 32716 5966 32768
rect 7006 32716 7012 32768
rect 7064 32716 7070 32768
rect 7116 32756 7144 32796
rect 7650 32784 7656 32836
rect 7708 32784 7714 32836
rect 8404 32833 8432 32864
rect 10045 32861 10057 32895
rect 10091 32861 10103 32895
rect 10045 32855 10103 32861
rect 7745 32827 7803 32833
rect 7745 32793 7757 32827
rect 7791 32793 7803 32827
rect 7745 32787 7803 32793
rect 8389 32827 8447 32833
rect 8389 32793 8401 32827
rect 8435 32824 8447 32827
rect 9766 32824 9772 32836
rect 8435 32796 9772 32824
rect 8435 32793 8447 32796
rect 8389 32787 8447 32793
rect 7760 32756 7788 32787
rect 9766 32784 9772 32796
rect 9824 32784 9830 32836
rect 10060 32824 10088 32855
rect 10502 32852 10508 32904
rect 10560 32852 10566 32904
rect 11790 32852 11796 32904
rect 11848 32892 11854 32904
rect 12158 32892 12164 32904
rect 11848 32864 12164 32892
rect 11848 32852 11854 32864
rect 12158 32852 12164 32864
rect 12216 32852 12222 32904
rect 12713 32895 12771 32901
rect 12713 32892 12725 32895
rect 12406 32864 12725 32892
rect 12406 32824 12434 32864
rect 12713 32861 12725 32864
rect 12759 32861 12771 32895
rect 12713 32855 12771 32861
rect 10060 32796 12434 32824
rect 7116 32728 7788 32756
rect 7834 32716 7840 32768
rect 7892 32756 7898 32768
rect 11882 32756 11888 32768
rect 7892 32728 11888 32756
rect 7892 32716 7898 32728
rect 11882 32716 11888 32728
rect 11940 32716 11946 32768
rect 12066 32716 12072 32768
rect 12124 32716 12130 32768
rect 12621 32759 12679 32765
rect 12621 32725 12633 32759
rect 12667 32756 12679 32759
rect 12820 32756 12848 32932
rect 12912 32932 13369 32960
rect 12912 32901 12940 32932
rect 13357 32929 13369 32932
rect 13403 32960 13415 32963
rect 13906 32960 13912 32972
rect 13403 32932 13912 32960
rect 13403 32929 13415 32932
rect 13357 32923 13415 32929
rect 13906 32920 13912 32932
rect 13964 32920 13970 32972
rect 12897 32895 12955 32901
rect 12897 32861 12909 32895
rect 12943 32861 12955 32895
rect 12897 32855 12955 32861
rect 12986 32852 12992 32904
rect 13044 32852 13050 32904
rect 13170 32852 13176 32904
rect 13228 32852 13234 32904
rect 13265 32895 13323 32901
rect 13265 32861 13277 32895
rect 13311 32892 13323 32895
rect 13311 32864 13584 32892
rect 13311 32861 13323 32864
rect 13265 32855 13323 32861
rect 13556 32768 13584 32864
rect 13354 32756 13360 32768
rect 12667 32728 13360 32756
rect 12667 32725 12679 32728
rect 12621 32719 12679 32725
rect 13354 32716 13360 32728
rect 13412 32716 13418 32768
rect 13538 32716 13544 32768
rect 13596 32716 13602 32768
rect 14016 32756 14044 33000
rect 14090 32920 14096 32972
rect 14148 32920 14154 32972
rect 14182 32852 14188 32904
rect 14240 32892 14246 32904
rect 15657 32895 15715 32901
rect 15657 32892 15669 32895
rect 14240 32864 15669 32892
rect 14240 32852 14246 32864
rect 15657 32861 15669 32864
rect 15703 32861 15715 32895
rect 15764 32892 15792 33068
rect 17957 33065 17969 33099
rect 18003 33096 18015 33099
rect 28350 33096 28356 33108
rect 18003 33068 28356 33096
rect 18003 33065 18015 33068
rect 17957 33059 18015 33065
rect 28350 33056 28356 33068
rect 28408 33056 28414 33108
rect 29822 33056 29828 33108
rect 29880 33096 29886 33108
rect 30929 33099 30987 33105
rect 30929 33096 30941 33099
rect 29880 33068 30941 33096
rect 29880 33056 29886 33068
rect 30929 33065 30941 33068
rect 30975 33065 30987 33099
rect 30929 33059 30987 33065
rect 32217 33099 32275 33105
rect 32217 33065 32229 33099
rect 32263 33096 32275 33099
rect 32398 33096 32404 33108
rect 32263 33068 32404 33096
rect 32263 33065 32275 33068
rect 32217 33059 32275 33065
rect 32398 33056 32404 33068
rect 32456 33056 32462 33108
rect 34514 33056 34520 33108
rect 34572 33056 34578 33108
rect 23750 32988 23756 33040
rect 23808 32988 23814 33040
rect 26881 33031 26939 33037
rect 26881 33028 26893 33031
rect 26160 33000 26893 33028
rect 18049 32963 18107 32969
rect 18049 32960 18061 32963
rect 17236 32932 18061 32960
rect 15841 32895 15899 32901
rect 15841 32892 15853 32895
rect 15764 32864 15853 32892
rect 15657 32855 15715 32861
rect 15841 32861 15853 32864
rect 15887 32892 15899 32895
rect 16666 32892 16672 32904
rect 15887 32864 16672 32892
rect 15887 32861 15899 32864
rect 15841 32855 15899 32861
rect 14360 32827 14418 32833
rect 14360 32793 14372 32827
rect 14406 32824 14418 32827
rect 14458 32824 14464 32836
rect 14406 32796 14464 32824
rect 14406 32793 14418 32796
rect 14360 32787 14418 32793
rect 14458 32784 14464 32796
rect 14516 32784 14522 32836
rect 15672 32824 15700 32855
rect 16666 32852 16672 32864
rect 16724 32892 16730 32904
rect 17236 32901 17264 32932
rect 18049 32929 18061 32932
rect 18095 32929 18107 32963
rect 18049 32923 18107 32929
rect 22094 32920 22100 32972
rect 22152 32960 22158 32972
rect 26160 32960 26188 33000
rect 26881 32997 26893 33000
rect 26927 33028 26939 33031
rect 27157 33031 27215 33037
rect 27157 33028 27169 33031
rect 26927 33000 27169 33028
rect 26927 32997 26939 33000
rect 26881 32991 26939 32997
rect 27157 32997 27169 33000
rect 27203 33028 27215 33031
rect 27433 33031 27491 33037
rect 27433 33028 27445 33031
rect 27203 33000 27445 33028
rect 27203 32997 27215 33000
rect 27157 32991 27215 32997
rect 27433 32997 27445 33000
rect 27479 32997 27491 33031
rect 27433 32991 27491 32997
rect 32766 32960 32772 32972
rect 22152 32932 24532 32960
rect 22152 32920 22158 32932
rect 16945 32895 17003 32901
rect 16945 32892 16957 32895
rect 16724 32864 16957 32892
rect 16724 32852 16730 32864
rect 16945 32861 16957 32864
rect 16991 32861 17003 32895
rect 16945 32855 17003 32861
rect 17221 32895 17279 32901
rect 17221 32861 17233 32895
rect 17267 32861 17279 32895
rect 17221 32855 17279 32861
rect 16209 32827 16267 32833
rect 16209 32824 16221 32827
rect 14568 32796 15599 32824
rect 15672 32796 16221 32824
rect 14568 32756 14596 32796
rect 14016 32728 14596 32756
rect 14826 32716 14832 32768
rect 14884 32756 14890 32768
rect 15102 32756 15108 32768
rect 14884 32728 15108 32756
rect 14884 32716 14890 32728
rect 15102 32716 15108 32728
rect 15160 32756 15166 32768
rect 15473 32759 15531 32765
rect 15473 32756 15485 32759
rect 15160 32728 15485 32756
rect 15160 32716 15166 32728
rect 15473 32725 15485 32728
rect 15519 32725 15531 32759
rect 15571 32756 15599 32796
rect 16209 32793 16221 32796
rect 16255 32793 16267 32827
rect 16209 32787 16267 32793
rect 16758 32784 16764 32836
rect 16816 32824 16822 32836
rect 17236 32824 17264 32855
rect 17402 32852 17408 32904
rect 17460 32852 17466 32904
rect 17497 32895 17555 32901
rect 17497 32861 17509 32895
rect 17543 32861 17555 32895
rect 17497 32855 17555 32861
rect 17589 32895 17647 32901
rect 17589 32861 17601 32895
rect 17635 32861 17647 32895
rect 17589 32855 17647 32861
rect 16816 32796 17264 32824
rect 16816 32784 16822 32796
rect 17512 32756 17540 32855
rect 15571 32728 17540 32756
rect 17604 32756 17632 32855
rect 17770 32852 17776 32904
rect 17828 32852 17834 32904
rect 18598 32852 18604 32904
rect 18656 32892 18662 32904
rect 19245 32895 19303 32901
rect 19245 32892 19257 32895
rect 18656 32864 19257 32892
rect 18656 32852 18662 32864
rect 19245 32861 19257 32864
rect 19291 32892 19303 32895
rect 21085 32895 21143 32901
rect 21085 32892 21097 32895
rect 19291 32864 21097 32892
rect 19291 32861 19303 32864
rect 19245 32855 19303 32861
rect 21085 32861 21097 32864
rect 21131 32892 21143 32895
rect 21131 32864 22094 32892
rect 21131 32861 21143 32864
rect 21085 32855 21143 32861
rect 19512 32827 19570 32833
rect 19512 32793 19524 32827
rect 19558 32824 19570 32827
rect 19610 32824 19616 32836
rect 19558 32796 19616 32824
rect 19558 32793 19570 32796
rect 19512 32787 19570 32793
rect 19610 32784 19616 32796
rect 19668 32784 19674 32836
rect 21174 32824 21180 32836
rect 19720 32796 21180 32824
rect 17678 32756 17684 32768
rect 17604 32728 17684 32756
rect 15473 32719 15531 32725
rect 17678 32716 17684 32728
rect 17736 32756 17742 32768
rect 18325 32759 18383 32765
rect 18325 32756 18337 32759
rect 17736 32728 18337 32756
rect 17736 32716 17742 32728
rect 18325 32725 18337 32728
rect 18371 32756 18383 32759
rect 19720 32756 19748 32796
rect 21174 32784 21180 32796
rect 21232 32784 21238 32836
rect 21352 32827 21410 32833
rect 21352 32793 21364 32827
rect 21398 32824 21410 32827
rect 21450 32824 21456 32836
rect 21398 32796 21456 32824
rect 21398 32793 21410 32796
rect 21352 32787 21410 32793
rect 21450 32784 21456 32796
rect 21508 32784 21514 32836
rect 22066 32824 22094 32864
rect 23566 32852 23572 32904
rect 23624 32852 23630 32904
rect 24394 32852 24400 32904
rect 24452 32852 24458 32904
rect 24504 32892 24532 32932
rect 25792 32932 26188 32960
rect 25792 32892 25820 32932
rect 24504 32864 25820 32892
rect 25866 32852 25872 32904
rect 25924 32852 25930 32904
rect 26160 32901 26188 32932
rect 32140 32932 32772 32960
rect 32140 32904 32168 32932
rect 32766 32920 32772 32932
rect 32824 32920 32830 32972
rect 33045 32963 33103 32969
rect 33045 32929 33057 32963
rect 33091 32960 33103 32963
rect 33410 32960 33416 32972
rect 33091 32932 33416 32960
rect 33091 32929 33103 32932
rect 33045 32923 33103 32929
rect 33410 32920 33416 32932
rect 33468 32920 33474 32972
rect 25962 32895 26020 32901
rect 25962 32861 25974 32895
rect 26008 32861 26020 32895
rect 25962 32855 26020 32861
rect 26145 32895 26203 32901
rect 26145 32861 26157 32895
rect 26191 32861 26203 32895
rect 26145 32855 26203 32861
rect 26375 32895 26433 32901
rect 26375 32861 26387 32895
rect 26421 32892 26433 32895
rect 28718 32892 28724 32904
rect 26421 32864 28724 32892
rect 26421 32861 26433 32864
rect 26375 32855 26433 32861
rect 22554 32824 22560 32836
rect 22066 32796 22560 32824
rect 22554 32784 22560 32796
rect 22612 32824 22618 32836
rect 24412 32824 24440 32852
rect 22612 32796 24440 32824
rect 22612 32784 22618 32796
rect 24486 32784 24492 32836
rect 24544 32824 24550 32836
rect 24642 32827 24700 32833
rect 24642 32824 24654 32827
rect 24544 32796 24654 32824
rect 24544 32784 24550 32796
rect 24642 32793 24654 32796
rect 24688 32793 24700 32827
rect 25976 32824 26004 32855
rect 28718 32852 28724 32864
rect 28776 32852 28782 32904
rect 29549 32895 29607 32901
rect 29549 32861 29561 32895
rect 29595 32892 29607 32895
rect 29638 32892 29644 32904
rect 29595 32864 29644 32892
rect 29595 32861 29607 32864
rect 29549 32855 29607 32861
rect 29638 32852 29644 32864
rect 29696 32892 29702 32904
rect 32122 32892 32128 32904
rect 29696 32864 32128 32892
rect 29696 32852 29702 32864
rect 32122 32852 32128 32864
rect 32180 32852 32186 32904
rect 32401 32895 32459 32901
rect 32401 32861 32413 32895
rect 32447 32861 32459 32895
rect 32677 32895 32735 32901
rect 32677 32892 32689 32895
rect 32401 32855 32459 32861
rect 32508 32864 32689 32892
rect 24642 32787 24700 32793
rect 25792 32796 26004 32824
rect 26237 32827 26295 32833
rect 25792 32768 25820 32796
rect 26237 32793 26249 32827
rect 26283 32824 26295 32827
rect 26602 32824 26608 32836
rect 26283 32796 26608 32824
rect 26283 32793 26295 32796
rect 26237 32787 26295 32793
rect 26602 32784 26608 32796
rect 26660 32784 26666 32836
rect 26697 32827 26755 32833
rect 26697 32793 26709 32827
rect 26743 32824 26755 32827
rect 26743 32796 27016 32824
rect 26743 32793 26755 32796
rect 26697 32787 26755 32793
rect 26988 32768 27016 32796
rect 28166 32784 28172 32836
rect 28224 32824 28230 32836
rect 29822 32833 29828 32836
rect 28813 32827 28871 32833
rect 28813 32824 28825 32827
rect 28224 32796 28825 32824
rect 28224 32784 28230 32796
rect 28813 32793 28825 32796
rect 28859 32793 28871 32827
rect 28813 32787 28871 32793
rect 29816 32787 29828 32833
rect 29822 32784 29828 32787
rect 29880 32784 29886 32836
rect 31018 32784 31024 32836
rect 31076 32824 31082 32836
rect 32416 32824 32444 32855
rect 31076 32796 32444 32824
rect 31076 32784 31082 32796
rect 18371 32728 19748 32756
rect 18371 32725 18383 32728
rect 18325 32719 18383 32725
rect 19978 32716 19984 32768
rect 20036 32756 20042 32768
rect 20438 32756 20444 32768
rect 20036 32728 20444 32756
rect 20036 32716 20042 32728
rect 20438 32716 20444 32728
rect 20496 32756 20502 32768
rect 20625 32759 20683 32765
rect 20625 32756 20637 32759
rect 20496 32728 20637 32756
rect 20496 32716 20502 32728
rect 20625 32725 20637 32728
rect 20671 32725 20683 32759
rect 20625 32719 20683 32725
rect 21266 32716 21272 32768
rect 21324 32756 21330 32768
rect 22465 32759 22523 32765
rect 22465 32756 22477 32759
rect 21324 32728 22477 32756
rect 21324 32716 21330 32728
rect 22465 32725 22477 32728
rect 22511 32725 22523 32759
rect 22465 32719 22523 32725
rect 25774 32716 25780 32768
rect 25832 32716 25838 32768
rect 26050 32716 26056 32768
rect 26108 32756 26114 32768
rect 26513 32759 26571 32765
rect 26513 32756 26525 32759
rect 26108 32728 26525 32756
rect 26108 32716 26114 32728
rect 26513 32725 26525 32728
rect 26559 32725 26571 32759
rect 26513 32719 26571 32725
rect 26970 32716 26976 32768
rect 27028 32716 27034 32768
rect 28626 32716 28632 32768
rect 28684 32716 28690 32768
rect 32508 32756 32536 32864
rect 32677 32861 32689 32864
rect 32723 32861 32735 32895
rect 32677 32855 32735 32861
rect 32585 32827 32643 32833
rect 32585 32793 32597 32827
rect 32631 32824 32643 32827
rect 33134 32824 33140 32836
rect 32631 32796 33140 32824
rect 32631 32793 32643 32796
rect 32585 32787 32643 32793
rect 33134 32784 33140 32796
rect 33192 32784 33198 32836
rect 33502 32784 33508 32836
rect 33560 32784 33566 32836
rect 34422 32756 34428 32768
rect 32508 32728 34428 32756
rect 34422 32716 34428 32728
rect 34480 32716 34486 32768
rect 1104 32666 35328 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35328 32666
rect 1104 32592 35328 32614
rect 7834 32552 7840 32564
rect 7668 32524 7840 32552
rect 4798 32484 4804 32496
rect 3436 32456 4804 32484
rect 3436 32360 3464 32456
rect 4798 32444 4804 32456
rect 4856 32444 4862 32496
rect 3688 32419 3746 32425
rect 3688 32385 3700 32419
rect 3734 32416 3746 32419
rect 3970 32416 3976 32428
rect 3734 32388 3976 32416
rect 3734 32385 3746 32388
rect 3688 32379 3746 32385
rect 3970 32376 3976 32388
rect 4028 32376 4034 32428
rect 5902 32376 5908 32428
rect 5960 32416 5966 32428
rect 6365 32419 6423 32425
rect 6365 32416 6377 32419
rect 5960 32388 6377 32416
rect 5960 32376 5966 32388
rect 6365 32385 6377 32388
rect 6411 32416 6423 32419
rect 7668 32416 7696 32524
rect 7834 32512 7840 32524
rect 7892 32512 7898 32564
rect 9122 32512 9128 32564
rect 9180 32552 9186 32564
rect 9585 32555 9643 32561
rect 9585 32552 9597 32555
rect 9180 32524 9597 32552
rect 9180 32512 9186 32524
rect 9585 32521 9597 32524
rect 9631 32521 9643 32555
rect 9585 32515 9643 32521
rect 9766 32512 9772 32564
rect 9824 32552 9830 32564
rect 10778 32552 10784 32564
rect 9824 32524 10784 32552
rect 9824 32512 9830 32524
rect 10778 32512 10784 32524
rect 10836 32512 10842 32564
rect 12986 32512 12992 32564
rect 13044 32552 13050 32564
rect 13725 32555 13783 32561
rect 13725 32552 13737 32555
rect 13044 32524 13737 32552
rect 13044 32512 13050 32524
rect 13725 32521 13737 32524
rect 13771 32521 13783 32555
rect 13725 32515 13783 32521
rect 13906 32512 13912 32564
rect 13964 32552 13970 32564
rect 14366 32552 14372 32564
rect 13964 32524 14372 32552
rect 13964 32512 13970 32524
rect 14366 32512 14372 32524
rect 14424 32512 14430 32564
rect 14458 32512 14464 32564
rect 14516 32512 14522 32564
rect 14826 32512 14832 32564
rect 14884 32512 14890 32564
rect 16206 32552 16212 32564
rect 14936 32524 16212 32552
rect 8202 32484 8208 32496
rect 7760 32456 8208 32484
rect 7760 32425 7788 32456
rect 8202 32444 8208 32456
rect 8260 32444 8266 32496
rect 9030 32444 9036 32496
rect 9088 32484 9094 32496
rect 10137 32487 10195 32493
rect 10137 32484 10149 32487
rect 9088 32456 10149 32484
rect 9088 32444 9094 32456
rect 10137 32453 10149 32456
rect 10183 32484 10195 32487
rect 11149 32487 11207 32493
rect 11149 32484 11161 32487
rect 10183 32456 11161 32484
rect 10183 32453 10195 32456
rect 10137 32447 10195 32453
rect 11149 32453 11161 32456
rect 11195 32484 11207 32487
rect 12710 32484 12716 32496
rect 11195 32456 12716 32484
rect 11195 32453 11207 32456
rect 11149 32447 11207 32453
rect 12710 32444 12716 32456
rect 12768 32444 12774 32496
rect 12894 32444 12900 32496
rect 12952 32484 12958 32496
rect 14182 32484 14188 32496
rect 12952 32456 14188 32484
rect 12952 32444 12958 32456
rect 14182 32444 14188 32456
rect 14240 32444 14246 32496
rect 14936 32484 14964 32524
rect 16206 32512 16212 32524
rect 16264 32512 16270 32564
rect 16574 32512 16580 32564
rect 16632 32552 16638 32564
rect 19518 32552 19524 32564
rect 16632 32524 19524 32552
rect 16632 32512 16638 32524
rect 19518 32512 19524 32524
rect 19576 32512 19582 32564
rect 19610 32512 19616 32564
rect 19668 32512 19674 32564
rect 19978 32512 19984 32564
rect 20036 32512 20042 32564
rect 20990 32512 20996 32564
rect 21048 32512 21054 32564
rect 21174 32512 21180 32564
rect 21232 32552 21238 32564
rect 24765 32555 24823 32561
rect 21232 32524 24716 32552
rect 21232 32512 21238 32524
rect 14292 32456 14964 32484
rect 6411 32388 7696 32416
rect 7745 32419 7803 32425
rect 6411 32385 6423 32388
rect 6365 32379 6423 32385
rect 7745 32385 7757 32419
rect 7791 32385 7803 32419
rect 7745 32379 7803 32385
rect 8012 32419 8070 32425
rect 8012 32385 8024 32419
rect 8058 32416 8070 32419
rect 8058 32388 9260 32416
rect 8058 32385 8070 32388
rect 8012 32379 8070 32385
rect 3418 32308 3424 32360
rect 3476 32308 3482 32360
rect 9232 32289 9260 32388
rect 9398 32376 9404 32428
rect 9456 32416 9462 32428
rect 10502 32416 10508 32428
rect 9456 32388 10508 32416
rect 9456 32376 9462 32388
rect 9490 32308 9496 32360
rect 9548 32348 9554 32360
rect 9876 32357 9904 32388
rect 10502 32376 10508 32388
rect 10560 32376 10566 32428
rect 12618 32425 12624 32428
rect 12612 32379 12624 32425
rect 12618 32376 12624 32379
rect 12676 32376 12682 32428
rect 14292 32416 14320 32456
rect 15102 32444 15108 32496
rect 15160 32484 15166 32496
rect 15381 32487 15439 32493
rect 15381 32484 15393 32487
rect 15160 32456 15393 32484
rect 15160 32444 15166 32456
rect 15381 32453 15393 32456
rect 15427 32484 15439 32487
rect 18230 32484 18236 32496
rect 15427 32456 18236 32484
rect 15427 32453 15439 32456
rect 15381 32447 15439 32453
rect 18230 32444 18236 32456
rect 18288 32444 18294 32496
rect 19242 32444 19248 32496
rect 19300 32484 19306 32496
rect 20073 32487 20131 32493
rect 20073 32484 20085 32487
rect 19300 32456 20085 32484
rect 19300 32444 19306 32456
rect 20073 32453 20085 32456
rect 20119 32453 20131 32487
rect 24688 32484 24716 32524
rect 24765 32521 24777 32555
rect 24811 32552 24823 32555
rect 25774 32552 25780 32564
rect 24811 32524 25780 32552
rect 24811 32521 24823 32524
rect 24765 32515 24823 32521
rect 25774 32512 25780 32524
rect 25832 32512 25838 32564
rect 27985 32555 28043 32561
rect 27985 32521 27997 32555
rect 28031 32552 28043 32555
rect 28258 32552 28264 32564
rect 28031 32524 28264 32552
rect 28031 32521 28043 32524
rect 27985 32515 28043 32521
rect 28258 32512 28264 32524
rect 28316 32512 28322 32564
rect 28350 32512 28356 32564
rect 28408 32552 28414 32564
rect 34146 32552 34152 32564
rect 28408 32524 34152 32552
rect 28408 32512 28414 32524
rect 34146 32512 34152 32524
rect 34204 32512 34210 32564
rect 24688 32456 27568 32484
rect 20073 32447 20131 32453
rect 13924 32388 14320 32416
rect 9677 32351 9735 32357
rect 9677 32348 9689 32351
rect 9548 32320 9689 32348
rect 9548 32308 9554 32320
rect 9677 32317 9689 32320
rect 9723 32317 9735 32351
rect 9677 32311 9735 32317
rect 9861 32351 9919 32357
rect 9861 32317 9873 32351
rect 9907 32317 9919 32351
rect 9861 32311 9919 32317
rect 10965 32351 11023 32357
rect 10965 32317 10977 32351
rect 11011 32348 11023 32351
rect 11054 32348 11060 32360
rect 11011 32320 11060 32348
rect 11011 32317 11023 32320
rect 10965 32311 11023 32317
rect 11054 32308 11060 32320
rect 11112 32348 11118 32360
rect 11514 32348 11520 32360
rect 11112 32320 11520 32348
rect 11112 32308 11118 32320
rect 11514 32308 11520 32320
rect 11572 32348 11578 32360
rect 12345 32351 12403 32357
rect 12345 32348 12357 32351
rect 11572 32320 12357 32348
rect 11572 32308 11578 32320
rect 12345 32317 12357 32320
rect 12391 32317 12403 32351
rect 12345 32311 12403 32317
rect 13354 32308 13360 32360
rect 13412 32348 13418 32360
rect 13924 32348 13952 32388
rect 17034 32376 17040 32428
rect 17092 32376 17098 32428
rect 21177 32419 21235 32425
rect 21177 32385 21189 32419
rect 21223 32385 21235 32419
rect 21177 32379 21235 32385
rect 14921 32351 14979 32357
rect 14921 32348 14933 32351
rect 13412 32320 13952 32348
rect 14292 32320 14933 32348
rect 13412 32308 13418 32320
rect 9217 32283 9275 32289
rect 9217 32249 9229 32283
rect 9263 32249 9275 32283
rect 9217 32243 9275 32249
rect 4798 32172 4804 32224
rect 4856 32172 4862 32224
rect 6549 32215 6607 32221
rect 6549 32181 6561 32215
rect 6595 32212 6607 32215
rect 6730 32212 6736 32224
rect 6595 32184 6736 32212
rect 6595 32181 6607 32184
rect 6549 32175 6607 32181
rect 6730 32172 6736 32184
rect 6788 32212 6794 32224
rect 7190 32212 7196 32224
rect 6788 32184 7196 32212
rect 6788 32172 6794 32184
rect 7190 32172 7196 32184
rect 7248 32172 7254 32224
rect 13078 32172 13084 32224
rect 13136 32212 13142 32224
rect 13630 32212 13636 32224
rect 13136 32184 13636 32212
rect 13136 32172 13142 32184
rect 13630 32172 13636 32184
rect 13688 32212 13694 32224
rect 14292 32212 14320 32320
rect 14921 32317 14933 32320
rect 14967 32317 14979 32351
rect 14921 32311 14979 32317
rect 15102 32308 15108 32360
rect 15160 32308 15166 32360
rect 16574 32348 16580 32360
rect 15396 32320 16580 32348
rect 14550 32240 14556 32292
rect 14608 32280 14614 32292
rect 15120 32280 15148 32308
rect 14608 32252 15148 32280
rect 14608 32240 14614 32252
rect 13688 32184 14320 32212
rect 13688 32172 13694 32184
rect 14458 32172 14464 32224
rect 14516 32212 14522 32224
rect 15396 32212 15424 32320
rect 16574 32308 16580 32320
rect 16632 32308 16638 32360
rect 17126 32308 17132 32360
rect 17184 32308 17190 32360
rect 17310 32308 17316 32360
rect 17368 32308 17374 32360
rect 19521 32351 19579 32357
rect 19521 32317 19533 32351
rect 19567 32348 19579 32351
rect 20165 32351 20223 32357
rect 20165 32348 20177 32351
rect 19567 32320 20177 32348
rect 19567 32317 19579 32320
rect 19521 32311 19579 32317
rect 20165 32317 20177 32320
rect 20211 32317 20223 32351
rect 21192 32348 21220 32379
rect 21266 32376 21272 32428
rect 21324 32376 21330 32428
rect 21358 32376 21364 32428
rect 21416 32416 21422 32428
rect 21453 32419 21511 32425
rect 21453 32416 21465 32419
rect 21416 32388 21465 32416
rect 21416 32376 21422 32388
rect 21453 32385 21465 32388
rect 21499 32385 21511 32419
rect 21453 32379 21511 32385
rect 21545 32419 21603 32425
rect 21545 32385 21557 32419
rect 21591 32416 21603 32419
rect 21591 32388 22140 32416
rect 21591 32385 21603 32388
rect 21545 32379 21603 32385
rect 21726 32348 21732 32360
rect 21192 32320 21732 32348
rect 20165 32311 20223 32317
rect 16114 32240 16120 32292
rect 16172 32280 16178 32292
rect 19536 32280 19564 32311
rect 21726 32308 21732 32320
rect 21784 32348 21790 32360
rect 21821 32351 21879 32357
rect 21821 32348 21833 32351
rect 21784 32320 21833 32348
rect 21784 32308 21790 32320
rect 21821 32317 21833 32320
rect 21867 32317 21879 32351
rect 21821 32311 21879 32317
rect 16172 32252 19564 32280
rect 16172 32240 16178 32252
rect 14516 32184 15424 32212
rect 14516 32172 14522 32184
rect 15562 32172 15568 32224
rect 15620 32212 15626 32224
rect 16669 32215 16727 32221
rect 16669 32212 16681 32215
rect 15620 32184 16681 32212
rect 15620 32172 15626 32184
rect 16669 32181 16681 32184
rect 16715 32181 16727 32215
rect 16669 32175 16727 32181
rect 17310 32172 17316 32224
rect 17368 32212 17374 32224
rect 17589 32215 17647 32221
rect 17589 32212 17601 32215
rect 17368 32184 17601 32212
rect 17368 32172 17374 32184
rect 17589 32181 17601 32184
rect 17635 32212 17647 32215
rect 20438 32212 20444 32224
rect 17635 32184 20444 32212
rect 17635 32181 17647 32184
rect 17589 32175 17647 32181
rect 20438 32172 20444 32184
rect 20496 32172 20502 32224
rect 22112 32221 22140 32388
rect 22554 32376 22560 32428
rect 22612 32376 22618 32428
rect 22830 32425 22836 32428
rect 22824 32379 22836 32425
rect 22830 32376 22836 32379
rect 22888 32376 22894 32428
rect 23750 32376 23756 32428
rect 23808 32416 23814 32428
rect 24857 32419 24915 32425
rect 24857 32416 24869 32419
rect 23808 32388 24869 32416
rect 23808 32376 23814 32388
rect 24857 32385 24869 32388
rect 24903 32385 24915 32419
rect 24857 32379 24915 32385
rect 25041 32351 25099 32357
rect 25041 32317 25053 32351
rect 25087 32348 25099 32351
rect 26142 32348 26148 32360
rect 25087 32320 26148 32348
rect 25087 32317 25099 32320
rect 25041 32311 25099 32317
rect 26142 32308 26148 32320
rect 26200 32308 26206 32360
rect 24397 32283 24455 32289
rect 23492 32252 24072 32280
rect 22097 32215 22155 32221
rect 22097 32181 22109 32215
rect 22143 32212 22155 32215
rect 23492 32212 23520 32252
rect 22143 32184 23520 32212
rect 22143 32181 22155 32184
rect 22097 32175 22155 32181
rect 23934 32172 23940 32224
rect 23992 32172 23998 32224
rect 24044 32212 24072 32252
rect 24397 32249 24409 32283
rect 24443 32280 24455 32283
rect 24486 32280 24492 32292
rect 24443 32252 24492 32280
rect 24443 32249 24455 32252
rect 24397 32243 24455 32249
rect 24486 32240 24492 32252
rect 24544 32240 24550 32292
rect 27540 32280 27568 32456
rect 27798 32444 27804 32496
rect 27856 32484 27862 32496
rect 28626 32484 28632 32496
rect 27856 32456 28632 32484
rect 27856 32444 27862 32456
rect 28626 32444 28632 32456
rect 28684 32484 28690 32496
rect 28813 32487 28871 32493
rect 28813 32484 28825 32487
rect 28684 32456 28825 32484
rect 28684 32444 28690 32456
rect 28813 32453 28825 32456
rect 28859 32453 28871 32487
rect 28813 32447 28871 32453
rect 29638 32444 29644 32496
rect 29696 32484 29702 32496
rect 29825 32487 29883 32493
rect 29825 32484 29837 32487
rect 29696 32456 29837 32484
rect 29696 32444 29702 32456
rect 29825 32453 29837 32456
rect 29871 32453 29883 32487
rect 29825 32447 29883 32453
rect 27614 32376 27620 32428
rect 27672 32416 27678 32428
rect 28166 32416 28172 32428
rect 27672 32388 28172 32416
rect 27672 32376 27678 32388
rect 28166 32376 28172 32388
rect 28224 32376 28230 32428
rect 28258 32376 28264 32428
rect 28316 32376 28322 32428
rect 28353 32419 28411 32425
rect 28353 32385 28365 32419
rect 28399 32385 28411 32419
rect 28353 32379 28411 32385
rect 28368 32348 28396 32379
rect 28534 32376 28540 32428
rect 28592 32376 28598 32428
rect 28442 32348 28448 32360
rect 28368 32320 28448 32348
rect 28442 32308 28448 32320
rect 28500 32348 28506 32360
rect 28629 32351 28687 32357
rect 28629 32348 28641 32351
rect 28500 32320 28641 32348
rect 28500 32308 28506 32320
rect 28629 32317 28641 32320
rect 28675 32317 28687 32351
rect 28629 32311 28687 32317
rect 29546 32280 29552 32292
rect 27540 32252 29552 32280
rect 29546 32240 29552 32252
rect 29604 32280 29610 32292
rect 30282 32280 30288 32292
rect 29604 32252 30288 32280
rect 29604 32240 29610 32252
rect 30282 32240 30288 32252
rect 30340 32240 30346 32292
rect 26694 32212 26700 32224
rect 24044 32184 26700 32212
rect 26694 32172 26700 32184
rect 26752 32172 26758 32224
rect 1104 32122 35328 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 35328 32122
rect 1104 32048 35328 32070
rect 6641 32011 6699 32017
rect 6641 31977 6653 32011
rect 6687 32008 6699 32011
rect 7098 32008 7104 32020
rect 6687 31980 7104 32008
rect 6687 31977 6699 31980
rect 6641 31971 6699 31977
rect 7098 31968 7104 31980
rect 7156 31968 7162 32020
rect 7374 31968 7380 32020
rect 7432 32008 7438 32020
rect 7561 32011 7619 32017
rect 7561 32008 7573 32011
rect 7432 31980 7573 32008
rect 7432 31968 7438 31980
rect 7561 31977 7573 31980
rect 7607 31977 7619 32011
rect 7561 31971 7619 31977
rect 8846 31968 8852 32020
rect 8904 32008 8910 32020
rect 9306 32008 9312 32020
rect 8904 31980 9312 32008
rect 8904 31968 8910 31980
rect 9306 31968 9312 31980
rect 9364 31968 9370 32020
rect 9582 31968 9588 32020
rect 9640 31968 9646 32020
rect 9769 32011 9827 32017
rect 9769 31977 9781 32011
rect 9815 32008 9827 32011
rect 9858 32008 9864 32020
rect 9815 31980 9864 32008
rect 9815 31977 9827 31980
rect 9769 31971 9827 31977
rect 9858 31968 9864 31980
rect 9916 31968 9922 32020
rect 11054 32008 11060 32020
rect 10152 31980 11060 32008
rect 6733 31943 6791 31949
rect 6733 31909 6745 31943
rect 6779 31909 6791 31943
rect 9490 31940 9496 31952
rect 6733 31903 6791 31909
rect 7576 31912 9496 31940
rect 4341 31875 4399 31881
rect 4341 31841 4353 31875
rect 4387 31872 4399 31875
rect 4706 31872 4712 31884
rect 4387 31844 4712 31872
rect 4387 31841 4399 31844
rect 4341 31835 4399 31841
rect 4706 31832 4712 31844
rect 4764 31832 4770 31884
rect 1394 31764 1400 31816
rect 1452 31764 1458 31816
rect 1673 31807 1731 31813
rect 1673 31773 1685 31807
rect 1719 31804 1731 31807
rect 1719 31776 2452 31804
rect 1719 31773 1731 31776
rect 1673 31767 1731 31773
rect 2424 31677 2452 31776
rect 4614 31764 4620 31816
rect 4672 31764 4678 31816
rect 5258 31764 5264 31816
rect 5316 31764 5322 31816
rect 5528 31807 5586 31813
rect 5528 31773 5540 31807
rect 5574 31804 5586 31807
rect 6748 31804 6776 31903
rect 7282 31832 7288 31884
rect 7340 31832 7346 31884
rect 7576 31872 7604 31912
rect 9490 31900 9496 31912
rect 9548 31900 9554 31952
rect 7392 31844 7604 31872
rect 5574 31776 6776 31804
rect 5574 31773 5586 31776
rect 5528 31767 5586 31773
rect 7190 31764 7196 31816
rect 7248 31804 7254 31816
rect 7392 31804 7420 31844
rect 8202 31832 8208 31884
rect 8260 31872 8266 31884
rect 10152 31881 10180 31980
rect 11054 31968 11060 31980
rect 11112 31968 11118 32020
rect 12618 31968 12624 32020
rect 12676 32008 12682 32020
rect 12805 32011 12863 32017
rect 12805 32008 12817 32011
rect 12676 31980 12817 32008
rect 12676 31968 12682 31980
rect 12805 31977 12817 31980
rect 12851 31977 12863 32011
rect 12805 31971 12863 31977
rect 16669 32011 16727 32017
rect 16669 31977 16681 32011
rect 16715 32008 16727 32011
rect 17126 32008 17132 32020
rect 16715 31980 17132 32008
rect 16715 31977 16727 31980
rect 16669 31971 16727 31977
rect 17126 31968 17132 31980
rect 17184 31968 17190 32020
rect 21450 31968 21456 32020
rect 21508 31968 21514 32020
rect 22094 31968 22100 32020
rect 22152 32008 22158 32020
rect 22152 31980 22416 32008
rect 22152 31968 22158 31980
rect 11609 31943 11667 31949
rect 11609 31909 11621 31943
rect 11655 31909 11667 31943
rect 11609 31903 11667 31909
rect 10137 31875 10195 31881
rect 10137 31872 10149 31875
rect 8260 31844 10149 31872
rect 8260 31832 8266 31844
rect 10137 31841 10149 31844
rect 10183 31841 10195 31875
rect 10137 31835 10195 31841
rect 7248 31776 7420 31804
rect 7248 31764 7254 31776
rect 7466 31764 7472 31816
rect 7524 31804 7530 31816
rect 7745 31807 7803 31813
rect 7745 31804 7757 31807
rect 7524 31776 7757 31804
rect 7524 31764 7530 31776
rect 7745 31773 7757 31776
rect 7791 31773 7803 31807
rect 7745 31767 7803 31773
rect 8110 31764 8116 31816
rect 8168 31764 8174 31816
rect 8754 31764 8760 31816
rect 8812 31804 8818 31816
rect 9122 31813 9128 31816
rect 8941 31807 8999 31813
rect 8941 31804 8953 31807
rect 8812 31776 8953 31804
rect 8812 31764 8818 31776
rect 8941 31773 8953 31776
rect 8987 31773 8999 31807
rect 8941 31767 8999 31773
rect 9089 31807 9128 31813
rect 9089 31773 9101 31807
rect 9089 31767 9128 31773
rect 9122 31764 9128 31767
rect 9180 31764 9186 31816
rect 9306 31764 9312 31816
rect 9364 31764 9370 31816
rect 9398 31764 9404 31816
rect 9456 31813 9462 31816
rect 9456 31767 9464 31813
rect 9858 31804 9864 31816
rect 9508 31776 9864 31804
rect 9456 31764 9462 31767
rect 7098 31696 7104 31748
rect 7156 31736 7162 31748
rect 7837 31739 7895 31745
rect 7837 31736 7849 31739
rect 7156 31708 7849 31736
rect 7156 31696 7162 31708
rect 7837 31705 7849 31708
rect 7883 31705 7895 31739
rect 7837 31699 7895 31705
rect 7929 31739 7987 31745
rect 7929 31705 7941 31739
rect 7975 31705 7987 31739
rect 7929 31699 7987 31705
rect 9217 31739 9275 31745
rect 9217 31705 9229 31739
rect 9263 31736 9275 31739
rect 9508 31736 9536 31776
rect 9858 31764 9864 31776
rect 9916 31764 9922 31816
rect 10404 31807 10462 31813
rect 10404 31773 10416 31807
rect 10450 31804 10462 31807
rect 11624 31804 11652 31903
rect 18230 31900 18236 31952
rect 18288 31940 18294 31952
rect 22388 31949 22416 31980
rect 22830 31968 22836 32020
rect 22888 32008 22894 32020
rect 23109 32011 23167 32017
rect 23109 32008 23121 32011
rect 22888 31980 23121 32008
rect 22888 31968 22894 31980
rect 23109 31977 23121 31980
rect 23155 31977 23167 32011
rect 23109 31971 23167 31977
rect 26050 31968 26056 32020
rect 26108 31968 26114 32020
rect 26237 32011 26295 32017
rect 26237 31977 26249 32011
rect 26283 32008 26295 32011
rect 27982 32008 27988 32020
rect 26283 31980 27988 32008
rect 26283 31977 26295 31980
rect 26237 31971 26295 31977
rect 27982 31968 27988 31980
rect 28040 31968 28046 32020
rect 28077 32011 28135 32017
rect 28077 31977 28089 32011
rect 28123 32008 28135 32011
rect 28534 32008 28540 32020
rect 28123 31980 28540 32008
rect 28123 31977 28135 31980
rect 28077 31971 28135 31977
rect 28534 31968 28540 31980
rect 28592 31968 28598 32020
rect 29549 32011 29607 32017
rect 29549 31977 29561 32011
rect 29595 32008 29607 32011
rect 29822 32008 29828 32020
rect 29595 31980 29828 32008
rect 29595 31977 29607 31980
rect 29549 31971 29607 31977
rect 29822 31968 29828 31980
rect 29880 31968 29886 32020
rect 22373 31943 22431 31949
rect 18288 31912 22324 31940
rect 18288 31900 18294 31912
rect 12253 31875 12311 31881
rect 12253 31841 12265 31875
rect 12299 31872 12311 31875
rect 12529 31875 12587 31881
rect 12529 31872 12541 31875
rect 12299 31844 12541 31872
rect 12299 31841 12311 31844
rect 12253 31835 12311 31841
rect 12529 31841 12541 31844
rect 12575 31872 12587 31875
rect 12710 31872 12716 31884
rect 12575 31844 12716 31872
rect 12575 31841 12587 31844
rect 12529 31835 12587 31841
rect 12710 31832 12716 31844
rect 12768 31832 12774 31884
rect 13449 31875 13507 31881
rect 13449 31841 13461 31875
rect 13495 31841 13507 31875
rect 13449 31835 13507 31841
rect 10450 31776 11652 31804
rect 11977 31807 12035 31813
rect 10450 31773 10462 31776
rect 10404 31767 10462 31773
rect 11977 31773 11989 31807
rect 12023 31804 12035 31807
rect 12066 31804 12072 31816
rect 12023 31776 12072 31804
rect 12023 31773 12035 31776
rect 11977 31767 12035 31773
rect 12066 31764 12072 31776
rect 12124 31764 12130 31816
rect 12986 31764 12992 31816
rect 13044 31804 13050 31816
rect 13173 31807 13231 31813
rect 13173 31804 13185 31807
rect 13044 31776 13185 31804
rect 13044 31764 13050 31776
rect 13173 31773 13185 31776
rect 13219 31773 13231 31807
rect 13173 31767 13231 31773
rect 9263 31708 9536 31736
rect 9263 31705 9275 31708
rect 9217 31699 9275 31705
rect 2409 31671 2467 31677
rect 2409 31637 2421 31671
rect 2455 31668 2467 31671
rect 7558 31668 7564 31680
rect 2455 31640 7564 31668
rect 2455 31637 2467 31640
rect 2409 31631 2467 31637
rect 7558 31628 7564 31640
rect 7616 31628 7622 31680
rect 7944 31668 7972 31699
rect 11882 31696 11888 31748
rect 11940 31736 11946 31748
rect 13265 31739 13323 31745
rect 13265 31736 13277 31739
rect 11940 31708 13277 31736
rect 11940 31696 11946 31708
rect 13265 31705 13277 31708
rect 13311 31705 13323 31739
rect 13464 31736 13492 31835
rect 20898 31832 20904 31884
rect 20956 31872 20962 31884
rect 21174 31872 21180 31884
rect 20956 31844 21180 31872
rect 20956 31832 20962 31844
rect 21174 31832 21180 31844
rect 21232 31872 21238 31884
rect 21913 31875 21971 31881
rect 21913 31872 21925 31875
rect 21232 31844 21925 31872
rect 21232 31832 21238 31844
rect 21913 31841 21925 31844
rect 21959 31841 21971 31875
rect 21913 31835 21971 31841
rect 22094 31832 22100 31884
rect 22152 31832 22158 31884
rect 15289 31807 15347 31813
rect 15289 31773 15301 31807
rect 15335 31804 15347 31807
rect 16666 31804 16672 31816
rect 15335 31776 16672 31804
rect 15335 31773 15347 31776
rect 15289 31767 15347 31773
rect 16666 31764 16672 31776
rect 16724 31804 16730 31816
rect 17221 31807 17279 31813
rect 17221 31804 17233 31807
rect 16724 31776 17233 31804
rect 16724 31764 16730 31776
rect 17221 31773 17233 31776
rect 17267 31773 17279 31807
rect 17221 31767 17279 31773
rect 21266 31764 21272 31816
rect 21324 31804 21330 31816
rect 21821 31807 21879 31813
rect 21821 31804 21833 31807
rect 21324 31776 21833 31804
rect 21324 31764 21330 31776
rect 21821 31773 21833 31776
rect 21867 31773 21879 31807
rect 22296 31804 22324 31912
rect 22373 31909 22385 31943
rect 22419 31940 22431 31943
rect 22922 31940 22928 31952
rect 22419 31912 22928 31940
rect 22419 31909 22431 31912
rect 22373 31903 22431 31909
rect 22922 31900 22928 31912
rect 22980 31900 22986 31952
rect 27890 31900 27896 31952
rect 27948 31940 27954 31952
rect 28169 31943 28227 31949
rect 28169 31940 28181 31943
rect 27948 31912 28181 31940
rect 27948 31900 27954 31912
rect 28169 31909 28181 31912
rect 28215 31909 28227 31943
rect 28169 31903 28227 31909
rect 23661 31875 23719 31881
rect 23661 31872 23673 31875
rect 22940 31844 23673 31872
rect 22940 31813 22968 31844
rect 23661 31841 23673 31844
rect 23707 31841 23719 31875
rect 23661 31835 23719 31841
rect 28813 31875 28871 31881
rect 28813 31841 28825 31875
rect 28859 31841 28871 31875
rect 28813 31835 28871 31841
rect 22925 31807 22983 31813
rect 22925 31804 22937 31807
rect 22296 31776 22937 31804
rect 21821 31767 21879 31773
rect 22925 31773 22937 31776
rect 22971 31773 22983 31807
rect 22925 31767 22983 31773
rect 23569 31807 23627 31813
rect 23569 31773 23581 31807
rect 23615 31804 23627 31807
rect 23750 31804 23756 31816
rect 23615 31776 23756 31804
rect 23615 31773 23627 31776
rect 23569 31767 23627 31773
rect 23750 31764 23756 31776
rect 23808 31764 23814 31816
rect 25866 31764 25872 31816
rect 25924 31764 25930 31816
rect 25958 31764 25964 31816
rect 26016 31764 26022 31816
rect 26697 31807 26755 31813
rect 26697 31773 26709 31807
rect 26743 31804 26755 31807
rect 26786 31804 26792 31816
rect 26743 31776 26792 31804
rect 26743 31773 26755 31776
rect 26697 31767 26755 31773
rect 26786 31764 26792 31776
rect 26844 31804 26850 31816
rect 26844 31776 27200 31804
rect 26844 31764 26850 31776
rect 27172 31754 27200 31776
rect 28534 31764 28540 31816
rect 28592 31764 28598 31816
rect 28828 31804 28856 31835
rect 29914 31832 29920 31884
rect 29972 31872 29978 31884
rect 30009 31875 30067 31881
rect 30009 31872 30021 31875
rect 29972 31844 30021 31872
rect 29972 31832 29978 31844
rect 30009 31841 30021 31844
rect 30055 31841 30067 31875
rect 30009 31835 30067 31841
rect 30098 31832 30104 31884
rect 30156 31872 30162 31884
rect 30193 31875 30251 31881
rect 30193 31872 30205 31875
rect 30156 31844 30205 31872
rect 30156 31832 30162 31844
rect 30193 31841 30205 31844
rect 30239 31872 30251 31875
rect 30929 31875 30987 31881
rect 30929 31872 30941 31875
rect 30239 31844 30941 31872
rect 30239 31841 30251 31844
rect 30193 31835 30251 31841
rect 30929 31841 30941 31844
rect 30975 31841 30987 31875
rect 30929 31835 30987 31841
rect 32766 31832 32772 31884
rect 32824 31832 32830 31884
rect 33045 31875 33103 31881
rect 33045 31841 33057 31875
rect 33091 31872 33103 31875
rect 33778 31872 33784 31884
rect 33091 31844 33784 31872
rect 33091 31841 33103 31844
rect 33045 31835 33103 31841
rect 33778 31832 33784 31844
rect 33836 31832 33842 31884
rect 29089 31807 29147 31813
rect 29089 31804 29101 31807
rect 28828 31776 29101 31804
rect 29089 31773 29101 31776
rect 29135 31804 29147 31807
rect 29454 31804 29460 31816
rect 29135 31776 29460 31804
rect 29135 31773 29147 31776
rect 29089 31767 29147 31773
rect 29454 31764 29460 31776
rect 29512 31764 29518 31816
rect 15562 31745 15568 31748
rect 13464 31708 13768 31736
rect 13265 31699 13323 31705
rect 8297 31671 8355 31677
rect 8297 31668 8309 31671
rect 7944 31640 8309 31668
rect 8297 31637 8309 31640
rect 8343 31668 8355 31671
rect 10686 31668 10692 31680
rect 8343 31640 10692 31668
rect 8343 31637 8355 31640
rect 8297 31631 8355 31637
rect 10686 31628 10692 31640
rect 10744 31628 10750 31680
rect 11517 31671 11575 31677
rect 11517 31637 11529 31671
rect 11563 31668 11575 31671
rect 12066 31668 12072 31680
rect 11563 31640 12072 31668
rect 11563 31637 11575 31640
rect 11517 31631 11575 31637
rect 12066 31628 12072 31640
rect 12124 31628 12130 31680
rect 13740 31677 13768 31708
rect 15556 31699 15568 31745
rect 15562 31696 15568 31699
rect 15620 31696 15626 31748
rect 17488 31739 17546 31745
rect 17488 31705 17500 31739
rect 17534 31736 17546 31739
rect 17770 31736 17776 31748
rect 17534 31708 17776 31736
rect 17534 31705 17546 31708
rect 17488 31699 17546 31705
rect 17770 31696 17776 31708
rect 17828 31696 17834 31748
rect 23014 31736 23020 31748
rect 17880 31708 23020 31736
rect 13725 31671 13783 31677
rect 13725 31637 13737 31671
rect 13771 31668 13783 31671
rect 16114 31668 16120 31680
rect 13771 31640 16120 31668
rect 13771 31637 13783 31640
rect 13725 31631 13783 31637
rect 16114 31628 16120 31640
rect 16172 31628 16178 31680
rect 17402 31628 17408 31680
rect 17460 31668 17466 31680
rect 17880 31668 17908 31708
rect 23014 31696 23020 31708
rect 23072 31696 23078 31748
rect 23106 31696 23112 31748
rect 23164 31736 23170 31748
rect 26964 31739 27022 31745
rect 23164 31708 23612 31736
rect 23164 31696 23170 31708
rect 17460 31640 17908 31668
rect 17460 31628 17466 31640
rect 18138 31628 18144 31680
rect 18196 31668 18202 31680
rect 18601 31671 18659 31677
rect 18601 31668 18613 31671
rect 18196 31640 18613 31668
rect 18196 31628 18202 31640
rect 18601 31637 18613 31640
rect 18647 31637 18659 31671
rect 18601 31631 18659 31637
rect 22738 31628 22744 31680
rect 22796 31668 22802 31680
rect 23290 31668 23296 31680
rect 22796 31640 23296 31668
rect 22796 31628 22802 31640
rect 23290 31628 23296 31640
rect 23348 31628 23354 31680
rect 23474 31628 23480 31680
rect 23532 31628 23538 31680
rect 23584 31668 23612 31708
rect 26964 31705 26976 31739
rect 27010 31736 27022 31739
rect 27062 31736 27068 31748
rect 27010 31708 27068 31736
rect 27010 31705 27022 31708
rect 26964 31699 27022 31705
rect 27062 31696 27068 31708
rect 27120 31696 27126 31748
rect 27172 31736 27375 31754
rect 27430 31736 27436 31748
rect 27172 31726 27436 31736
rect 27347 31708 27436 31726
rect 27430 31696 27436 31708
rect 27488 31696 27494 31748
rect 27522 31696 27528 31748
rect 27580 31736 27586 31748
rect 27580 31708 27936 31736
rect 27580 31696 27586 31708
rect 27798 31668 27804 31680
rect 23584 31640 27804 31668
rect 27798 31628 27804 31640
rect 27856 31628 27862 31680
rect 27908 31668 27936 31708
rect 28166 31696 28172 31748
rect 28224 31736 28230 31748
rect 28629 31739 28687 31745
rect 28629 31736 28641 31739
rect 28224 31708 28641 31736
rect 28224 31696 28230 31708
rect 28629 31705 28641 31708
rect 28675 31736 28687 31739
rect 28902 31736 28908 31748
rect 28675 31708 28908 31736
rect 28675 31705 28687 31708
rect 28629 31699 28687 31705
rect 28902 31696 28908 31708
rect 28960 31736 28966 31748
rect 29917 31739 29975 31745
rect 29917 31736 29929 31739
rect 28960 31708 29929 31736
rect 28960 31696 28966 31708
rect 29917 31705 29929 31708
rect 29963 31705 29975 31739
rect 30745 31739 30803 31745
rect 30745 31736 30757 31739
rect 29917 31699 29975 31705
rect 30024 31708 30757 31736
rect 30024 31668 30052 31708
rect 30745 31705 30757 31708
rect 30791 31705 30803 31739
rect 30745 31699 30803 31705
rect 33502 31696 33508 31748
rect 33560 31696 33566 31748
rect 27908 31640 30052 31668
rect 30374 31628 30380 31680
rect 30432 31628 30438 31680
rect 30834 31628 30840 31680
rect 30892 31628 30898 31680
rect 34514 31628 34520 31680
rect 34572 31628 34578 31680
rect 1104 31578 35328 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35328 31578
rect 1104 31504 35328 31526
rect 1394 31424 1400 31476
rect 1452 31424 1458 31476
rect 2593 31467 2651 31473
rect 2593 31433 2605 31467
rect 2639 31464 2651 31467
rect 5166 31464 5172 31476
rect 2639 31436 5172 31464
rect 2639 31433 2651 31436
rect 2593 31427 2651 31433
rect 5166 31424 5172 31436
rect 5224 31464 5230 31476
rect 5353 31467 5411 31473
rect 5353 31464 5365 31467
rect 5224 31436 5365 31464
rect 5224 31424 5230 31436
rect 5353 31433 5365 31436
rect 5399 31433 5411 31467
rect 5353 31427 5411 31433
rect 6365 31467 6423 31473
rect 6365 31433 6377 31467
rect 6411 31464 6423 31467
rect 6914 31464 6920 31476
rect 6411 31436 6920 31464
rect 6411 31433 6423 31436
rect 6365 31427 6423 31433
rect 6914 31424 6920 31436
rect 6972 31464 6978 31476
rect 8110 31464 8116 31476
rect 6972 31436 8116 31464
rect 6972 31424 6978 31436
rect 8110 31424 8116 31436
rect 8168 31424 8174 31476
rect 9306 31424 9312 31476
rect 9364 31464 9370 31476
rect 9493 31467 9551 31473
rect 9493 31464 9505 31467
rect 9364 31436 9505 31464
rect 9364 31424 9370 31436
rect 9493 31433 9505 31436
rect 9539 31433 9551 31467
rect 9493 31427 9551 31433
rect 9585 31467 9643 31473
rect 9585 31433 9597 31467
rect 9631 31433 9643 31467
rect 9585 31427 9643 31433
rect 3418 31356 3424 31408
rect 3476 31396 3482 31408
rect 7282 31396 7288 31408
rect 3476 31368 4016 31396
rect 3476 31356 3482 31368
rect 3988 31337 4016 31368
rect 6196 31368 7288 31396
rect 3717 31331 3775 31337
rect 3717 31297 3729 31331
rect 3763 31328 3775 31331
rect 3973 31331 4031 31337
rect 3763 31300 3924 31328
rect 3763 31297 3775 31300
rect 3717 31291 3775 31297
rect 3896 31260 3924 31300
rect 3973 31297 3985 31331
rect 4019 31297 4031 31331
rect 3973 31291 4031 31297
rect 4062 31288 4068 31340
rect 4120 31288 4126 31340
rect 4341 31331 4399 31337
rect 4341 31297 4353 31331
rect 4387 31328 4399 31331
rect 4614 31328 4620 31340
rect 4387 31300 4620 31328
rect 4387 31297 4399 31300
rect 4341 31291 4399 31297
rect 4614 31288 4620 31300
rect 4672 31288 4678 31340
rect 3896 31232 4016 31260
rect 3988 31192 4016 31232
rect 4706 31220 4712 31272
rect 4764 31260 4770 31272
rect 5350 31260 5356 31272
rect 4764 31232 5356 31260
rect 4764 31220 4770 31232
rect 5350 31220 5356 31232
rect 5408 31260 5414 31272
rect 5445 31263 5503 31269
rect 5445 31260 5457 31263
rect 5408 31232 5457 31260
rect 5408 31220 5414 31232
rect 5445 31229 5457 31232
rect 5491 31229 5503 31263
rect 5445 31223 5503 31229
rect 5629 31263 5687 31269
rect 5629 31229 5641 31263
rect 5675 31260 5687 31263
rect 6196 31260 6224 31368
rect 7282 31356 7288 31368
rect 7340 31356 7346 31408
rect 8380 31399 8438 31405
rect 8380 31365 8392 31399
rect 8426 31396 8438 31399
rect 9600 31396 9628 31427
rect 9674 31424 9680 31476
rect 9732 31464 9738 31476
rect 10045 31467 10103 31473
rect 10045 31464 10057 31467
rect 9732 31436 10057 31464
rect 9732 31424 9738 31436
rect 10045 31433 10057 31436
rect 10091 31433 10103 31467
rect 12342 31464 12348 31476
rect 10045 31427 10103 31433
rect 11716 31436 12348 31464
rect 8426 31368 9628 31396
rect 8426 31365 8438 31368
rect 8380 31359 8438 31365
rect 6270 31288 6276 31340
rect 6328 31328 6334 31340
rect 7478 31331 7536 31337
rect 7478 31328 7490 31331
rect 6328 31300 7490 31328
rect 6328 31288 6334 31300
rect 7478 31297 7490 31300
rect 7524 31297 7536 31331
rect 7478 31291 7536 31297
rect 7745 31331 7803 31337
rect 7745 31297 7757 31331
rect 7791 31328 7803 31331
rect 8113 31331 8171 31337
rect 8113 31328 8125 31331
rect 7791 31300 8125 31328
rect 7791 31297 7803 31300
rect 7745 31291 7803 31297
rect 8113 31297 8125 31300
rect 8159 31328 8171 31331
rect 8202 31328 8208 31340
rect 8159 31300 8208 31328
rect 8159 31297 8171 31300
rect 8113 31291 8171 31297
rect 8202 31288 8208 31300
rect 8260 31288 8266 31340
rect 9306 31288 9312 31340
rect 9364 31328 9370 31340
rect 9953 31331 10011 31337
rect 9953 31328 9965 31331
rect 9364 31300 9965 31328
rect 9364 31288 9370 31300
rect 9953 31297 9965 31300
rect 9999 31297 10011 31331
rect 9953 31291 10011 31297
rect 10870 31288 10876 31340
rect 10928 31288 10934 31340
rect 11054 31288 11060 31340
rect 11112 31288 11118 31340
rect 11149 31331 11207 31337
rect 11149 31297 11161 31331
rect 11195 31328 11207 31331
rect 11238 31328 11244 31340
rect 11195 31300 11244 31328
rect 11195 31297 11207 31300
rect 11149 31291 11207 31297
rect 11238 31288 11244 31300
rect 11296 31288 11302 31340
rect 11716 31337 11744 31436
rect 12342 31424 12348 31436
rect 12400 31464 12406 31476
rect 15654 31464 15660 31476
rect 12400 31436 15660 31464
rect 12400 31424 12406 31436
rect 15654 31424 15660 31436
rect 15712 31464 15718 31476
rect 16482 31464 16488 31476
rect 15712 31436 16488 31464
rect 15712 31424 15718 31436
rect 16482 31424 16488 31436
rect 16540 31424 16546 31476
rect 17402 31424 17408 31476
rect 17460 31424 17466 31476
rect 17770 31424 17776 31476
rect 17828 31424 17834 31476
rect 21082 31424 21088 31476
rect 21140 31424 21146 31476
rect 21453 31467 21511 31473
rect 21453 31433 21465 31467
rect 21499 31464 21511 31467
rect 25590 31464 25596 31476
rect 21499 31436 25596 31464
rect 21499 31433 21511 31436
rect 21453 31427 21511 31433
rect 11790 31356 11796 31408
rect 11848 31356 11854 31408
rect 11885 31399 11943 31405
rect 11885 31365 11897 31399
rect 11931 31396 11943 31399
rect 12710 31396 12716 31408
rect 11931 31368 12716 31396
rect 11931 31365 11943 31368
rect 11885 31359 11943 31365
rect 12710 31356 12716 31368
rect 12768 31356 12774 31408
rect 16758 31396 16764 31408
rect 16684 31368 16764 31396
rect 11696 31331 11754 31337
rect 11696 31297 11708 31331
rect 11742 31297 11754 31331
rect 12066 31328 12072 31340
rect 12027 31300 12072 31328
rect 11696 31291 11754 31297
rect 12066 31288 12072 31300
rect 12124 31288 12130 31340
rect 12161 31331 12219 31337
rect 12161 31297 12173 31331
rect 12207 31328 12219 31331
rect 12526 31328 12532 31340
rect 12207 31300 12532 31328
rect 12207 31297 12219 31300
rect 12161 31291 12219 31297
rect 12526 31288 12532 31300
rect 12584 31328 12590 31340
rect 13538 31328 13544 31340
rect 12584 31300 13544 31328
rect 12584 31288 12590 31300
rect 13538 31288 13544 31300
rect 13596 31288 13602 31340
rect 16684 31337 16712 31368
rect 16758 31356 16764 31368
rect 16816 31396 16822 31408
rect 17586 31396 17592 31408
rect 16816 31368 17592 31396
rect 16816 31356 16822 31368
rect 17586 31356 17592 31368
rect 17644 31356 17650 31408
rect 18233 31399 18291 31405
rect 18233 31365 18245 31399
rect 18279 31396 18291 31399
rect 19702 31396 19708 31408
rect 18279 31368 19708 31396
rect 18279 31365 18291 31368
rect 18233 31359 18291 31365
rect 19702 31356 19708 31368
rect 19760 31356 19766 31408
rect 20809 31399 20867 31405
rect 20809 31365 20821 31399
rect 20855 31396 20867 31399
rect 21266 31396 21272 31408
rect 20855 31368 21272 31396
rect 20855 31365 20867 31368
rect 20809 31359 20867 31365
rect 21266 31356 21272 31368
rect 21324 31356 21330 31408
rect 16669 31331 16727 31337
rect 16669 31297 16681 31331
rect 16715 31297 16727 31331
rect 16669 31291 16727 31297
rect 16850 31288 16856 31340
rect 16908 31288 16914 31340
rect 17126 31288 17132 31340
rect 17184 31328 17190 31340
rect 17221 31331 17279 31337
rect 17221 31328 17233 31331
rect 17184 31300 17233 31328
rect 17184 31288 17190 31300
rect 17221 31297 17233 31300
rect 17267 31297 17279 31331
rect 17221 31291 17279 31297
rect 17310 31288 17316 31340
rect 17368 31328 17374 31340
rect 17368 31300 17816 31328
rect 17368 31288 17374 31300
rect 5675 31232 6224 31260
rect 10137 31263 10195 31269
rect 5675 31229 5687 31232
rect 5629 31223 5687 31229
rect 10137 31229 10149 31263
rect 10183 31229 10195 31263
rect 16945 31263 17003 31269
rect 16945 31260 16957 31263
rect 10137 31223 10195 31229
rect 11900 31232 16957 31260
rect 4985 31195 5043 31201
rect 4985 31192 4997 31195
rect 3988 31164 4997 31192
rect 4985 31161 4997 31164
rect 5031 31161 5043 31195
rect 4985 31155 5043 31161
rect 9674 31152 9680 31204
rect 9732 31192 9738 31204
rect 10152 31192 10180 31223
rect 11517 31195 11575 31201
rect 11517 31192 11529 31195
rect 9732 31164 10180 31192
rect 11164 31164 11529 31192
rect 9732 31152 9738 31164
rect 4614 31084 4620 31136
rect 4672 31124 4678 31136
rect 10410 31124 10416 31136
rect 4672 31096 10416 31124
rect 4672 31084 4678 31096
rect 10410 31084 10416 31096
rect 10468 31084 10474 31136
rect 11164 31133 11192 31164
rect 11517 31161 11529 31164
rect 11563 31161 11575 31195
rect 11517 31155 11575 31161
rect 11149 31127 11207 31133
rect 11149 31093 11161 31127
rect 11195 31093 11207 31127
rect 11149 31087 11207 31093
rect 11333 31127 11391 31133
rect 11333 31093 11345 31127
rect 11379 31124 11391 31127
rect 11900 31124 11928 31232
rect 16945 31229 16957 31232
rect 16991 31229 17003 31263
rect 16945 31223 17003 31229
rect 17037 31263 17095 31269
rect 17037 31229 17049 31263
rect 17083 31260 17095 31263
rect 17678 31260 17684 31272
rect 17083 31232 17684 31260
rect 17083 31229 17095 31232
rect 17037 31223 17095 31229
rect 17678 31220 17684 31232
rect 17736 31220 17742 31272
rect 17788 31260 17816 31300
rect 18138 31288 18144 31340
rect 18196 31288 18202 31340
rect 18598 31288 18604 31340
rect 18656 31288 18662 31340
rect 18868 31331 18926 31337
rect 18868 31297 18880 31331
rect 18914 31328 18926 31331
rect 19242 31328 19248 31340
rect 18914 31300 19248 31328
rect 18914 31297 18926 31300
rect 18868 31291 18926 31297
rect 19242 31288 19248 31300
rect 19300 31288 19306 31340
rect 20533 31331 20591 31337
rect 20533 31328 20545 31331
rect 19996 31300 20545 31328
rect 18322 31260 18328 31272
rect 17788 31232 18328 31260
rect 18322 31220 18328 31232
rect 18380 31220 18386 31272
rect 11379 31096 11928 31124
rect 11379 31093 11391 31096
rect 11333 31087 11391 31093
rect 12342 31084 12348 31136
rect 12400 31084 12406 31136
rect 12526 31084 12532 31136
rect 12584 31084 12590 31136
rect 12710 31084 12716 31136
rect 12768 31084 12774 31136
rect 17696 31133 17724 31220
rect 19996 31136 20024 31300
rect 20533 31297 20545 31300
rect 20579 31297 20591 31331
rect 20533 31291 20591 31297
rect 20717 31331 20775 31337
rect 20717 31297 20729 31331
rect 20763 31297 20775 31331
rect 20717 31291 20775 31297
rect 20901 31331 20959 31337
rect 20901 31297 20913 31331
rect 20947 31328 20959 31331
rect 21468 31328 21496 31427
rect 25590 31424 25596 31436
rect 25648 31424 25654 31476
rect 25866 31424 25872 31476
rect 25924 31464 25930 31476
rect 26053 31467 26111 31473
rect 26053 31464 26065 31467
rect 25924 31436 26065 31464
rect 25924 31424 25930 31436
rect 26053 31433 26065 31436
rect 26099 31433 26111 31467
rect 26789 31467 26847 31473
rect 26789 31464 26801 31467
rect 26053 31427 26111 31433
rect 26160 31436 26801 31464
rect 24670 31396 24676 31408
rect 23124 31368 24676 31396
rect 23124 31328 23152 31368
rect 24670 31356 24676 31368
rect 24728 31356 24734 31408
rect 20947 31300 21496 31328
rect 22848 31300 23152 31328
rect 23201 31331 23259 31337
rect 20947 31297 20959 31300
rect 20901 31291 20959 31297
rect 20732 31260 20760 31291
rect 21269 31263 21327 31269
rect 21269 31260 21281 31263
rect 20732 31232 21281 31260
rect 21269 31229 21281 31232
rect 21315 31260 21327 31263
rect 22848 31260 22876 31300
rect 23201 31297 23213 31331
rect 23247 31328 23259 31331
rect 24848 31331 24906 31337
rect 23247 31300 23612 31328
rect 23247 31297 23259 31300
rect 23201 31291 23259 31297
rect 23584 31272 23612 31300
rect 24848 31297 24860 31331
rect 24894 31328 24906 31331
rect 25130 31328 25136 31340
rect 24894 31300 25136 31328
rect 24894 31297 24906 31300
rect 24848 31291 24906 31297
rect 25130 31288 25136 31300
rect 25188 31288 25194 31340
rect 26160 31328 26188 31436
rect 26789 31433 26801 31436
rect 26835 31464 26847 31467
rect 27614 31464 27620 31476
rect 26835 31436 27620 31464
rect 26835 31433 26847 31436
rect 26789 31427 26847 31433
rect 27614 31424 27620 31436
rect 27672 31424 27678 31476
rect 28258 31424 28264 31476
rect 28316 31464 28322 31476
rect 28810 31464 28816 31476
rect 28316 31436 28816 31464
rect 28316 31424 28322 31436
rect 28810 31424 28816 31436
rect 28868 31464 28874 31476
rect 29457 31467 29515 31473
rect 29457 31464 29469 31467
rect 28868 31436 29469 31464
rect 28868 31424 28874 31436
rect 29457 31433 29469 31436
rect 29503 31433 29515 31467
rect 29457 31427 29515 31433
rect 30834 31424 30840 31476
rect 30892 31464 30898 31476
rect 31389 31467 31447 31473
rect 31389 31464 31401 31467
rect 30892 31436 31401 31464
rect 30892 31424 30898 31436
rect 31389 31433 31401 31436
rect 31435 31433 31447 31467
rect 31389 31427 31447 31433
rect 33778 31424 33784 31476
rect 33836 31464 33842 31476
rect 33965 31467 34023 31473
rect 33965 31464 33977 31467
rect 33836 31436 33977 31464
rect 33836 31424 33842 31436
rect 33965 31433 33977 31436
rect 34011 31433 34023 31467
rect 33965 31427 34023 31433
rect 27430 31356 27436 31408
rect 27488 31396 27494 31408
rect 30276 31399 30334 31405
rect 27488 31368 29684 31396
rect 27488 31356 27494 31368
rect 26237 31331 26295 31337
rect 26237 31328 26249 31331
rect 26160 31300 26249 31328
rect 26237 31297 26249 31300
rect 26283 31297 26295 31331
rect 26237 31291 26295 31297
rect 26329 31331 26387 31337
rect 26329 31297 26341 31331
rect 26375 31297 26387 31331
rect 26329 31291 26387 31297
rect 21315 31232 22876 31260
rect 22925 31263 22983 31269
rect 21315 31229 21327 31232
rect 21269 31223 21327 31229
rect 22925 31229 22937 31263
rect 22971 31260 22983 31263
rect 23293 31263 23351 31269
rect 23293 31260 23305 31263
rect 22971 31232 23305 31260
rect 22971 31229 22983 31232
rect 22925 31223 22983 31229
rect 23293 31229 23305 31232
rect 23339 31260 23351 31263
rect 23382 31260 23388 31272
rect 23339 31232 23388 31260
rect 23339 31229 23351 31232
rect 23293 31223 23351 31229
rect 23382 31220 23388 31232
rect 23440 31220 23446 31272
rect 23566 31220 23572 31272
rect 23624 31220 23630 31272
rect 24394 31220 24400 31272
rect 24452 31260 24458 31272
rect 24581 31263 24639 31269
rect 24581 31260 24593 31263
rect 24452 31232 24593 31260
rect 24452 31220 24458 31232
rect 24581 31229 24593 31232
rect 24627 31229 24639 31263
rect 26344 31260 26372 31291
rect 26510 31288 26516 31340
rect 26568 31288 26574 31340
rect 26605 31331 26663 31337
rect 26605 31297 26617 31331
rect 26651 31328 26663 31331
rect 26786 31328 26792 31340
rect 26651 31300 26792 31328
rect 26651 31297 26663 31300
rect 26605 31291 26663 31297
rect 26786 31288 26792 31300
rect 26844 31288 26850 31340
rect 28092 31337 28120 31368
rect 29656 31340 29684 31368
rect 30276 31365 30288 31399
rect 30322 31396 30334 31399
rect 30374 31396 30380 31408
rect 30322 31368 30380 31396
rect 30322 31365 30334 31368
rect 30276 31359 30334 31365
rect 30374 31356 30380 31368
rect 30432 31356 30438 31408
rect 34333 31399 34391 31405
rect 34333 31365 34345 31399
rect 34379 31396 34391 31399
rect 34379 31368 34560 31396
rect 34379 31365 34391 31368
rect 34333 31359 34391 31365
rect 34532 31340 34560 31368
rect 34790 31356 34796 31408
rect 34848 31356 34854 31408
rect 28350 31337 28356 31340
rect 28077 31331 28135 31337
rect 28077 31297 28089 31331
rect 28123 31297 28135 31331
rect 28077 31291 28135 31297
rect 28344 31291 28356 31337
rect 28350 31288 28356 31291
rect 28408 31288 28414 31340
rect 29638 31288 29644 31340
rect 29696 31328 29702 31340
rect 30009 31331 30067 31337
rect 30009 31328 30021 31331
rect 29696 31300 30021 31328
rect 29696 31288 29702 31300
rect 30009 31297 30021 31300
rect 30055 31297 30067 31331
rect 30009 31291 30067 31297
rect 34149 31331 34207 31337
rect 34149 31297 34161 31331
rect 34195 31297 34207 31331
rect 34149 31291 34207 31297
rect 24581 31223 24639 31229
rect 25976 31232 26372 31260
rect 17681 31127 17739 31133
rect 17681 31093 17693 31127
rect 17727 31124 17739 31127
rect 17862 31124 17868 31136
rect 17727 31096 17868 31124
rect 17727 31093 17739 31096
rect 17681 31087 17739 31093
rect 17862 31084 17868 31096
rect 17920 31084 17926 31136
rect 19978 31084 19984 31136
rect 20036 31084 20042 31136
rect 23017 31127 23075 31133
rect 23017 31093 23029 31127
rect 23063 31124 23075 31127
rect 23290 31124 23296 31136
rect 23063 31096 23296 31124
rect 23063 31093 23075 31096
rect 23017 31087 23075 31093
rect 23290 31084 23296 31096
rect 23348 31084 23354 31136
rect 23584 31124 23612 31220
rect 25976 31136 26004 31232
rect 25222 31124 25228 31136
rect 23584 31096 25228 31124
rect 25222 31084 25228 31096
rect 25280 31084 25286 31136
rect 25958 31084 25964 31136
rect 26016 31084 26022 31136
rect 26786 31084 26792 31136
rect 26844 31124 26850 31136
rect 26973 31127 27031 31133
rect 26973 31124 26985 31127
rect 26844 31096 26985 31124
rect 26844 31084 26850 31096
rect 26973 31093 26985 31096
rect 27019 31093 27031 31127
rect 26973 31087 27031 31093
rect 27062 31084 27068 31136
rect 27120 31124 27126 31136
rect 34164 31124 34192 31291
rect 34422 31288 34428 31340
rect 34480 31288 34486 31340
rect 34514 31288 34520 31340
rect 34572 31288 34578 31340
rect 27120 31096 34192 31124
rect 27120 31084 27126 31096
rect 1104 31034 35328 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 35328 31034
rect 1104 30960 35328 30982
rect 3970 30880 3976 30932
rect 4028 30880 4034 30932
rect 6270 30880 6276 30932
rect 6328 30880 6334 30932
rect 7558 30880 7564 30932
rect 7616 30920 7622 30932
rect 23382 30920 23388 30932
rect 7616 30892 23388 30920
rect 7616 30880 7622 30892
rect 23382 30880 23388 30892
rect 23440 30880 23446 30932
rect 23474 30880 23480 30932
rect 23532 30920 23538 30932
rect 23934 30920 23940 30932
rect 23532 30892 23940 30920
rect 23532 30880 23538 30892
rect 23934 30880 23940 30892
rect 23992 30920 23998 30932
rect 23992 30892 24808 30920
rect 23992 30880 23998 30892
rect 5445 30855 5503 30861
rect 5445 30821 5457 30855
rect 5491 30852 5503 30855
rect 10870 30852 10876 30864
rect 5491 30824 10876 30852
rect 5491 30821 5503 30824
rect 5445 30815 5503 30821
rect 10870 30812 10876 30824
rect 10928 30812 10934 30864
rect 15654 30812 15660 30864
rect 15712 30852 15718 30864
rect 15933 30855 15991 30861
rect 15933 30852 15945 30855
rect 15712 30824 15945 30852
rect 15712 30812 15718 30824
rect 15933 30821 15945 30824
rect 15979 30852 15991 30855
rect 16114 30852 16120 30864
rect 15979 30824 16120 30852
rect 15979 30821 15991 30824
rect 15933 30815 15991 30821
rect 16114 30812 16120 30824
rect 16172 30812 16178 30864
rect 18322 30812 18328 30864
rect 18380 30852 18386 30864
rect 18601 30855 18659 30861
rect 18601 30852 18613 30855
rect 18380 30824 18613 30852
rect 18380 30812 18386 30824
rect 18601 30821 18613 30824
rect 18647 30821 18659 30855
rect 18601 30815 18659 30821
rect 4614 30744 4620 30796
rect 4672 30744 4678 30796
rect 6730 30744 6736 30796
rect 6788 30744 6794 30796
rect 6825 30787 6883 30793
rect 6825 30753 6837 30787
rect 6871 30784 6883 30787
rect 18616 30784 18644 30815
rect 19242 30812 19248 30864
rect 19300 30812 19306 30864
rect 19794 30784 19800 30796
rect 6871 30756 7604 30784
rect 18616 30756 19800 30784
rect 6871 30753 6883 30756
rect 6825 30747 6883 30753
rect 4433 30719 4491 30725
rect 4433 30685 4445 30719
rect 4479 30716 4491 30719
rect 4706 30716 4712 30728
rect 4479 30688 4712 30716
rect 4479 30685 4491 30688
rect 4433 30679 4491 30685
rect 4706 30676 4712 30688
rect 4764 30676 4770 30728
rect 4798 30676 4804 30728
rect 4856 30676 4862 30728
rect 4890 30676 4896 30728
rect 4948 30716 4954 30728
rect 4948 30688 4993 30716
rect 4948 30676 4954 30688
rect 5166 30676 5172 30728
rect 5224 30676 5230 30728
rect 5307 30719 5365 30725
rect 5307 30685 5319 30719
rect 5353 30716 5365 30719
rect 6641 30719 6699 30725
rect 5353 30688 6592 30716
rect 5353 30685 5365 30688
rect 5307 30679 5365 30685
rect 4341 30651 4399 30657
rect 4341 30617 4353 30651
rect 4387 30648 4399 30651
rect 4908 30648 4936 30676
rect 4387 30620 4936 30648
rect 5077 30651 5135 30657
rect 4387 30617 4399 30620
rect 4341 30611 4399 30617
rect 5077 30617 5089 30651
rect 5123 30617 5135 30651
rect 5077 30611 5135 30617
rect 5092 30580 5120 30611
rect 5629 30583 5687 30589
rect 5629 30580 5641 30583
rect 5092 30552 5641 30580
rect 5629 30549 5641 30552
rect 5675 30580 5687 30583
rect 5810 30580 5816 30592
rect 5675 30552 5816 30580
rect 5675 30549 5687 30552
rect 5629 30543 5687 30549
rect 5810 30540 5816 30552
rect 5868 30540 5874 30592
rect 6564 30580 6592 30688
rect 6641 30685 6653 30719
rect 6687 30716 6699 30719
rect 6914 30716 6920 30728
rect 6687 30688 6920 30716
rect 6687 30685 6699 30688
rect 6641 30679 6699 30685
rect 6914 30676 6920 30688
rect 6972 30676 6978 30728
rect 7466 30648 7472 30660
rect 6932 30620 7472 30648
rect 6932 30580 6960 30620
rect 7466 30608 7472 30620
rect 7524 30608 7530 30660
rect 6564 30552 6960 30580
rect 7193 30583 7251 30589
rect 7193 30549 7205 30583
rect 7239 30580 7251 30583
rect 7576 30580 7604 30756
rect 19794 30744 19800 30756
rect 19852 30744 19858 30796
rect 19889 30787 19947 30793
rect 19889 30753 19901 30787
rect 19935 30784 19947 30787
rect 19935 30756 20208 30784
rect 19935 30753 19947 30756
rect 19889 30747 19947 30753
rect 11330 30676 11336 30728
rect 11388 30716 11394 30728
rect 12253 30719 12311 30725
rect 12253 30716 12265 30719
rect 11388 30688 12265 30716
rect 11388 30676 11394 30688
rect 12253 30685 12265 30688
rect 12299 30685 12311 30719
rect 12253 30679 12311 30685
rect 12894 30676 12900 30728
rect 12952 30716 12958 30728
rect 13262 30716 13268 30728
rect 12952 30688 13268 30716
rect 12952 30676 12958 30688
rect 13262 30676 13268 30688
rect 13320 30716 13326 30728
rect 13817 30719 13875 30725
rect 13817 30716 13829 30719
rect 13320 30688 13829 30716
rect 13320 30676 13326 30688
rect 13817 30685 13829 30688
rect 13863 30685 13875 30719
rect 13817 30679 13875 30685
rect 14093 30719 14151 30725
rect 14093 30685 14105 30719
rect 14139 30716 14151 30719
rect 15102 30716 15108 30728
rect 14139 30688 15108 30716
rect 14139 30685 14151 30688
rect 14093 30679 14151 30685
rect 15102 30676 15108 30688
rect 15160 30676 15166 30728
rect 15286 30676 15292 30728
rect 15344 30716 15350 30728
rect 15470 30716 15476 30728
rect 15344 30688 15476 30716
rect 15344 30676 15350 30688
rect 15470 30676 15476 30688
rect 15528 30676 15534 30728
rect 15565 30719 15623 30725
rect 15565 30685 15577 30719
rect 15611 30685 15623 30719
rect 15565 30679 15623 30685
rect 19613 30719 19671 30725
rect 19613 30685 19625 30719
rect 19659 30716 19671 30719
rect 19978 30716 19984 30728
rect 19659 30688 19984 30716
rect 19659 30685 19671 30688
rect 19613 30679 19671 30685
rect 12520 30651 12578 30657
rect 12520 30617 12532 30651
rect 12566 30648 12578 30651
rect 12802 30648 12808 30660
rect 12566 30620 12808 30648
rect 12566 30617 12578 30620
rect 12520 30611 12578 30617
rect 12802 30608 12808 30620
rect 12860 30608 12866 30660
rect 14360 30651 14418 30657
rect 13556 30620 13860 30648
rect 10318 30580 10324 30592
rect 7239 30552 10324 30580
rect 7239 30549 7251 30552
rect 7193 30543 7251 30549
rect 10318 30540 10324 30552
rect 10376 30540 10382 30592
rect 10410 30540 10416 30592
rect 10468 30580 10474 30592
rect 13556 30580 13584 30620
rect 10468 30552 13584 30580
rect 10468 30540 10474 30552
rect 13630 30540 13636 30592
rect 13688 30540 13694 30592
rect 13832 30580 13860 30620
rect 14360 30617 14372 30651
rect 14406 30648 14418 30651
rect 14550 30648 14556 30660
rect 14406 30620 14556 30648
rect 14406 30617 14418 30620
rect 14360 30611 14418 30617
rect 14550 30608 14556 30620
rect 14608 30608 14614 30660
rect 15580 30648 15608 30679
rect 19978 30676 19984 30688
rect 20036 30676 20042 30728
rect 14660 30620 15608 30648
rect 14660 30580 14688 30620
rect 13832 30552 14688 30580
rect 15473 30583 15531 30589
rect 15473 30549 15485 30583
rect 15519 30580 15531 30583
rect 15562 30580 15568 30592
rect 15519 30552 15568 30580
rect 15519 30549 15531 30552
rect 15473 30543 15531 30549
rect 15562 30540 15568 30552
rect 15620 30540 15626 30592
rect 15746 30540 15752 30592
rect 15804 30540 15810 30592
rect 17586 30540 17592 30592
rect 17644 30540 17650 30592
rect 19702 30540 19708 30592
rect 19760 30540 19766 30592
rect 20180 30589 20208 30756
rect 20441 30719 20499 30725
rect 20441 30685 20453 30719
rect 20487 30716 20499 30719
rect 21818 30716 21824 30728
rect 20487 30688 21824 30716
rect 20487 30685 20499 30688
rect 20441 30679 20499 30685
rect 21818 30676 21824 30688
rect 21876 30716 21882 30728
rect 22281 30719 22339 30725
rect 22281 30716 22293 30719
rect 21876 30688 22293 30716
rect 21876 30676 21882 30688
rect 22281 30685 22293 30688
rect 22327 30685 22339 30719
rect 22281 30679 22339 30685
rect 23658 30676 23664 30728
rect 23716 30716 23722 30728
rect 24780 30725 24808 30892
rect 25130 30880 25136 30932
rect 25188 30880 25194 30932
rect 25222 30880 25228 30932
rect 25280 30920 25286 30932
rect 27522 30920 27528 30932
rect 25280 30892 27528 30920
rect 25280 30880 25286 30892
rect 27522 30880 27528 30892
rect 27580 30880 27586 30932
rect 28350 30880 28356 30932
rect 28408 30920 28414 30932
rect 28445 30923 28503 30929
rect 28445 30920 28457 30923
rect 28408 30892 28457 30920
rect 28408 30880 28414 30892
rect 28445 30889 28457 30892
rect 28491 30889 28503 30923
rect 31757 30923 31815 30929
rect 31757 30920 31769 30923
rect 28445 30883 28503 30889
rect 31588 30892 31769 30920
rect 25041 30855 25099 30861
rect 25041 30821 25053 30855
rect 25087 30852 25099 30855
rect 25866 30852 25872 30864
rect 25087 30824 25872 30852
rect 25087 30821 25099 30824
rect 25041 30815 25099 30821
rect 25866 30812 25872 30824
rect 25924 30812 25930 30864
rect 31588 30861 31616 30892
rect 31757 30889 31769 30892
rect 31803 30889 31815 30923
rect 31757 30883 31815 30889
rect 31389 30855 31447 30861
rect 28276 30824 29040 30852
rect 25314 30744 25320 30796
rect 25372 30784 25378 30796
rect 28276 30793 28304 30824
rect 25685 30787 25743 30793
rect 25685 30784 25697 30787
rect 25372 30756 25697 30784
rect 25372 30744 25378 30756
rect 25685 30753 25697 30756
rect 25731 30784 25743 30787
rect 28261 30787 28319 30793
rect 28261 30784 28273 30787
rect 25731 30756 28273 30784
rect 25731 30753 25743 30756
rect 25685 30747 25743 30753
rect 28261 30753 28273 30756
rect 28307 30753 28319 30787
rect 28261 30747 28319 30753
rect 28902 30744 28908 30796
rect 28960 30744 28966 30796
rect 29012 30793 29040 30824
rect 31389 30821 31401 30855
rect 31435 30852 31447 30855
rect 31573 30855 31631 30861
rect 31573 30852 31585 30855
rect 31435 30824 31585 30852
rect 31435 30821 31447 30824
rect 31389 30815 31447 30821
rect 31573 30821 31585 30824
rect 31619 30821 31631 30855
rect 31573 30815 31631 30821
rect 28997 30787 29055 30793
rect 28997 30753 29009 30787
rect 29043 30753 29055 30787
rect 28997 30747 29055 30753
rect 30282 30744 30288 30796
rect 30340 30784 30346 30796
rect 30745 30787 30803 30793
rect 30745 30784 30757 30787
rect 30340 30756 30757 30784
rect 30340 30744 30346 30756
rect 30745 30753 30757 30756
rect 30791 30784 30803 30787
rect 31404 30784 31432 30815
rect 30791 30756 31432 30784
rect 30791 30753 30803 30756
rect 30745 30747 30803 30753
rect 24397 30719 24455 30725
rect 24397 30716 24409 30719
rect 23716 30688 24409 30716
rect 23716 30676 23722 30688
rect 24397 30685 24409 30688
rect 24443 30685 24455 30719
rect 24397 30679 24455 30685
rect 24490 30719 24548 30725
rect 24490 30685 24502 30719
rect 24536 30685 24548 30719
rect 24490 30679 24548 30685
rect 24765 30719 24823 30725
rect 24765 30685 24777 30719
rect 24811 30685 24823 30719
rect 24765 30679 24823 30685
rect 20686 30651 20744 30657
rect 20686 30617 20698 30651
rect 20732 30617 20744 30651
rect 20686 30611 20744 30617
rect 22548 30651 22606 30657
rect 22548 30617 22560 30651
rect 22594 30648 22606 30651
rect 22830 30648 22836 30660
rect 22594 30620 22836 30648
rect 22594 30617 22606 30620
rect 22548 30611 22606 30617
rect 20165 30583 20223 30589
rect 20165 30549 20177 30583
rect 20211 30580 20223 30583
rect 20530 30580 20536 30592
rect 20211 30552 20536 30580
rect 20211 30549 20223 30552
rect 20165 30543 20223 30549
rect 20530 30540 20536 30552
rect 20588 30540 20594 30592
rect 20712 30580 20740 30611
rect 22830 30608 22836 30620
rect 22888 30608 22894 30660
rect 20806 30580 20812 30592
rect 20712 30552 20812 30580
rect 20806 30540 20812 30552
rect 20864 30540 20870 30592
rect 21266 30540 21272 30592
rect 21324 30580 21330 30592
rect 21821 30583 21879 30589
rect 21821 30580 21833 30583
rect 21324 30552 21833 30580
rect 21324 30540 21330 30552
rect 21821 30549 21833 30552
rect 21867 30549 21879 30583
rect 21821 30543 21879 30549
rect 23198 30540 23204 30592
rect 23256 30580 23262 30592
rect 23661 30583 23719 30589
rect 23661 30580 23673 30583
rect 23256 30552 23673 30580
rect 23256 30540 23262 30552
rect 23661 30549 23673 30552
rect 23707 30580 23719 30583
rect 24504 30580 24532 30679
rect 24854 30676 24860 30728
rect 24912 30725 24918 30728
rect 24912 30716 24920 30725
rect 25501 30719 25559 30725
rect 24912 30688 24957 30716
rect 24912 30679 24920 30688
rect 25501 30685 25513 30719
rect 25547 30716 25559 30719
rect 25958 30716 25964 30728
rect 25547 30688 25964 30716
rect 25547 30685 25559 30688
rect 25501 30679 25559 30685
rect 24912 30676 24918 30679
rect 25958 30676 25964 30688
rect 26016 30676 26022 30728
rect 28810 30676 28816 30728
rect 28868 30676 28874 30728
rect 29270 30676 29276 30728
rect 29328 30716 29334 30728
rect 30377 30719 30435 30725
rect 30377 30716 30389 30719
rect 29328 30688 30389 30716
rect 29328 30676 29334 30688
rect 30377 30685 30389 30688
rect 30423 30685 30435 30719
rect 30377 30679 30435 30685
rect 30561 30719 30619 30725
rect 30561 30685 30573 30719
rect 30607 30685 30619 30719
rect 30561 30679 30619 30685
rect 30653 30719 30711 30725
rect 30653 30685 30665 30719
rect 30699 30685 30711 30719
rect 30653 30679 30711 30685
rect 24670 30608 24676 30660
rect 24728 30608 24734 30660
rect 25593 30651 25651 30657
rect 25593 30617 25605 30651
rect 25639 30648 25651 30651
rect 25682 30648 25688 30660
rect 25639 30620 25688 30648
rect 25639 30617 25651 30620
rect 25593 30611 25651 30617
rect 25682 30608 25688 30620
rect 25740 30608 25746 30660
rect 25774 30608 25780 30660
rect 25832 30648 25838 30660
rect 26145 30651 26203 30657
rect 26145 30648 26157 30651
rect 25832 30620 26157 30648
rect 25832 30608 25838 30620
rect 26145 30617 26157 30620
rect 26191 30617 26203 30651
rect 26145 30611 26203 30617
rect 27982 30608 27988 30660
rect 28040 30648 28046 30660
rect 28040 30620 28396 30648
rect 28040 30608 28046 30620
rect 23707 30552 24532 30580
rect 23707 30549 23719 30552
rect 23661 30543 23719 30549
rect 24854 30540 24860 30592
rect 24912 30580 24918 30592
rect 25958 30580 25964 30592
rect 24912 30552 25964 30580
rect 24912 30540 24918 30552
rect 25958 30540 25964 30552
rect 26016 30540 26022 30592
rect 27614 30540 27620 30592
rect 27672 30580 27678 30592
rect 27890 30580 27896 30592
rect 27672 30552 27896 30580
rect 27672 30540 27678 30552
rect 27890 30540 27896 30552
rect 27948 30540 27954 30592
rect 28368 30580 28396 30620
rect 28994 30608 29000 30660
rect 29052 30648 29058 30660
rect 30576 30648 30604 30679
rect 29052 30620 30604 30648
rect 29052 30608 29058 30620
rect 30668 30580 30696 30679
rect 30834 30676 30840 30728
rect 30892 30716 30898 30728
rect 30929 30719 30987 30725
rect 30929 30716 30941 30719
rect 30892 30688 30941 30716
rect 30892 30676 30898 30688
rect 30929 30685 30941 30688
rect 30975 30685 30987 30719
rect 30929 30679 30987 30685
rect 31202 30676 31208 30728
rect 31260 30716 31266 30728
rect 31941 30719 31999 30725
rect 31941 30716 31953 30719
rect 31260 30688 31953 30716
rect 31260 30676 31266 30688
rect 31941 30685 31953 30688
rect 31987 30685 31999 30719
rect 31941 30679 31999 30685
rect 34057 30719 34115 30725
rect 34057 30685 34069 30719
rect 34103 30716 34115 30719
rect 34146 30716 34152 30728
rect 34103 30688 34152 30716
rect 34103 30685 34115 30688
rect 34057 30679 34115 30685
rect 34146 30676 34152 30688
rect 34204 30676 34210 30728
rect 31113 30651 31171 30657
rect 31113 30617 31125 30651
rect 31159 30648 31171 30651
rect 33042 30648 33048 30660
rect 31159 30620 33048 30648
rect 31159 30617 31171 30620
rect 31113 30611 31171 30617
rect 33042 30608 33048 30620
rect 33100 30608 33106 30660
rect 34333 30651 34391 30657
rect 34333 30617 34345 30651
rect 34379 30648 34391 30651
rect 34514 30648 34520 30660
rect 34379 30620 34520 30648
rect 34379 30617 34391 30620
rect 34333 30611 34391 30617
rect 34514 30608 34520 30620
rect 34572 30608 34578 30660
rect 28368 30552 30696 30580
rect 1104 30490 35328 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35328 30490
rect 1104 30416 35328 30438
rect 4614 30336 4620 30388
rect 4672 30336 4678 30388
rect 4798 30336 4804 30388
rect 4856 30336 4862 30388
rect 5169 30379 5227 30385
rect 5169 30345 5181 30379
rect 5215 30376 5227 30379
rect 5215 30348 12756 30376
rect 5215 30345 5227 30348
rect 5169 30339 5227 30345
rect 4632 30308 4660 30336
rect 4890 30308 4896 30320
rect 4632 30280 4896 30308
rect 4890 30268 4896 30280
rect 4948 30308 4954 30320
rect 5184 30308 5212 30339
rect 4948 30280 5212 30308
rect 4948 30268 4954 30280
rect 5350 30268 5356 30320
rect 5408 30308 5414 30320
rect 9214 30308 9220 30320
rect 5408 30280 9220 30308
rect 5408 30268 5414 30280
rect 9214 30268 9220 30280
rect 9272 30308 9278 30320
rect 9309 30311 9367 30317
rect 9309 30308 9321 30311
rect 9272 30280 9321 30308
rect 9272 30268 9278 30280
rect 9309 30277 9321 30280
rect 9355 30277 9367 30311
rect 9309 30271 9367 30277
rect 10505 30311 10563 30317
rect 10505 30277 10517 30311
rect 10551 30308 10563 30311
rect 11054 30308 11060 30320
rect 10551 30280 11060 30308
rect 10551 30277 10563 30280
rect 10505 30271 10563 30277
rect 1302 30200 1308 30252
rect 1360 30240 1366 30252
rect 1397 30243 1455 30249
rect 1397 30240 1409 30243
rect 1360 30212 1409 30240
rect 1360 30200 1366 30212
rect 1397 30209 1409 30212
rect 1443 30240 1455 30243
rect 1673 30243 1731 30249
rect 1673 30240 1685 30243
rect 1443 30212 1685 30240
rect 1443 30209 1455 30212
rect 1397 30203 1455 30209
rect 1673 30209 1685 30212
rect 1719 30209 1731 30243
rect 1673 30203 1731 30209
rect 3602 30200 3608 30252
rect 3660 30240 3666 30252
rect 4249 30243 4307 30249
rect 4249 30240 4261 30243
rect 3660 30212 4261 30240
rect 3660 30200 3666 30212
rect 4249 30209 4261 30212
rect 4295 30209 4307 30243
rect 4249 30203 4307 30209
rect 4433 30243 4491 30249
rect 4433 30209 4445 30243
rect 4479 30209 4491 30243
rect 4433 30203 4491 30209
rect 4525 30243 4583 30249
rect 4525 30209 4537 30243
rect 4571 30209 4583 30243
rect 4525 30203 4583 30209
rect 4617 30243 4675 30249
rect 4617 30209 4629 30243
rect 4663 30240 4675 30243
rect 5442 30240 5448 30252
rect 4663 30212 5448 30240
rect 4663 30209 4675 30212
rect 4617 30203 4675 30209
rect 1581 30039 1639 30045
rect 1581 30005 1593 30039
rect 1627 30036 1639 30039
rect 2866 30036 2872 30048
rect 1627 30008 2872 30036
rect 1627 30005 1639 30008
rect 1581 29999 1639 30005
rect 2866 29996 2872 30008
rect 2924 29996 2930 30048
rect 4448 30036 4476 30203
rect 4540 30104 4568 30203
rect 5442 30200 5448 30212
rect 5500 30240 5506 30252
rect 9401 30243 9459 30249
rect 5500 30212 9352 30240
rect 5500 30200 5506 30212
rect 9324 30184 9352 30212
rect 9401 30209 9413 30243
rect 9447 30240 9459 30243
rect 9766 30240 9772 30252
rect 9447 30212 9772 30240
rect 9447 30209 9459 30212
rect 9401 30203 9459 30209
rect 9766 30200 9772 30212
rect 9824 30240 9830 30252
rect 10321 30243 10379 30249
rect 10321 30240 10333 30243
rect 9824 30212 10333 30240
rect 9824 30200 9830 30212
rect 10321 30209 10333 30212
rect 10367 30209 10379 30243
rect 10321 30203 10379 30209
rect 9306 30132 9312 30184
rect 9364 30132 9370 30184
rect 9582 30132 9588 30184
rect 9640 30132 9646 30184
rect 10226 30132 10232 30184
rect 10284 30172 10290 30184
rect 10520 30172 10548 30271
rect 11054 30268 11060 30280
rect 11112 30268 11118 30320
rect 12728 30308 12756 30348
rect 12802 30336 12808 30388
rect 12860 30336 12866 30388
rect 14458 30376 14464 30388
rect 12912 30348 14464 30376
rect 12912 30308 12940 30348
rect 14458 30336 14464 30348
rect 14516 30336 14522 30388
rect 14550 30336 14556 30388
rect 14608 30336 14614 30388
rect 15013 30379 15071 30385
rect 15013 30345 15025 30379
rect 15059 30376 15071 30379
rect 15286 30376 15292 30388
rect 15059 30348 15292 30376
rect 15059 30345 15071 30348
rect 15013 30339 15071 30345
rect 15286 30336 15292 30348
rect 15344 30376 15350 30388
rect 15746 30376 15752 30388
rect 15344 30348 15752 30376
rect 15344 30336 15350 30348
rect 15746 30336 15752 30348
rect 15804 30336 15810 30388
rect 16298 30336 16304 30388
rect 16356 30376 16362 30388
rect 19337 30379 19395 30385
rect 16356 30348 18460 30376
rect 16356 30336 16362 30348
rect 12728 30280 12940 30308
rect 13078 30268 13084 30320
rect 13136 30308 13142 30320
rect 13173 30311 13231 30317
rect 13173 30308 13185 30311
rect 13136 30280 13185 30308
rect 13136 30268 13142 30280
rect 13173 30277 13185 30280
rect 13219 30277 13231 30311
rect 13173 30271 13231 30277
rect 13265 30311 13323 30317
rect 13265 30277 13277 30311
rect 13311 30308 13323 30311
rect 13630 30308 13636 30320
rect 13311 30280 13636 30308
rect 13311 30277 13323 30280
rect 13265 30271 13323 30277
rect 13630 30268 13636 30280
rect 13688 30308 13694 30320
rect 13909 30311 13967 30317
rect 13909 30308 13921 30311
rect 13688 30280 13921 30308
rect 13688 30268 13694 30280
rect 13909 30277 13921 30280
rect 13955 30277 13967 30311
rect 13909 30271 13967 30277
rect 14001 30311 14059 30317
rect 14001 30277 14013 30311
rect 14047 30308 14059 30311
rect 14274 30308 14280 30320
rect 14047 30280 14280 30308
rect 14047 30277 14059 30280
rect 14001 30271 14059 30277
rect 14274 30268 14280 30280
rect 14332 30268 14338 30320
rect 14921 30311 14979 30317
rect 14921 30277 14933 30311
rect 14967 30308 14979 30311
rect 14967 30280 15608 30308
rect 14967 30277 14979 30280
rect 14921 30271 14979 30277
rect 15580 30252 15608 30280
rect 18138 30268 18144 30320
rect 18196 30308 18202 30320
rect 18325 30311 18383 30317
rect 18325 30308 18337 30311
rect 18196 30280 18337 30308
rect 18196 30268 18202 30280
rect 18325 30277 18337 30280
rect 18371 30277 18383 30311
rect 18325 30271 18383 30277
rect 18432 30252 18460 30348
rect 19337 30345 19349 30379
rect 19383 30376 19395 30379
rect 19702 30376 19708 30388
rect 19383 30348 19708 30376
rect 19383 30345 19395 30348
rect 19337 30339 19395 30345
rect 19702 30336 19708 30348
rect 19760 30336 19766 30388
rect 20806 30336 20812 30388
rect 20864 30336 20870 30388
rect 21266 30336 21272 30388
rect 21324 30336 21330 30388
rect 22830 30336 22836 30388
rect 22888 30336 22894 30388
rect 23198 30336 23204 30388
rect 23256 30336 23262 30388
rect 24670 30336 24676 30388
rect 24728 30376 24734 30388
rect 25774 30376 25780 30388
rect 24728 30348 25780 30376
rect 24728 30336 24734 30348
rect 25774 30336 25780 30348
rect 25832 30336 25838 30388
rect 27893 30379 27951 30385
rect 27893 30345 27905 30379
rect 27939 30345 27951 30379
rect 27893 30339 27951 30345
rect 18506 30268 18512 30320
rect 18564 30308 18570 30320
rect 20898 30308 20904 30320
rect 18564 30280 20904 30308
rect 18564 30268 18570 30280
rect 20898 30268 20904 30280
rect 20956 30268 20962 30320
rect 21174 30268 21180 30320
rect 21232 30268 21238 30320
rect 24486 30308 24492 30320
rect 21284 30280 24492 30308
rect 10594 30200 10600 30252
rect 10652 30200 10658 30252
rect 10686 30200 10692 30252
rect 10744 30240 10750 30252
rect 11149 30243 11207 30249
rect 11149 30240 11161 30243
rect 10744 30212 11161 30240
rect 10744 30200 10750 30212
rect 11149 30209 11161 30212
rect 11195 30240 11207 30243
rect 11882 30240 11888 30252
rect 11195 30212 11888 30240
rect 11195 30209 11207 30212
rect 11149 30203 11207 30209
rect 11882 30200 11888 30212
rect 11940 30200 11946 30252
rect 12710 30200 12716 30252
rect 12768 30240 12774 30252
rect 13817 30243 13875 30249
rect 13817 30240 13829 30243
rect 12768 30212 13829 30240
rect 12768 30200 12774 30212
rect 13817 30209 13829 30212
rect 13863 30209 13875 30243
rect 13817 30203 13875 30209
rect 10284 30144 10548 30172
rect 10796 30144 12434 30172
rect 10284 30132 10290 30144
rect 4614 30104 4620 30116
rect 4540 30076 4620 30104
rect 4614 30064 4620 30076
rect 4672 30064 4678 30116
rect 9030 30064 9036 30116
rect 9088 30104 9094 30116
rect 10796 30104 10824 30144
rect 9088 30076 10824 30104
rect 10873 30107 10931 30113
rect 9088 30064 9094 30076
rect 10873 30073 10885 30107
rect 10919 30104 10931 30107
rect 11238 30104 11244 30116
rect 10919 30076 11244 30104
rect 10919 30073 10931 30076
rect 10873 30067 10931 30073
rect 11238 30064 11244 30076
rect 11296 30064 11302 30116
rect 4798 30036 4804 30048
rect 4448 30008 4804 30036
rect 4798 29996 4804 30008
rect 4856 30036 4862 30048
rect 4893 30039 4951 30045
rect 4893 30036 4905 30039
rect 4856 30008 4905 30036
rect 4856 29996 4862 30008
rect 4893 30005 4905 30008
rect 4939 30005 4951 30039
rect 4893 29999 4951 30005
rect 8938 29996 8944 30048
rect 8996 29996 9002 30048
rect 9582 29996 9588 30048
rect 9640 30036 9646 30048
rect 9861 30039 9919 30045
rect 9861 30036 9873 30039
rect 9640 30008 9873 30036
rect 9640 29996 9646 30008
rect 9861 30005 9873 30008
rect 9907 30036 9919 30039
rect 11054 30036 11060 30048
rect 9907 30008 11060 30036
rect 9907 30005 9919 30008
rect 9861 29999 9919 30005
rect 11054 29996 11060 30008
rect 11112 29996 11118 30048
rect 12406 30036 12434 30144
rect 13262 30132 13268 30184
rect 13320 30172 13326 30184
rect 13357 30175 13415 30181
rect 13357 30172 13369 30175
rect 13320 30144 13369 30172
rect 13320 30132 13326 30144
rect 13357 30141 13369 30144
rect 13403 30141 13415 30175
rect 13832 30172 13860 30203
rect 14090 30200 14096 30252
rect 14148 30240 14154 30252
rect 14185 30243 14243 30249
rect 14185 30240 14197 30243
rect 14148 30212 14197 30240
rect 14148 30200 14154 30212
rect 14185 30209 14197 30212
rect 14231 30209 14243 30243
rect 14185 30203 14243 30209
rect 15194 30200 15200 30252
rect 15252 30240 15258 30252
rect 15473 30243 15531 30249
rect 15473 30240 15485 30243
rect 15252 30212 15485 30240
rect 15252 30200 15258 30212
rect 15473 30209 15485 30212
rect 15519 30209 15531 30243
rect 15473 30203 15531 30209
rect 15562 30200 15568 30252
rect 15620 30240 15626 30252
rect 15749 30243 15807 30249
rect 15620 30212 15665 30240
rect 15620 30200 15626 30212
rect 15749 30209 15761 30243
rect 15795 30209 15807 30243
rect 15749 30203 15807 30209
rect 15105 30175 15163 30181
rect 13832 30144 14504 30172
rect 13357 30135 13415 30141
rect 13170 30064 13176 30116
rect 13228 30104 13234 30116
rect 13633 30107 13691 30113
rect 13633 30104 13645 30107
rect 13228 30076 13645 30104
rect 13228 30064 13234 30076
rect 13633 30073 13645 30076
rect 13679 30073 13691 30107
rect 13633 30067 13691 30073
rect 14274 30036 14280 30048
rect 12406 30008 14280 30036
rect 14274 29996 14280 30008
rect 14332 29996 14338 30048
rect 14476 30045 14504 30144
rect 15105 30141 15117 30175
rect 15151 30172 15163 30175
rect 15654 30172 15660 30184
rect 15151 30144 15660 30172
rect 15151 30141 15163 30144
rect 15105 30135 15163 30141
rect 15654 30132 15660 30144
rect 15712 30132 15718 30184
rect 15764 30172 15792 30203
rect 15838 30200 15844 30252
rect 15896 30200 15902 30252
rect 15979 30243 16037 30249
rect 15979 30209 15991 30243
rect 16025 30240 16037 30243
rect 16206 30240 16212 30252
rect 16025 30212 16212 30240
rect 16025 30209 16037 30212
rect 15979 30203 16037 30209
rect 16206 30200 16212 30212
rect 16264 30200 16270 30252
rect 18049 30243 18107 30249
rect 18049 30209 18061 30243
rect 18095 30209 18107 30243
rect 18049 30203 18107 30209
rect 18233 30243 18291 30249
rect 18233 30209 18245 30243
rect 18279 30240 18291 30243
rect 18279 30212 18368 30240
rect 18279 30209 18291 30212
rect 18233 30203 18291 30209
rect 16301 30175 16359 30181
rect 16301 30172 16313 30175
rect 15764 30144 16313 30172
rect 16301 30141 16313 30144
rect 16347 30172 16359 30175
rect 16574 30172 16580 30184
rect 16347 30144 16580 30172
rect 16347 30141 16359 30144
rect 16301 30135 16359 30141
rect 16574 30132 16580 30144
rect 16632 30172 16638 30184
rect 17034 30172 17040 30184
rect 16632 30144 17040 30172
rect 16632 30132 16638 30144
rect 17034 30132 17040 30144
rect 17092 30132 17098 30184
rect 16117 30107 16175 30113
rect 16117 30073 16129 30107
rect 16163 30104 16175 30107
rect 16850 30104 16856 30116
rect 16163 30076 16856 30104
rect 16163 30073 16175 30076
rect 16117 30067 16175 30073
rect 16850 30064 16856 30076
rect 16908 30064 16914 30116
rect 18064 30104 18092 30203
rect 18340 30172 18368 30212
rect 18414 30200 18420 30252
rect 18472 30200 18478 30252
rect 18877 30243 18935 30249
rect 18877 30209 18889 30243
rect 18923 30240 18935 30243
rect 21284 30240 21312 30280
rect 24486 30268 24492 30280
rect 24544 30268 24550 30320
rect 27908 30308 27936 30339
rect 28261 30311 28319 30317
rect 28261 30308 28273 30311
rect 26804 30280 28273 30308
rect 21913 30243 21971 30249
rect 21913 30240 21925 30243
rect 18923 30212 21312 30240
rect 21560 30212 21925 30240
rect 18923 30209 18935 30212
rect 18877 30203 18935 30209
rect 18892 30172 18920 30203
rect 18340 30144 18920 30172
rect 19153 30175 19211 30181
rect 19153 30141 19165 30175
rect 19199 30141 19211 30175
rect 19153 30135 19211 30141
rect 19245 30175 19303 30181
rect 19245 30141 19257 30175
rect 19291 30172 19303 30175
rect 20622 30172 20628 30184
rect 19291 30144 20628 30172
rect 19291 30141 19303 30144
rect 19245 30135 19303 30141
rect 18322 30104 18328 30116
rect 18064 30076 18328 30104
rect 18322 30064 18328 30076
rect 18380 30064 18386 30116
rect 18601 30107 18659 30113
rect 18601 30073 18613 30107
rect 18647 30104 18659 30107
rect 18690 30104 18696 30116
rect 18647 30076 18696 30104
rect 18647 30073 18659 30076
rect 18601 30067 18659 30073
rect 18690 30064 18696 30076
rect 18748 30064 18754 30116
rect 19168 30104 19196 30135
rect 20622 30132 20628 30144
rect 20680 30132 20686 30184
rect 21453 30175 21511 30181
rect 21453 30141 21465 30175
rect 21499 30172 21511 30175
rect 21560 30172 21588 30212
rect 21913 30209 21925 30212
rect 21959 30240 21971 30243
rect 23014 30240 23020 30252
rect 21959 30212 23020 30240
rect 21959 30209 21971 30212
rect 21913 30203 21971 30209
rect 23014 30200 23020 30212
rect 23072 30200 23078 30252
rect 26804 30240 26832 30280
rect 23400 30212 26832 30240
rect 26973 30243 27031 30249
rect 21499 30144 21588 30172
rect 21499 30141 21511 30144
rect 21453 30135 21511 30141
rect 21634 30132 21640 30184
rect 21692 30172 21698 30184
rect 21692 30144 22094 30172
rect 21692 30132 21698 30144
rect 21910 30104 21916 30116
rect 19168 30076 21916 30104
rect 21910 30064 21916 30076
rect 21968 30064 21974 30116
rect 22066 30104 22094 30144
rect 23290 30132 23296 30184
rect 23348 30132 23354 30184
rect 23400 30104 23428 30212
rect 26973 30209 26985 30243
rect 27019 30209 27031 30243
rect 26973 30203 27031 30209
rect 23477 30175 23535 30181
rect 23477 30141 23489 30175
rect 23523 30172 23535 30175
rect 26988 30172 27016 30203
rect 27062 30200 27068 30252
rect 27120 30200 27126 30252
rect 27249 30243 27307 30249
rect 27249 30209 27261 30243
rect 27295 30209 27307 30243
rect 27249 30203 27307 30209
rect 27154 30172 27160 30184
rect 23523 30144 23796 30172
rect 26988 30144 27160 30172
rect 23523 30141 23535 30144
rect 23477 30135 23535 30141
rect 22066 30076 23428 30104
rect 14461 30039 14519 30045
rect 14461 30005 14473 30039
rect 14507 30036 14519 30039
rect 14550 30036 14556 30048
rect 14507 30008 14556 30036
rect 14507 30005 14519 30008
rect 14461 29999 14519 30005
rect 14550 29996 14556 30008
rect 14608 29996 14614 30048
rect 16298 29996 16304 30048
rect 16356 30036 16362 30048
rect 16393 30039 16451 30045
rect 16393 30036 16405 30039
rect 16356 30008 16405 30036
rect 16356 29996 16362 30008
rect 16393 30005 16405 30008
rect 16439 30005 16451 30039
rect 16393 29999 16451 30005
rect 19334 29996 19340 30048
rect 19392 30036 19398 30048
rect 19705 30039 19763 30045
rect 19705 30036 19717 30039
rect 19392 30008 19717 30036
rect 19392 29996 19398 30008
rect 19705 30005 19717 30008
rect 19751 30005 19763 30039
rect 19705 29999 19763 30005
rect 20714 29996 20720 30048
rect 20772 30036 20778 30048
rect 23768 30045 23796 30144
rect 27154 30132 27160 30144
rect 27212 30132 27218 30184
rect 24486 30064 24492 30116
rect 24544 30104 24550 30116
rect 26697 30107 26755 30113
rect 26697 30104 26709 30107
rect 24544 30076 26709 30104
rect 24544 30064 24550 30076
rect 26697 30073 26709 30076
rect 26743 30104 26755 30107
rect 27264 30104 27292 30203
rect 27338 30200 27344 30252
rect 27396 30200 27402 30252
rect 27448 30249 27476 30280
rect 28261 30277 28273 30280
rect 28307 30308 28319 30311
rect 28445 30311 28503 30317
rect 28445 30308 28457 30311
rect 28307 30280 28457 30308
rect 28307 30277 28319 30280
rect 28261 30271 28319 30277
rect 28445 30277 28457 30280
rect 28491 30277 28503 30311
rect 28445 30271 28503 30277
rect 33965 30311 34023 30317
rect 33965 30277 33977 30311
rect 34011 30308 34023 30311
rect 34146 30308 34152 30320
rect 34011 30280 34152 30308
rect 34011 30277 34023 30280
rect 33965 30271 34023 30277
rect 34146 30268 34152 30280
rect 34204 30268 34210 30320
rect 27438 30243 27496 30249
rect 27438 30209 27450 30243
rect 27484 30209 27496 30243
rect 27709 30243 27767 30249
rect 27709 30240 27721 30243
rect 27438 30203 27496 30209
rect 27540 30212 27721 30240
rect 27540 30104 27568 30212
rect 27709 30209 27721 30212
rect 27755 30240 27767 30243
rect 28077 30243 28135 30249
rect 28077 30240 28089 30243
rect 27755 30212 28089 30240
rect 27755 30209 27767 30212
rect 27709 30203 27767 30209
rect 28077 30209 28089 30212
rect 28123 30209 28135 30243
rect 28077 30203 28135 30209
rect 29273 30243 29331 30249
rect 29273 30209 29285 30243
rect 29319 30240 29331 30243
rect 29319 30212 29684 30240
rect 29319 30209 29331 30212
rect 29273 30203 29331 30209
rect 26743 30076 27292 30104
rect 27448 30076 27568 30104
rect 27617 30107 27675 30113
rect 26743 30073 26755 30076
rect 26697 30067 26755 30073
rect 23753 30039 23811 30045
rect 23753 30036 23765 30039
rect 20772 30008 23765 30036
rect 20772 29996 20778 30008
rect 23753 30005 23765 30008
rect 23799 30036 23811 30039
rect 24026 30036 24032 30048
rect 23799 30008 24032 30036
rect 23799 30005 23811 30008
rect 23753 29999 23811 30005
rect 24026 29996 24032 30008
rect 24084 29996 24090 30048
rect 25041 30039 25099 30045
rect 25041 30005 25053 30039
rect 25087 30036 25099 30039
rect 25314 30036 25320 30048
rect 25087 30008 25320 30036
rect 25087 30005 25099 30008
rect 25041 29999 25099 30005
rect 25314 29996 25320 30008
rect 25372 29996 25378 30048
rect 25590 29996 25596 30048
rect 25648 30036 25654 30048
rect 26050 30036 26056 30048
rect 25648 30008 26056 30036
rect 25648 29996 25654 30008
rect 26050 29996 26056 30008
rect 26108 30036 26114 30048
rect 27448 30036 27476 30076
rect 27617 30073 27629 30107
rect 27663 30104 27675 30107
rect 28994 30104 29000 30116
rect 27663 30076 29000 30104
rect 27663 30073 27675 30076
rect 27617 30067 27675 30073
rect 28994 30064 29000 30076
rect 29052 30064 29058 30116
rect 26108 30008 27476 30036
rect 26108 29996 26114 30008
rect 27522 29996 27528 30048
rect 27580 30036 27586 30048
rect 29086 30036 29092 30048
rect 27580 30008 29092 30036
rect 27580 29996 27586 30008
rect 29086 29996 29092 30008
rect 29144 30036 29150 30048
rect 29656 30045 29684 30212
rect 33042 30200 33048 30252
rect 33100 30240 33106 30252
rect 33781 30243 33839 30249
rect 33781 30240 33793 30243
rect 33100 30212 33793 30240
rect 33100 30200 33106 30212
rect 33781 30209 33793 30212
rect 33827 30209 33839 30243
rect 33781 30203 33839 30209
rect 34057 30243 34115 30249
rect 34057 30209 34069 30243
rect 34103 30240 34115 30243
rect 34238 30240 34244 30252
rect 34103 30212 34244 30240
rect 34103 30209 34115 30212
rect 34057 30203 34115 30209
rect 34238 30200 34244 30212
rect 34296 30200 34302 30252
rect 34149 30175 34207 30181
rect 34149 30172 34161 30175
rect 33428 30144 34161 30172
rect 33428 30048 33456 30144
rect 34149 30141 34161 30144
rect 34195 30141 34207 30175
rect 34149 30135 34207 30141
rect 34425 30175 34483 30181
rect 34425 30141 34437 30175
rect 34471 30141 34483 30175
rect 34425 30135 34483 30141
rect 33502 30064 33508 30116
rect 33560 30104 33566 30116
rect 34440 30104 34468 30135
rect 33560 30076 34468 30104
rect 33560 30064 33566 30076
rect 29365 30039 29423 30045
rect 29365 30036 29377 30039
rect 29144 30008 29377 30036
rect 29144 29996 29150 30008
rect 29365 30005 29377 30008
rect 29411 30005 29423 30039
rect 29365 29999 29423 30005
rect 29641 30039 29699 30045
rect 29641 30005 29653 30039
rect 29687 30036 29699 30039
rect 30190 30036 30196 30048
rect 29687 30008 30196 30036
rect 29687 30005 29699 30008
rect 29641 29999 29699 30005
rect 30190 29996 30196 30008
rect 30248 29996 30254 30048
rect 33410 29996 33416 30048
rect 33468 29996 33474 30048
rect 33594 29996 33600 30048
rect 33652 29996 33658 30048
rect 1104 29946 35328 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 35328 29946
rect 1104 29872 35328 29894
rect 3602 29792 3608 29844
rect 3660 29792 3666 29844
rect 8754 29792 8760 29844
rect 8812 29792 8818 29844
rect 10594 29792 10600 29844
rect 10652 29832 10658 29844
rect 10965 29835 11023 29841
rect 10965 29832 10977 29835
rect 10652 29804 10977 29832
rect 10652 29792 10658 29804
rect 10965 29801 10977 29804
rect 11011 29801 11023 29835
rect 10965 29795 11023 29801
rect 11054 29792 11060 29844
rect 11112 29832 11118 29844
rect 11112 29804 12434 29832
rect 11112 29792 11118 29804
rect 5258 29656 5264 29708
rect 5316 29656 5322 29708
rect 9217 29699 9275 29705
rect 9217 29696 9229 29699
rect 8404 29668 9229 29696
rect 2222 29588 2228 29640
rect 2280 29628 2286 29640
rect 3789 29631 3847 29637
rect 3789 29628 3801 29631
rect 2280 29600 3801 29628
rect 2280 29588 2286 29600
rect 3789 29597 3801 29600
rect 3835 29628 3847 29631
rect 5276 29628 5304 29656
rect 8404 29637 8432 29668
rect 9217 29665 9229 29668
rect 9263 29665 9275 29699
rect 9217 29659 9275 29665
rect 6733 29631 6791 29637
rect 6733 29628 6745 29631
rect 3835 29600 6745 29628
rect 3835 29597 3847 29600
rect 3789 29591 3847 29597
rect 6733 29597 6745 29600
rect 6779 29597 6791 29631
rect 8205 29631 8263 29637
rect 8205 29628 8217 29631
rect 6733 29591 6791 29597
rect 6932 29600 8217 29628
rect 2492 29563 2550 29569
rect 2492 29529 2504 29563
rect 2538 29560 2550 29563
rect 3050 29560 3056 29572
rect 2538 29532 3056 29560
rect 2538 29529 2550 29532
rect 2492 29523 2550 29529
rect 3050 29520 3056 29532
rect 3108 29520 3114 29572
rect 4056 29563 4114 29569
rect 4056 29529 4068 29563
rect 4102 29560 4114 29563
rect 4246 29560 4252 29572
rect 4102 29532 4252 29560
rect 4102 29529 4114 29532
rect 4056 29523 4114 29529
rect 4246 29520 4252 29532
rect 4304 29520 4310 29572
rect 4522 29520 4528 29572
rect 4580 29560 4586 29572
rect 4890 29560 4896 29572
rect 4580 29532 4896 29560
rect 4580 29520 4586 29532
rect 4890 29520 4896 29532
rect 4948 29520 4954 29572
rect 5528 29563 5586 29569
rect 5528 29529 5540 29563
rect 5574 29560 5586 29563
rect 6270 29560 6276 29572
rect 5574 29532 6276 29560
rect 5574 29529 5586 29532
rect 5528 29523 5586 29529
rect 6270 29520 6276 29532
rect 6328 29520 6334 29572
rect 4614 29452 4620 29504
rect 4672 29492 4678 29504
rect 5169 29495 5227 29501
rect 5169 29492 5181 29495
rect 4672 29464 5181 29492
rect 4672 29452 4678 29464
rect 5169 29461 5181 29464
rect 5215 29461 5227 29495
rect 5169 29455 5227 29461
rect 6641 29495 6699 29501
rect 6641 29461 6653 29495
rect 6687 29492 6699 29495
rect 6730 29492 6736 29504
rect 6687 29464 6736 29492
rect 6687 29461 6699 29464
rect 6641 29455 6699 29461
rect 6730 29452 6736 29464
rect 6788 29492 6794 29504
rect 6932 29492 6960 29600
rect 8205 29597 8217 29600
rect 8251 29597 8263 29631
rect 8205 29591 8263 29597
rect 8389 29631 8447 29637
rect 8389 29597 8401 29631
rect 8435 29597 8447 29631
rect 8389 29591 8447 29597
rect 8570 29588 8576 29640
rect 8628 29628 8634 29640
rect 9030 29628 9036 29640
rect 8628 29600 9036 29628
rect 8628 29588 8634 29600
rect 9030 29588 9036 29600
rect 9088 29588 9094 29640
rect 7000 29563 7058 29569
rect 7000 29529 7012 29563
rect 7046 29560 7058 29563
rect 7374 29560 7380 29572
rect 7046 29532 7380 29560
rect 7046 29529 7058 29532
rect 7000 29523 7058 29529
rect 7374 29520 7380 29532
rect 7432 29520 7438 29572
rect 8481 29563 8539 29569
rect 8481 29529 8493 29563
rect 8527 29529 8539 29563
rect 8481 29523 8539 29529
rect 6788 29464 6960 29492
rect 6788 29452 6794 29464
rect 7742 29452 7748 29504
rect 7800 29492 7806 29504
rect 8113 29495 8171 29501
rect 8113 29492 8125 29495
rect 7800 29464 8125 29492
rect 7800 29452 7806 29464
rect 8113 29461 8125 29464
rect 8159 29492 8171 29495
rect 8496 29492 8524 29523
rect 8159 29464 8524 29492
rect 9232 29492 9260 29659
rect 11330 29656 11336 29708
rect 11388 29656 11394 29708
rect 12406 29696 12434 29804
rect 14366 29792 14372 29844
rect 14424 29792 14430 29844
rect 15013 29835 15071 29841
rect 15013 29801 15025 29835
rect 15059 29832 15071 29835
rect 15194 29832 15200 29844
rect 15059 29804 15200 29832
rect 15059 29801 15071 29804
rect 15013 29795 15071 29801
rect 15194 29792 15200 29804
rect 15252 29792 15258 29844
rect 18414 29792 18420 29844
rect 18472 29832 18478 29844
rect 18693 29835 18751 29841
rect 18693 29832 18705 29835
rect 18472 29804 18705 29832
rect 18472 29792 18478 29804
rect 18693 29801 18705 29804
rect 18739 29832 18751 29835
rect 20530 29832 20536 29844
rect 18739 29804 20536 29832
rect 18739 29801 18751 29804
rect 18693 29795 18751 29801
rect 20530 29792 20536 29804
rect 20588 29792 20594 29844
rect 20622 29792 20628 29844
rect 20680 29792 20686 29844
rect 21269 29835 21327 29841
rect 20824 29804 21220 29832
rect 12713 29767 12771 29773
rect 12713 29733 12725 29767
rect 12759 29764 12771 29767
rect 12759 29736 13768 29764
rect 12759 29733 12771 29736
rect 12713 29727 12771 29733
rect 13357 29699 13415 29705
rect 13357 29696 13369 29699
rect 12406 29668 13369 29696
rect 13357 29665 13369 29668
rect 13403 29696 13415 29699
rect 13633 29699 13691 29705
rect 13633 29696 13645 29699
rect 13403 29668 13645 29696
rect 13403 29665 13415 29668
rect 13357 29659 13415 29665
rect 13633 29665 13645 29668
rect 13679 29665 13691 29699
rect 13633 29659 13691 29665
rect 9582 29588 9588 29640
rect 9640 29628 9646 29640
rect 11348 29628 11376 29656
rect 9640 29600 11376 29628
rect 9640 29588 9646 29600
rect 13078 29588 13084 29640
rect 13136 29628 13142 29640
rect 13173 29631 13231 29637
rect 13173 29628 13185 29631
rect 13136 29600 13185 29628
rect 13136 29588 13142 29600
rect 13173 29597 13185 29600
rect 13219 29597 13231 29631
rect 13173 29591 13231 29597
rect 13265 29631 13323 29637
rect 13265 29597 13277 29631
rect 13311 29628 13323 29631
rect 13740 29628 13768 29736
rect 14274 29656 14280 29708
rect 14332 29696 14338 29708
rect 15197 29699 15255 29705
rect 15197 29696 15209 29699
rect 14332 29668 15209 29696
rect 14332 29656 14338 29668
rect 14090 29628 14096 29640
rect 13311 29600 14096 29628
rect 13311 29597 13323 29600
rect 13265 29591 13323 29597
rect 14090 29588 14096 29600
rect 14148 29588 14154 29640
rect 14642 29588 14648 29640
rect 14700 29588 14706 29640
rect 14844 29637 14872 29668
rect 15197 29665 15209 29668
rect 15243 29696 15255 29699
rect 15243 29668 15516 29696
rect 15243 29665 15255 29668
rect 15197 29659 15255 29665
rect 14829 29631 14887 29637
rect 14829 29597 14841 29631
rect 14875 29597 14887 29631
rect 14829 29591 14887 29597
rect 15102 29588 15108 29640
rect 15160 29628 15166 29640
rect 15381 29631 15439 29637
rect 15381 29628 15393 29631
rect 15160 29600 15393 29628
rect 15160 29588 15166 29600
rect 15381 29597 15393 29600
rect 15427 29597 15439 29631
rect 15488 29628 15516 29668
rect 16666 29656 16672 29708
rect 16724 29696 16730 29708
rect 16945 29699 17003 29705
rect 16945 29696 16957 29699
rect 16724 29668 16957 29696
rect 16724 29656 16730 29668
rect 16945 29665 16957 29668
rect 16991 29665 17003 29699
rect 16945 29659 17003 29665
rect 15488 29600 19196 29628
rect 15381 29591 15439 29597
rect 9852 29563 9910 29569
rect 9852 29529 9864 29563
rect 9898 29560 9910 29563
rect 10134 29560 10140 29572
rect 9898 29532 10140 29560
rect 9898 29529 9910 29532
rect 9852 29523 9910 29529
rect 10134 29520 10140 29532
rect 10192 29520 10198 29572
rect 11600 29563 11658 29569
rect 11600 29529 11612 29563
rect 11646 29560 11658 29563
rect 15648 29563 15706 29569
rect 11646 29532 12848 29560
rect 11646 29529 11658 29532
rect 11600 29523 11658 29529
rect 10502 29492 10508 29504
rect 9232 29464 10508 29492
rect 8159 29461 8171 29464
rect 8113 29455 8171 29461
rect 10502 29452 10508 29464
rect 10560 29452 10566 29504
rect 12820 29501 12848 29532
rect 15648 29529 15660 29563
rect 15694 29560 15706 29563
rect 15746 29560 15752 29572
rect 15694 29532 15752 29560
rect 15694 29529 15706 29532
rect 15648 29523 15706 29529
rect 15746 29520 15752 29532
rect 15804 29520 15810 29572
rect 17212 29563 17270 29569
rect 17212 29529 17224 29563
rect 17258 29560 17270 29563
rect 17402 29560 17408 29572
rect 17258 29532 17408 29560
rect 17258 29529 17270 29532
rect 17212 29523 17270 29529
rect 17402 29520 17408 29532
rect 17460 29520 17466 29572
rect 19168 29560 19196 29600
rect 19242 29588 19248 29640
rect 19300 29588 19306 29640
rect 19334 29588 19340 29640
rect 19392 29628 19398 29640
rect 19512 29631 19570 29637
rect 19512 29628 19524 29631
rect 19392 29600 19524 29628
rect 19392 29588 19398 29600
rect 19512 29597 19524 29600
rect 19558 29597 19570 29631
rect 20640 29628 20668 29792
rect 20717 29631 20775 29637
rect 20717 29628 20729 29631
rect 20640 29600 20729 29628
rect 19512 29591 19570 29597
rect 20717 29597 20729 29600
rect 20763 29597 20775 29631
rect 20717 29591 20775 29597
rect 20824 29560 20852 29804
rect 21082 29764 21088 29776
rect 21008 29736 21088 29764
rect 21008 29637 21036 29736
rect 21082 29724 21088 29736
rect 21140 29724 21146 29776
rect 21192 29764 21220 29804
rect 21269 29801 21281 29835
rect 21315 29832 21327 29835
rect 21358 29832 21364 29844
rect 21315 29804 21364 29832
rect 21315 29801 21327 29804
rect 21269 29795 21327 29801
rect 21358 29792 21364 29804
rect 21416 29792 21422 29844
rect 23658 29792 23664 29844
rect 23716 29792 23722 29844
rect 25038 29792 25044 29844
rect 25096 29832 25102 29844
rect 25777 29835 25835 29841
rect 25777 29832 25789 29835
rect 25096 29804 25789 29832
rect 25096 29792 25102 29804
rect 25777 29801 25789 29804
rect 25823 29832 25835 29835
rect 27062 29832 27068 29844
rect 25823 29804 27068 29832
rect 25823 29801 25835 29804
rect 25777 29795 25835 29801
rect 27062 29792 27068 29804
rect 27120 29792 27126 29844
rect 27154 29792 27160 29844
rect 27212 29792 27218 29844
rect 27338 29792 27344 29844
rect 27396 29832 27402 29844
rect 27433 29835 27491 29841
rect 27433 29832 27445 29835
rect 27396 29804 27445 29832
rect 27396 29792 27402 29804
rect 27433 29801 27445 29804
rect 27479 29801 27491 29835
rect 29549 29835 29607 29841
rect 29549 29832 29561 29835
rect 27433 29795 27491 29801
rect 28000 29804 29561 29832
rect 27172 29764 27200 29792
rect 28000 29764 28028 29804
rect 29549 29801 29561 29804
rect 29595 29801 29607 29835
rect 29549 29795 29607 29801
rect 29914 29792 29920 29844
rect 29972 29832 29978 29844
rect 30561 29835 30619 29841
rect 30561 29832 30573 29835
rect 29972 29804 30573 29832
rect 29972 29792 29978 29804
rect 30561 29801 30573 29804
rect 30607 29801 30619 29835
rect 30561 29795 30619 29801
rect 34146 29792 34152 29844
rect 34204 29832 34210 29844
rect 34517 29835 34575 29841
rect 34517 29832 34529 29835
rect 34204 29804 34529 29832
rect 34204 29792 34210 29804
rect 34517 29801 34529 29804
rect 34563 29801 34575 29835
rect 34517 29795 34575 29801
rect 21192 29736 24348 29764
rect 27172 29736 28028 29764
rect 21192 29696 21220 29736
rect 21361 29699 21419 29705
rect 21361 29696 21373 29699
rect 21192 29668 21373 29696
rect 20993 29631 21051 29637
rect 20993 29597 21005 29631
rect 21039 29597 21051 29631
rect 20993 29591 21051 29597
rect 21085 29631 21143 29637
rect 21085 29597 21097 29631
rect 21131 29628 21143 29631
rect 21192 29628 21220 29668
rect 21361 29665 21373 29668
rect 21407 29665 21419 29699
rect 21361 29659 21419 29665
rect 22002 29656 22008 29708
rect 22060 29696 22066 29708
rect 22557 29699 22615 29705
rect 22557 29696 22569 29699
rect 22060 29668 22569 29696
rect 22060 29656 22066 29668
rect 22557 29665 22569 29668
rect 22603 29665 22615 29699
rect 22557 29659 22615 29665
rect 21131 29600 21220 29628
rect 22465 29631 22523 29637
rect 21131 29597 21143 29600
rect 21085 29591 21143 29597
rect 22465 29597 22477 29631
rect 22511 29628 22523 29631
rect 23109 29631 23167 29637
rect 23109 29628 23121 29631
rect 22511 29600 23121 29628
rect 22511 29597 22523 29600
rect 22465 29591 22523 29597
rect 23109 29597 23121 29600
rect 23155 29628 23167 29631
rect 23198 29628 23204 29640
rect 23155 29600 23204 29628
rect 23155 29597 23167 29600
rect 23109 29591 23167 29597
rect 23198 29588 23204 29600
rect 23256 29588 23262 29640
rect 23477 29631 23535 29637
rect 23477 29597 23489 29631
rect 23523 29628 23535 29631
rect 23566 29628 23572 29640
rect 23523 29600 23572 29628
rect 23523 29597 23535 29600
rect 23477 29591 23535 29597
rect 23566 29588 23572 29600
rect 23624 29588 23630 29640
rect 24320 29628 24348 29736
rect 29362 29724 29368 29776
rect 29420 29764 29426 29776
rect 29420 29736 30144 29764
rect 29420 29724 29426 29736
rect 24394 29656 24400 29708
rect 24452 29656 24458 29708
rect 27246 29656 27252 29708
rect 27304 29696 27310 29708
rect 27985 29699 28043 29705
rect 27985 29696 27997 29699
rect 27304 29668 27997 29696
rect 27304 29656 27310 29668
rect 27985 29665 27997 29668
rect 28031 29665 28043 29699
rect 27985 29659 28043 29665
rect 25498 29628 25504 29640
rect 24320 29600 25504 29628
rect 25498 29588 25504 29600
rect 25556 29588 25562 29640
rect 26053 29631 26111 29637
rect 26053 29597 26065 29631
rect 26099 29628 26111 29631
rect 27264 29628 27292 29656
rect 26099 29600 27292 29628
rect 26099 29597 26111 29600
rect 26053 29591 26111 29597
rect 29546 29588 29552 29640
rect 29604 29628 29610 29640
rect 30116 29637 30144 29736
rect 33045 29699 33103 29705
rect 33045 29665 33057 29699
rect 33091 29696 33103 29699
rect 33594 29696 33600 29708
rect 33091 29668 33600 29696
rect 33091 29665 33103 29668
rect 33045 29659 33103 29665
rect 33594 29656 33600 29668
rect 33652 29656 33658 29708
rect 29733 29631 29791 29637
rect 29733 29628 29745 29631
rect 29604 29600 29745 29628
rect 29604 29588 29610 29600
rect 29733 29597 29745 29600
rect 29779 29628 29791 29631
rect 30101 29631 30159 29637
rect 29779 29600 30052 29628
rect 29779 29597 29791 29600
rect 29733 29591 29791 29597
rect 19168 29532 20852 29560
rect 20901 29563 20959 29569
rect 20901 29529 20913 29563
rect 20947 29560 20959 29563
rect 23293 29563 23351 29569
rect 23293 29560 23305 29563
rect 20947 29532 23305 29560
rect 20947 29529 20959 29532
rect 20901 29523 20959 29529
rect 23293 29529 23305 29532
rect 23339 29529 23351 29563
rect 23293 29523 23351 29529
rect 23385 29563 23443 29569
rect 23385 29529 23397 29563
rect 23431 29560 23443 29563
rect 23658 29560 23664 29572
rect 23431 29532 23664 29560
rect 23431 29529 23443 29532
rect 23385 29523 23443 29529
rect 12805 29495 12863 29501
rect 12805 29461 12817 29495
rect 12851 29461 12863 29495
rect 12805 29455 12863 29461
rect 15838 29452 15844 29504
rect 15896 29492 15902 29504
rect 16761 29495 16819 29501
rect 16761 29492 16773 29495
rect 15896 29464 16773 29492
rect 15896 29452 15902 29464
rect 16761 29461 16773 29464
rect 16807 29461 16819 29495
rect 16761 29455 16819 29461
rect 18322 29452 18328 29504
rect 18380 29452 18386 29504
rect 19886 29452 19892 29504
rect 19944 29492 19950 29504
rect 20916 29492 20944 29523
rect 23658 29520 23664 29532
rect 23716 29520 23722 29572
rect 24670 29569 24676 29572
rect 24664 29523 24676 29569
rect 24670 29520 24676 29523
rect 24728 29520 24734 29572
rect 26320 29563 26378 29569
rect 26320 29529 26332 29563
rect 26366 29560 26378 29563
rect 26970 29560 26976 29572
rect 26366 29532 26976 29560
rect 26366 29529 26378 29532
rect 26320 29523 26378 29529
rect 26970 29520 26976 29532
rect 27028 29520 27034 29572
rect 28252 29563 28310 29569
rect 28252 29529 28264 29563
rect 28298 29560 28310 29563
rect 28534 29560 28540 29572
rect 28298 29532 28540 29560
rect 28298 29529 28310 29532
rect 28252 29523 28310 29529
rect 28534 29520 28540 29532
rect 28592 29520 28598 29572
rect 29822 29520 29828 29572
rect 29880 29520 29886 29572
rect 29914 29520 29920 29572
rect 29972 29520 29978 29572
rect 30024 29560 30052 29600
rect 30101 29597 30113 29631
rect 30147 29597 30159 29631
rect 30101 29591 30159 29597
rect 32766 29588 32772 29640
rect 32824 29588 32830 29640
rect 30377 29563 30435 29569
rect 30377 29560 30389 29563
rect 30024 29532 30389 29560
rect 30377 29529 30389 29532
rect 30423 29529 30435 29563
rect 30377 29523 30435 29529
rect 33502 29520 33508 29572
rect 33560 29520 33566 29572
rect 19944 29464 20944 29492
rect 22005 29495 22063 29501
rect 19944 29452 19950 29464
rect 22005 29461 22017 29495
rect 22051 29492 22063 29495
rect 22094 29492 22100 29504
rect 22051 29464 22100 29492
rect 22051 29461 22063 29464
rect 22005 29455 22063 29461
rect 22094 29452 22100 29464
rect 22152 29452 22158 29504
rect 22370 29452 22376 29504
rect 22428 29452 22434 29504
rect 23014 29452 23020 29504
rect 23072 29492 23078 29504
rect 26418 29492 26424 29504
rect 23072 29464 26424 29492
rect 23072 29452 23078 29464
rect 26418 29452 26424 29464
rect 26476 29492 26482 29504
rect 27522 29492 27528 29504
rect 26476 29464 27528 29492
rect 26476 29452 26482 29464
rect 27522 29452 27528 29464
rect 27580 29452 27586 29504
rect 29086 29452 29092 29504
rect 29144 29492 29150 29504
rect 30193 29495 30251 29501
rect 30193 29492 30205 29495
rect 29144 29464 30205 29492
rect 29144 29452 29150 29464
rect 30193 29461 30205 29464
rect 30239 29461 30251 29495
rect 30193 29455 30251 29461
rect 1104 29402 35328 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35328 29402
rect 1104 29328 35328 29350
rect 3050 29248 3056 29300
rect 3108 29248 3114 29300
rect 3421 29291 3479 29297
rect 3421 29257 3433 29291
rect 3467 29288 3479 29291
rect 3602 29288 3608 29300
rect 3467 29260 3608 29288
rect 3467 29257 3479 29260
rect 3421 29251 3479 29257
rect 3602 29248 3608 29260
rect 3660 29248 3666 29300
rect 4246 29248 4252 29300
rect 4304 29248 4310 29300
rect 4614 29248 4620 29300
rect 4672 29248 4678 29300
rect 4706 29248 4712 29300
rect 4764 29248 4770 29300
rect 6730 29248 6736 29300
rect 6788 29248 6794 29300
rect 6822 29248 6828 29300
rect 6880 29248 6886 29300
rect 7374 29248 7380 29300
rect 7432 29248 7438 29300
rect 7742 29248 7748 29300
rect 7800 29248 7806 29300
rect 9674 29288 9680 29300
rect 7944 29260 9680 29288
rect 3513 29223 3571 29229
rect 3513 29189 3525 29223
rect 3559 29220 3571 29223
rect 4724 29220 4752 29248
rect 3559 29192 4752 29220
rect 5261 29223 5319 29229
rect 3559 29189 3571 29192
rect 3513 29183 3571 29189
rect 5261 29189 5273 29223
rect 5307 29220 5319 29223
rect 6362 29220 6368 29232
rect 5307 29192 6368 29220
rect 5307 29189 5319 29192
rect 5261 29183 5319 29189
rect 6362 29180 6368 29192
rect 6420 29180 6426 29232
rect 6840 29220 6868 29248
rect 7837 29223 7895 29229
rect 7837 29220 7849 29223
rect 6840 29192 7849 29220
rect 7837 29189 7849 29192
rect 7883 29189 7895 29223
rect 7837 29183 7895 29189
rect 5626 29152 5632 29164
rect 4908 29124 5632 29152
rect 3694 29044 3700 29096
rect 3752 29044 3758 29096
rect 4908 29093 4936 29124
rect 5626 29112 5632 29124
rect 5684 29152 5690 29164
rect 7944 29152 7972 29260
rect 9674 29248 9680 29260
rect 9732 29248 9738 29300
rect 9766 29248 9772 29300
rect 9824 29248 9830 29300
rect 10134 29248 10140 29300
rect 10192 29248 10198 29300
rect 10505 29291 10563 29297
rect 10505 29257 10517 29291
rect 10551 29288 10563 29291
rect 10594 29288 10600 29300
rect 10551 29260 10600 29288
rect 10551 29257 10563 29260
rect 10505 29251 10563 29257
rect 10594 29248 10600 29260
rect 10652 29248 10658 29300
rect 14461 29291 14519 29297
rect 14461 29257 14473 29291
rect 14507 29257 14519 29291
rect 14461 29251 14519 29257
rect 14921 29291 14979 29297
rect 14921 29257 14933 29291
rect 14967 29288 14979 29291
rect 15286 29288 15292 29300
rect 14967 29260 15292 29288
rect 14967 29257 14979 29260
rect 14921 29251 14979 29257
rect 8202 29180 8208 29232
rect 8260 29220 8266 29232
rect 9582 29220 9588 29232
rect 8260 29192 9588 29220
rect 8260 29180 8266 29192
rect 8404 29161 8432 29192
rect 9582 29180 9588 29192
rect 9640 29180 9646 29232
rect 13256 29223 13314 29229
rect 13256 29189 13268 29223
rect 13302 29220 13314 29223
rect 14476 29220 14504 29251
rect 15286 29248 15292 29260
rect 15344 29248 15350 29300
rect 15746 29248 15752 29300
rect 15804 29248 15810 29300
rect 15838 29248 15844 29300
rect 15896 29288 15902 29300
rect 16117 29291 16175 29297
rect 16117 29288 16129 29291
rect 15896 29260 16129 29288
rect 15896 29248 15902 29260
rect 16117 29257 16129 29260
rect 16163 29257 16175 29291
rect 16117 29251 16175 29257
rect 17402 29248 17408 29300
rect 17460 29248 17466 29300
rect 17773 29291 17831 29297
rect 17773 29257 17785 29291
rect 17819 29288 17831 29291
rect 18322 29288 18328 29300
rect 17819 29260 18328 29288
rect 17819 29257 17831 29260
rect 17773 29251 17831 29257
rect 18322 29248 18328 29260
rect 18380 29248 18386 29300
rect 19168 29260 22324 29288
rect 13302 29192 14504 29220
rect 15304 29220 15332 29248
rect 16209 29223 16267 29229
rect 16209 29220 16221 29223
rect 15304 29192 16221 29220
rect 13302 29189 13314 29192
rect 13256 29183 13314 29189
rect 16209 29189 16221 29192
rect 16255 29189 16267 29223
rect 16209 29183 16267 29189
rect 18233 29223 18291 29229
rect 18233 29189 18245 29223
rect 18279 29220 18291 29223
rect 19168 29220 19196 29260
rect 18279 29192 19196 29220
rect 18279 29189 18291 29192
rect 18233 29183 18291 29189
rect 5684 29124 7972 29152
rect 8389 29155 8447 29161
rect 5684 29112 5690 29124
rect 8389 29121 8401 29155
rect 8435 29121 8447 29155
rect 8389 29115 8447 29121
rect 8656 29155 8714 29161
rect 8656 29121 8668 29155
rect 8702 29152 8714 29155
rect 8938 29152 8944 29164
rect 8702 29124 8944 29152
rect 8702 29121 8714 29124
rect 8656 29115 8714 29121
rect 8938 29112 8944 29124
rect 8996 29112 9002 29164
rect 10597 29155 10655 29161
rect 10597 29121 10609 29155
rect 10643 29152 10655 29155
rect 11974 29152 11980 29164
rect 10643 29124 11980 29152
rect 10643 29121 10655 29124
rect 10597 29115 10655 29121
rect 11974 29112 11980 29124
rect 12032 29112 12038 29164
rect 14642 29152 14648 29164
rect 12406 29124 14320 29152
rect 4893 29087 4951 29093
rect 4893 29053 4905 29087
rect 4939 29053 4951 29087
rect 4893 29047 4951 29053
rect 5258 29044 5264 29096
rect 5316 29084 5322 29096
rect 5534 29084 5540 29096
rect 5316 29056 5540 29084
rect 5316 29044 5322 29056
rect 5534 29044 5540 29056
rect 5592 29084 5598 29096
rect 5997 29087 6055 29093
rect 5997 29084 6009 29087
rect 5592 29056 6009 29084
rect 5592 29044 5598 29056
rect 5997 29053 6009 29056
rect 6043 29053 6055 29087
rect 5997 29047 6055 29053
rect 6178 29044 6184 29096
rect 6236 29084 6242 29096
rect 6917 29087 6975 29093
rect 6917 29084 6929 29087
rect 6236 29056 6929 29084
rect 6236 29044 6242 29056
rect 6917 29053 6929 29056
rect 6963 29053 6975 29087
rect 6917 29047 6975 29053
rect 8021 29087 8079 29093
rect 8021 29053 8033 29087
rect 8067 29053 8079 29087
rect 8021 29047 8079 29053
rect 3786 28976 3792 29028
rect 3844 29016 3850 29028
rect 3973 29019 4031 29025
rect 3973 29016 3985 29019
rect 3844 28988 3985 29016
rect 3844 28976 3850 28988
rect 3973 28985 3985 28988
rect 4019 29016 4031 29019
rect 6196 29016 6224 29044
rect 4019 28988 6224 29016
rect 4019 28985 4031 28988
rect 3973 28979 4031 28985
rect 6270 28976 6276 29028
rect 6328 29016 6334 29028
rect 6365 29019 6423 29025
rect 6365 29016 6377 29019
rect 6328 28988 6377 29016
rect 6328 28976 6334 28988
rect 6365 28985 6377 28988
rect 6411 28985 6423 29019
rect 8036 29016 8064 29047
rect 10410 29044 10416 29096
rect 10468 29084 10474 29096
rect 10689 29087 10747 29093
rect 10689 29084 10701 29087
rect 10468 29056 10701 29084
rect 10468 29044 10474 29056
rect 10689 29053 10701 29056
rect 10735 29084 10747 29087
rect 10965 29087 11023 29093
rect 10965 29084 10977 29087
rect 10735 29056 10977 29084
rect 10735 29053 10747 29056
rect 10689 29047 10747 29053
rect 10965 29053 10977 29056
rect 11011 29053 11023 29087
rect 10965 29047 11023 29053
rect 8297 29019 8355 29025
rect 8297 29016 8309 29019
rect 8036 28988 8309 29016
rect 6365 28979 6423 28985
rect 8297 28985 8309 28988
rect 8343 29016 8355 29019
rect 12406 29016 12434 29124
rect 12986 29044 12992 29096
rect 13044 29044 13050 29096
rect 8343 28988 8432 29016
rect 8343 28985 8355 28988
rect 8297 28979 8355 28985
rect 8404 28948 8432 28988
rect 9324 28988 12434 29016
rect 8662 28948 8668 28960
rect 8404 28920 8668 28948
rect 8662 28908 8668 28920
rect 8720 28948 8726 28960
rect 9324 28948 9352 28988
rect 8720 28920 9352 28948
rect 14292 28948 14320 29124
rect 14384 29124 14648 29152
rect 14384 29025 14412 29124
rect 14642 29112 14648 29124
rect 14700 29152 14706 29164
rect 14829 29155 14887 29161
rect 14829 29152 14841 29155
rect 14700 29124 14841 29152
rect 14700 29112 14706 29124
rect 14829 29121 14841 29124
rect 14875 29121 14887 29155
rect 14829 29115 14887 29121
rect 15013 29087 15071 29093
rect 15013 29053 15025 29087
rect 15059 29084 15071 29087
rect 15289 29087 15347 29093
rect 15289 29084 15301 29087
rect 15059 29056 15301 29084
rect 15059 29053 15071 29056
rect 15013 29047 15071 29053
rect 15289 29053 15301 29056
rect 15335 29053 15347 29087
rect 15289 29047 15347 29053
rect 14369 29019 14427 29025
rect 14369 28985 14381 29019
rect 14415 28985 14427 29019
rect 15028 29016 15056 29047
rect 16022 29044 16028 29096
rect 16080 29084 16086 29096
rect 16301 29087 16359 29093
rect 16301 29084 16313 29087
rect 16080 29056 16313 29084
rect 16080 29044 16086 29056
rect 16301 29053 16313 29056
rect 16347 29084 16359 29087
rect 16669 29087 16727 29093
rect 16669 29084 16681 29087
rect 16347 29056 16681 29084
rect 16347 29053 16359 29056
rect 16301 29047 16359 29053
rect 16669 29053 16681 29056
rect 16715 29053 16727 29087
rect 16669 29047 16727 29053
rect 17865 29087 17923 29093
rect 17865 29053 17877 29087
rect 17911 29053 17923 29087
rect 17865 29047 17923 29053
rect 18049 29087 18107 29093
rect 18049 29053 18061 29087
rect 18095 29084 18107 29087
rect 18248 29084 18276 29183
rect 19242 29180 19248 29232
rect 19300 29220 19306 29232
rect 22094 29229 22100 29232
rect 19300 29192 21864 29220
rect 19300 29180 19306 29192
rect 19720 29161 19748 29192
rect 21836 29164 21864 29192
rect 22088 29183 22100 29229
rect 22094 29180 22100 29183
rect 22152 29180 22158 29232
rect 19705 29155 19763 29161
rect 19705 29121 19717 29155
rect 19751 29121 19763 29155
rect 19705 29115 19763 29121
rect 19972 29155 20030 29161
rect 19972 29121 19984 29155
rect 20018 29152 20030 29155
rect 20254 29152 20260 29164
rect 20018 29124 20260 29152
rect 20018 29121 20030 29124
rect 19972 29115 20030 29121
rect 20254 29112 20260 29124
rect 20312 29112 20318 29164
rect 21818 29112 21824 29164
rect 21876 29112 21882 29164
rect 22296 29152 22324 29260
rect 23198 29248 23204 29300
rect 23256 29248 23262 29300
rect 24670 29248 24676 29300
rect 24728 29248 24734 29300
rect 25038 29248 25044 29300
rect 25096 29248 25102 29300
rect 25133 29291 25191 29297
rect 25133 29257 25145 29291
rect 25179 29288 25191 29291
rect 25682 29288 25688 29300
rect 25179 29260 25688 29288
rect 25179 29257 25191 29260
rect 25133 29251 25191 29257
rect 22370 29180 22376 29232
rect 22428 29220 22434 29232
rect 23290 29220 23296 29232
rect 22428 29192 23296 29220
rect 22428 29180 22434 29192
rect 23290 29180 23296 29192
rect 23348 29220 23354 29232
rect 23753 29223 23811 29229
rect 23753 29220 23765 29223
rect 23348 29192 23765 29220
rect 23348 29180 23354 29192
rect 23753 29189 23765 29192
rect 23799 29220 23811 29223
rect 25148 29220 25176 29251
rect 25682 29248 25688 29260
rect 25740 29248 25746 29300
rect 26970 29248 26976 29300
rect 27028 29248 27034 29300
rect 27338 29248 27344 29300
rect 27396 29288 27402 29300
rect 27433 29291 27491 29297
rect 27433 29288 27445 29291
rect 27396 29260 27445 29288
rect 27396 29248 27402 29260
rect 27433 29257 27445 29260
rect 27479 29257 27491 29291
rect 27433 29251 27491 29257
rect 28534 29248 28540 29300
rect 28592 29248 28598 29300
rect 28905 29291 28963 29297
rect 28905 29257 28917 29291
rect 28951 29288 28963 29291
rect 29362 29288 29368 29300
rect 28951 29260 29368 29288
rect 28951 29257 28963 29260
rect 28905 29251 28963 29257
rect 29362 29248 29368 29260
rect 29420 29248 29426 29300
rect 29822 29248 29828 29300
rect 29880 29288 29886 29300
rect 30837 29291 30895 29297
rect 30837 29288 30849 29291
rect 29880 29260 30849 29288
rect 29880 29248 29886 29260
rect 30837 29257 30849 29260
rect 30883 29257 30895 29291
rect 30837 29251 30895 29257
rect 32766 29220 32772 29232
rect 23799 29192 25176 29220
rect 29472 29192 32772 29220
rect 23799 29189 23811 29192
rect 23753 29183 23811 29189
rect 22296 29124 22876 29152
rect 21634 29084 21640 29096
rect 18095 29056 18276 29084
rect 20732 29056 21640 29084
rect 18095 29053 18107 29056
rect 18049 29047 18107 29053
rect 14369 28979 14427 28985
rect 14476 28988 15056 29016
rect 17880 29016 17908 29047
rect 19702 29016 19708 29028
rect 17880 28988 19708 29016
rect 14476 28948 14504 28988
rect 19702 28976 19708 28988
rect 19760 28976 19766 29028
rect 20732 29016 20760 29056
rect 21634 29044 21640 29056
rect 21692 29044 21698 29096
rect 20640 28988 20760 29016
rect 14292 28920 14504 28948
rect 8720 28908 8726 28920
rect 19150 28908 19156 28960
rect 19208 28948 19214 28960
rect 20640 28948 20668 28988
rect 21082 28976 21088 29028
rect 21140 28976 21146 29028
rect 22848 29016 22876 29124
rect 23658 29112 23664 29164
rect 23716 29112 23722 29164
rect 27341 29155 27399 29161
rect 27341 29121 27353 29155
rect 27387 29152 27399 29155
rect 27430 29152 27436 29164
rect 27387 29124 27436 29152
rect 27387 29121 27399 29124
rect 27341 29115 27399 29121
rect 27430 29112 27436 29124
rect 27488 29152 27494 29164
rect 29472 29161 29500 29192
rect 32766 29180 32772 29192
rect 32824 29180 32830 29232
rect 29730 29161 29736 29164
rect 28997 29155 29055 29161
rect 28997 29152 29009 29155
rect 27488 29124 29009 29152
rect 27488 29112 27494 29124
rect 28997 29121 29009 29124
rect 29043 29121 29055 29155
rect 28997 29115 29055 29121
rect 29457 29155 29515 29161
rect 29457 29121 29469 29155
rect 29503 29121 29515 29155
rect 29457 29115 29515 29121
rect 29724 29115 29736 29161
rect 29730 29112 29736 29115
rect 29788 29112 29794 29164
rect 23474 29044 23480 29096
rect 23532 29084 23538 29096
rect 23845 29087 23903 29093
rect 23845 29084 23857 29087
rect 23532 29056 23857 29084
rect 23532 29044 23538 29056
rect 23845 29053 23857 29056
rect 23891 29053 23903 29087
rect 23845 29047 23903 29053
rect 24581 29087 24639 29093
rect 24581 29053 24593 29087
rect 24627 29084 24639 29087
rect 25317 29087 25375 29093
rect 25317 29084 25329 29087
rect 24627 29056 25329 29084
rect 24627 29053 24639 29056
rect 24581 29047 24639 29053
rect 25317 29053 25329 29056
rect 25363 29084 25375 29087
rect 25866 29084 25872 29096
rect 25363 29056 25872 29084
rect 25363 29053 25375 29056
rect 25317 29047 25375 29053
rect 24596 29016 24624 29047
rect 25866 29044 25872 29056
rect 25924 29044 25930 29096
rect 27522 29044 27528 29096
rect 27580 29084 27586 29096
rect 27801 29087 27859 29093
rect 27801 29084 27813 29087
rect 27580 29056 27813 29084
rect 27580 29044 27586 29056
rect 27801 29053 27813 29056
rect 27847 29053 27859 29087
rect 27801 29047 27859 29053
rect 29086 29044 29092 29096
rect 29144 29044 29150 29096
rect 22848 28988 24624 29016
rect 19208 28920 20668 28948
rect 19208 28908 19214 28920
rect 20714 28908 20720 28960
rect 20772 28948 20778 28960
rect 23014 28948 23020 28960
rect 20772 28920 23020 28948
rect 20772 28908 20778 28920
rect 23014 28908 23020 28920
rect 23072 28908 23078 28960
rect 23290 28908 23296 28960
rect 23348 28908 23354 28960
rect 1104 28858 35328 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 35328 28858
rect 1104 28784 35328 28806
rect 6362 28704 6368 28756
rect 6420 28704 6426 28756
rect 20254 28704 20260 28756
rect 20312 28704 20318 28756
rect 23474 28744 23480 28756
rect 22066 28716 23480 28744
rect 6178 28636 6184 28688
rect 6236 28676 6242 28688
rect 6457 28679 6515 28685
rect 6457 28676 6469 28679
rect 6236 28648 6469 28676
rect 6236 28636 6242 28648
rect 6457 28645 6469 28648
rect 6503 28645 6515 28679
rect 6457 28639 6515 28645
rect 20346 28636 20352 28688
rect 20404 28676 20410 28688
rect 20404 28648 20852 28676
rect 20404 28636 20410 28648
rect 19702 28568 19708 28620
rect 19760 28608 19766 28620
rect 20824 28617 20852 28648
rect 20717 28611 20775 28617
rect 20717 28608 20729 28611
rect 19760 28580 20729 28608
rect 19760 28568 19766 28580
rect 20717 28577 20729 28580
rect 20763 28577 20775 28611
rect 20717 28571 20775 28577
rect 20809 28611 20867 28617
rect 20809 28577 20821 28611
rect 20855 28608 20867 28611
rect 22066 28608 22094 28716
rect 23474 28704 23480 28716
rect 23532 28704 23538 28756
rect 23658 28704 23664 28756
rect 23716 28744 23722 28756
rect 24121 28747 24179 28753
rect 24121 28744 24133 28747
rect 23716 28716 24133 28744
rect 23716 28704 23722 28716
rect 24121 28713 24133 28716
rect 24167 28713 24179 28747
rect 24121 28707 24179 28713
rect 29730 28704 29736 28756
rect 29788 28704 29794 28756
rect 20855 28580 22094 28608
rect 20855 28577 20867 28580
rect 20809 28571 20867 28577
rect 27154 28568 27160 28620
rect 27212 28568 27218 28620
rect 29362 28568 29368 28620
rect 29420 28608 29426 28620
rect 30285 28611 30343 28617
rect 30285 28608 30297 28611
rect 29420 28580 30297 28608
rect 29420 28568 29426 28580
rect 30285 28577 30297 28580
rect 30331 28577 30343 28611
rect 30285 28571 30343 28577
rect 5534 28500 5540 28552
rect 5592 28500 5598 28552
rect 8202 28500 8208 28552
rect 8260 28540 8266 28552
rect 14369 28543 14427 28549
rect 14369 28540 14381 28543
rect 8260 28512 14381 28540
rect 8260 28500 8266 28512
rect 14369 28509 14381 28512
rect 14415 28509 14427 28543
rect 14369 28503 14427 28509
rect 14645 28543 14703 28549
rect 14645 28509 14657 28543
rect 14691 28540 14703 28543
rect 15010 28540 15016 28552
rect 14691 28512 15016 28540
rect 14691 28509 14703 28512
rect 14645 28503 14703 28509
rect 15010 28500 15016 28512
rect 15068 28540 15074 28552
rect 17405 28543 17463 28549
rect 17405 28540 17417 28543
rect 15068 28512 17417 28540
rect 15068 28500 15074 28512
rect 17405 28509 17417 28512
rect 17451 28509 17463 28543
rect 17405 28503 17463 28509
rect 20625 28543 20683 28549
rect 20625 28509 20637 28543
rect 20671 28540 20683 28543
rect 21082 28540 21088 28552
rect 20671 28512 21088 28540
rect 20671 28509 20683 28512
rect 20625 28503 20683 28509
rect 21082 28500 21088 28512
rect 21140 28500 21146 28552
rect 21818 28500 21824 28552
rect 21876 28540 21882 28552
rect 22278 28540 22284 28552
rect 21876 28512 22284 28540
rect 21876 28500 21882 28512
rect 22278 28500 22284 28512
rect 22336 28540 22342 28552
rect 22741 28543 22799 28549
rect 22741 28540 22753 28543
rect 22336 28512 22753 28540
rect 22336 28500 22342 28512
rect 22741 28509 22753 28512
rect 22787 28509 22799 28543
rect 22741 28503 22799 28509
rect 23008 28543 23066 28549
rect 23008 28509 23020 28543
rect 23054 28540 23066 28543
rect 23290 28540 23296 28552
rect 23054 28512 23296 28540
rect 23054 28509 23066 28512
rect 23008 28503 23066 28509
rect 23290 28500 23296 28512
rect 23348 28500 23354 28552
rect 23382 28500 23388 28552
rect 23440 28540 23446 28552
rect 23440 28512 29684 28540
rect 23440 28500 23446 28512
rect 27424 28475 27482 28481
rect 27424 28441 27436 28475
rect 27470 28472 27482 28475
rect 27614 28472 27620 28484
rect 27470 28444 27620 28472
rect 27470 28441 27482 28444
rect 27424 28435 27482 28441
rect 27614 28432 27620 28444
rect 27672 28432 27678 28484
rect 28166 28472 28172 28484
rect 27908 28444 28172 28472
rect 3418 28364 3424 28416
rect 3476 28364 3482 28416
rect 5258 28364 5264 28416
rect 5316 28404 5322 28416
rect 10226 28404 10232 28416
rect 5316 28376 10232 28404
rect 5316 28364 5322 28376
rect 10226 28364 10232 28376
rect 10284 28364 10290 28416
rect 17218 28364 17224 28416
rect 17276 28364 17282 28416
rect 22738 28364 22744 28416
rect 22796 28404 22802 28416
rect 27908 28404 27936 28444
rect 28166 28432 28172 28444
rect 28224 28432 28230 28484
rect 29656 28481 29684 28512
rect 29822 28500 29828 28552
rect 29880 28540 29886 28552
rect 30101 28543 30159 28549
rect 30101 28540 30113 28543
rect 29880 28512 30113 28540
rect 29880 28500 29886 28512
rect 30101 28509 30113 28512
rect 30147 28509 30159 28543
rect 30101 28503 30159 28509
rect 29641 28475 29699 28481
rect 29641 28441 29653 28475
rect 29687 28472 29699 28475
rect 30193 28475 30251 28481
rect 30193 28472 30205 28475
rect 29687 28444 30205 28472
rect 29687 28441 29699 28444
rect 29641 28435 29699 28441
rect 30193 28441 30205 28444
rect 30239 28441 30251 28475
rect 30193 28435 30251 28441
rect 22796 28376 27936 28404
rect 22796 28364 22802 28376
rect 27982 28364 27988 28416
rect 28040 28404 28046 28416
rect 28537 28407 28595 28413
rect 28537 28404 28549 28407
rect 28040 28376 28549 28404
rect 28040 28364 28046 28376
rect 28537 28373 28549 28376
rect 28583 28373 28595 28407
rect 28537 28367 28595 28373
rect 29362 28364 29368 28416
rect 29420 28364 29426 28416
rect 1104 28314 35328 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35328 28314
rect 1104 28240 35328 28262
rect 1581 28203 1639 28209
rect 1581 28169 1593 28203
rect 1627 28200 1639 28203
rect 7929 28203 7987 28209
rect 7929 28200 7941 28203
rect 1627 28172 6040 28200
rect 1627 28169 1639 28172
rect 1581 28163 1639 28169
rect 2866 28092 2872 28144
rect 2924 28132 2930 28144
rect 3053 28135 3111 28141
rect 3053 28132 3065 28135
rect 2924 28104 3065 28132
rect 2924 28092 2930 28104
rect 3053 28101 3065 28104
rect 3099 28101 3111 28135
rect 3053 28095 3111 28101
rect 4525 28135 4583 28141
rect 4525 28101 4537 28135
rect 4571 28132 4583 28135
rect 4706 28132 4712 28144
rect 4571 28104 4712 28132
rect 4571 28101 4583 28104
rect 4525 28095 4583 28101
rect 4706 28092 4712 28104
rect 4764 28092 4770 28144
rect 4985 28135 5043 28141
rect 4985 28101 4997 28135
rect 5031 28132 5043 28135
rect 5258 28132 5264 28144
rect 5031 28104 5264 28132
rect 5031 28101 5043 28104
rect 4985 28095 5043 28101
rect 1302 28024 1308 28076
rect 1360 28064 1366 28076
rect 1397 28067 1455 28073
rect 1397 28064 1409 28067
rect 1360 28036 1409 28064
rect 1360 28024 1366 28036
rect 1397 28033 1409 28036
rect 1443 28064 1455 28067
rect 1673 28067 1731 28073
rect 1673 28064 1685 28067
rect 1443 28036 1685 28064
rect 1443 28033 1455 28036
rect 1397 28027 1455 28033
rect 1673 28033 1685 28036
rect 1719 28033 1731 28067
rect 1673 28027 1731 28033
rect 2777 28067 2835 28073
rect 2777 28033 2789 28067
rect 2823 28064 2835 28067
rect 3237 28067 3295 28073
rect 3237 28064 3249 28067
rect 2823 28036 3249 28064
rect 2823 28033 2835 28036
rect 2777 28027 2835 28033
rect 3237 28033 3249 28036
rect 3283 28064 3295 28067
rect 3418 28064 3424 28076
rect 3283 28036 3424 28064
rect 3283 28033 3295 28036
rect 3237 28027 3295 28033
rect 3418 28024 3424 28036
rect 3476 28064 3482 28076
rect 4154 28064 4160 28076
rect 3476 28036 4160 28064
rect 3476 28024 3482 28036
rect 4154 28024 4160 28036
rect 4212 28024 4218 28076
rect 4246 28024 4252 28076
rect 4304 28024 4310 28076
rect 4433 28067 4491 28073
rect 4433 28033 4445 28067
rect 4479 28033 4491 28067
rect 4433 28027 4491 28033
rect 4617 28067 4675 28073
rect 4617 28033 4629 28067
rect 4663 28064 4675 28067
rect 4890 28064 4896 28076
rect 4663 28036 4896 28064
rect 4663 28033 4675 28036
rect 4617 28027 4675 28033
rect 3786 27956 3792 28008
rect 3844 27996 3850 28008
rect 3881 27999 3939 28005
rect 3881 27996 3893 27999
rect 3844 27968 3893 27996
rect 3844 27956 3850 27968
rect 3881 27965 3893 27968
rect 3927 27965 3939 27999
rect 4448 27996 4476 28027
rect 4890 28024 4896 28036
rect 4948 28064 4954 28076
rect 5000 28064 5028 28095
rect 5258 28092 5264 28104
rect 5316 28092 5322 28144
rect 6012 28073 6040 28172
rect 7392 28172 7941 28200
rect 7392 28141 7420 28172
rect 7929 28169 7941 28172
rect 7975 28200 7987 28203
rect 10042 28200 10048 28212
rect 7975 28172 10048 28200
rect 7975 28169 7987 28172
rect 7929 28163 7987 28169
rect 10042 28160 10048 28172
rect 10100 28160 10106 28212
rect 14182 28160 14188 28212
rect 14240 28200 14246 28212
rect 16025 28203 16083 28209
rect 16025 28200 16037 28203
rect 14240 28172 14412 28200
rect 14240 28160 14246 28172
rect 14384 28141 14412 28172
rect 15672 28172 16037 28200
rect 7377 28135 7435 28141
rect 7377 28101 7389 28135
rect 7423 28101 7435 28135
rect 7377 28095 7435 28101
rect 14369 28135 14427 28141
rect 14369 28101 14381 28135
rect 14415 28101 14427 28135
rect 14369 28095 14427 28101
rect 15470 28092 15476 28144
rect 15528 28132 15534 28144
rect 15672 28141 15700 28172
rect 16025 28169 16037 28172
rect 16071 28200 16083 28203
rect 16206 28200 16212 28212
rect 16071 28172 16212 28200
rect 16071 28169 16083 28172
rect 16025 28163 16083 28169
rect 16206 28160 16212 28172
rect 16264 28160 16270 28212
rect 23106 28200 23112 28212
rect 22756 28172 23112 28200
rect 22756 28141 22784 28172
rect 23106 28160 23112 28172
rect 23164 28200 23170 28212
rect 24762 28200 24768 28212
rect 23164 28172 24768 28200
rect 23164 28160 23170 28172
rect 24762 28160 24768 28172
rect 24820 28160 24826 28212
rect 26789 28203 26847 28209
rect 26789 28169 26801 28203
rect 26835 28200 26847 28203
rect 26878 28200 26884 28212
rect 26835 28172 26884 28200
rect 26835 28169 26847 28172
rect 26789 28163 26847 28169
rect 26878 28160 26884 28172
rect 26936 28200 26942 28212
rect 27062 28200 27068 28212
rect 26936 28172 27068 28200
rect 26936 28160 26942 28172
rect 27062 28160 27068 28172
rect 27120 28200 27126 28212
rect 27120 28172 27200 28200
rect 27120 28160 27126 28172
rect 27172 28141 27200 28172
rect 27614 28160 27620 28212
rect 27672 28160 27678 28212
rect 27982 28160 27988 28212
rect 28040 28160 28046 28212
rect 15657 28135 15715 28141
rect 15657 28132 15669 28135
rect 15528 28104 15669 28132
rect 15528 28092 15534 28104
rect 15657 28101 15669 28104
rect 15703 28101 15715 28135
rect 15657 28095 15715 28101
rect 15841 28135 15899 28141
rect 15841 28101 15853 28135
rect 15887 28132 15899 28135
rect 16301 28135 16359 28141
rect 16301 28132 16313 28135
rect 15887 28104 16313 28132
rect 15887 28101 15899 28104
rect 15841 28095 15899 28101
rect 16301 28101 16313 28104
rect 16347 28132 16359 28135
rect 22741 28135 22799 28141
rect 16347 28104 20760 28132
rect 16347 28101 16359 28104
rect 16301 28095 16359 28101
rect 4948 28036 5028 28064
rect 5997 28067 6055 28073
rect 4948 28024 4954 28036
rect 5997 28033 6009 28067
rect 6043 28033 6055 28067
rect 5997 28027 6055 28033
rect 6086 28024 6092 28076
rect 6144 28064 6150 28076
rect 6733 28067 6791 28073
rect 6733 28064 6745 28067
rect 6144 28036 6745 28064
rect 6144 28024 6150 28036
rect 6733 28033 6745 28036
rect 6779 28064 6791 28067
rect 7193 28067 7251 28073
rect 7193 28064 7205 28067
rect 6779 28036 7205 28064
rect 6779 28033 6791 28036
rect 6733 28027 6791 28033
rect 7193 28033 7205 28036
rect 7239 28033 7251 28067
rect 7193 28027 7251 28033
rect 7466 28024 7472 28076
rect 7524 28024 7530 28076
rect 7558 28024 7564 28076
rect 7616 28024 7622 28076
rect 12158 28024 12164 28076
rect 12216 28064 12222 28076
rect 12630 28067 12688 28073
rect 12630 28064 12642 28067
rect 12216 28036 12642 28064
rect 12216 28024 12222 28036
rect 12630 28033 12642 28036
rect 12676 28033 12688 28067
rect 12630 28027 12688 28033
rect 16666 28024 16672 28076
rect 16724 28024 16730 28076
rect 16758 28024 16764 28076
rect 16816 28064 16822 28076
rect 16925 28067 16983 28073
rect 16925 28064 16937 28067
rect 16816 28036 16937 28064
rect 16816 28024 16822 28036
rect 16925 28033 16937 28036
rect 16971 28033 16983 28067
rect 16925 28027 16983 28033
rect 20070 28024 20076 28076
rect 20128 28024 20134 28076
rect 4798 27996 4804 28008
rect 4448 27968 4804 27996
rect 3881 27959 3939 27965
rect 4798 27956 4804 27968
rect 4856 27996 4862 28008
rect 6825 27999 6883 28005
rect 4856 27968 5212 27996
rect 4856 27956 4862 27968
rect 4798 27820 4804 27872
rect 4856 27820 4862 27872
rect 5184 27869 5212 27968
rect 6825 27965 6837 27999
rect 6871 27965 6883 27999
rect 6825 27959 6883 27965
rect 7009 27999 7067 28005
rect 7009 27965 7021 27999
rect 7055 27996 7067 27999
rect 8113 27999 8171 28005
rect 8113 27996 8125 27999
rect 7055 27968 8125 27996
rect 7055 27965 7067 27968
rect 7009 27959 7067 27965
rect 8113 27965 8125 27968
rect 8159 27996 8171 27999
rect 9950 27996 9956 28008
rect 8159 27968 9956 27996
rect 8159 27965 8171 27968
rect 8113 27959 8171 27965
rect 6181 27931 6239 27937
rect 6181 27897 6193 27931
rect 6227 27928 6239 27931
rect 6840 27928 6868 27959
rect 9950 27956 9956 27968
rect 10008 27956 10014 28008
rect 12897 27999 12955 28005
rect 12897 27965 12909 27999
rect 12943 27996 12955 27999
rect 12986 27996 12992 28008
rect 12943 27968 12992 27996
rect 12943 27965 12955 27968
rect 12897 27959 12955 27965
rect 12986 27956 12992 27968
rect 13044 27996 13050 28008
rect 14550 27996 14556 28008
rect 13044 27968 14556 27996
rect 13044 27956 13050 27968
rect 14550 27956 14556 27968
rect 14608 27996 14614 28008
rect 15102 27996 15108 28008
rect 14608 27968 15108 27996
rect 14608 27956 14614 27968
rect 15102 27956 15108 27968
rect 15160 27956 15166 28008
rect 20162 27956 20168 28008
rect 20220 27956 20226 28008
rect 20349 27999 20407 28005
rect 20349 27965 20361 27999
rect 20395 27996 20407 27999
rect 20438 27996 20444 28008
rect 20395 27968 20444 27996
rect 20395 27965 20407 27968
rect 20349 27959 20407 27965
rect 20438 27956 20444 27968
rect 20496 27996 20502 28008
rect 20496 27968 20668 27996
rect 20496 27956 20502 27968
rect 7190 27928 7196 27940
rect 6227 27900 7196 27928
rect 6227 27897 6239 27900
rect 6181 27891 6239 27897
rect 7190 27888 7196 27900
rect 7248 27888 7254 27940
rect 7745 27931 7803 27937
rect 7745 27897 7757 27931
rect 7791 27928 7803 27931
rect 9030 27928 9036 27940
rect 7791 27900 9036 27928
rect 7791 27897 7803 27900
rect 7745 27891 7803 27897
rect 9030 27888 9036 27900
rect 9088 27888 9094 27940
rect 20640 27872 20668 27968
rect 20732 27928 20760 28104
rect 22741 28101 22753 28135
rect 22787 28101 22799 28135
rect 22741 28095 22799 28101
rect 27157 28135 27215 28141
rect 27157 28101 27169 28135
rect 27203 28101 27215 28135
rect 27157 28095 27215 28101
rect 27249 28135 27307 28141
rect 27249 28101 27261 28135
rect 27295 28132 27307 28135
rect 28000 28132 28028 28160
rect 27295 28104 28028 28132
rect 27295 28101 27307 28104
rect 27249 28095 27307 28101
rect 21637 28067 21695 28073
rect 21637 28033 21649 28067
rect 21683 28064 21695 28067
rect 22646 28064 22652 28076
rect 21683 28036 22652 28064
rect 21683 28033 21695 28036
rect 21637 28027 21695 28033
rect 22646 28024 22652 28036
rect 22704 28024 22710 28076
rect 25308 28067 25366 28073
rect 25308 28033 25320 28067
rect 25354 28064 25366 28067
rect 25590 28064 25596 28076
rect 25354 28036 25596 28064
rect 25354 28033 25366 28036
rect 25308 28027 25366 28033
rect 25590 28024 25596 28036
rect 25648 28024 25654 28076
rect 26418 28024 26424 28076
rect 26476 28064 26482 28076
rect 26973 28067 27031 28073
rect 26973 28064 26985 28067
rect 26476 28036 26985 28064
rect 26476 28024 26482 28036
rect 26973 28033 26985 28036
rect 27019 28033 27031 28067
rect 26973 28027 27031 28033
rect 27341 28067 27399 28073
rect 27341 28033 27353 28067
rect 27387 28064 27399 28067
rect 28994 28064 29000 28076
rect 27387 28036 29000 28064
rect 27387 28033 27399 28036
rect 27341 28027 27399 28033
rect 28994 28024 29000 28036
rect 29052 28024 29058 28076
rect 34514 28024 34520 28076
rect 34572 28024 34578 28076
rect 22005 27999 22063 28005
rect 22005 27965 22017 27999
rect 22051 27996 22063 27999
rect 22278 27996 22284 28008
rect 22051 27968 22284 27996
rect 22051 27965 22063 27968
rect 22005 27959 22063 27965
rect 22278 27956 22284 27968
rect 22336 27956 22342 28008
rect 24118 27956 24124 28008
rect 24176 27996 24182 28008
rect 25041 27999 25099 28005
rect 25041 27996 25053 27999
rect 24176 27968 25053 27996
rect 24176 27956 24182 27968
rect 25041 27965 25053 27968
rect 25087 27965 25099 27999
rect 28077 27999 28135 28005
rect 28077 27996 28089 27999
rect 25041 27959 25099 27965
rect 26528 27968 28089 27996
rect 23290 27928 23296 27940
rect 20732 27900 23296 27928
rect 23290 27888 23296 27900
rect 23348 27928 23354 27940
rect 23842 27928 23848 27940
rect 23348 27900 23848 27928
rect 23348 27888 23354 27900
rect 23842 27888 23848 27900
rect 23900 27888 23906 27940
rect 26528 27872 26556 27968
rect 28077 27965 28089 27968
rect 28123 27965 28135 27999
rect 28077 27959 28135 27965
rect 28092 27928 28120 27959
rect 28166 27956 28172 28008
rect 28224 27996 28230 28008
rect 28445 27999 28503 28005
rect 28445 27996 28457 27999
rect 28224 27968 28457 27996
rect 28224 27956 28230 27968
rect 28445 27965 28457 27968
rect 28491 27965 28503 27999
rect 28445 27959 28503 27965
rect 34793 27999 34851 28005
rect 34793 27965 34805 27999
rect 34839 27996 34851 27999
rect 35342 27996 35348 28008
rect 34839 27968 35348 27996
rect 34839 27965 34851 27968
rect 34793 27959 34851 27965
rect 35342 27956 35348 27968
rect 35400 27956 35406 28008
rect 29365 27931 29423 27937
rect 29365 27928 29377 27931
rect 28092 27900 29377 27928
rect 29365 27897 29377 27900
rect 29411 27928 29423 27931
rect 29914 27928 29920 27940
rect 29411 27900 29920 27928
rect 29411 27897 29423 27900
rect 29365 27891 29423 27897
rect 29914 27888 29920 27900
rect 29972 27888 29978 27940
rect 5169 27863 5227 27869
rect 5169 27829 5181 27863
rect 5215 27860 5227 27863
rect 5350 27860 5356 27872
rect 5215 27832 5356 27860
rect 5215 27829 5227 27832
rect 5169 27823 5227 27829
rect 5350 27820 5356 27832
rect 5408 27820 5414 27872
rect 6270 27820 6276 27872
rect 6328 27860 6334 27872
rect 6365 27863 6423 27869
rect 6365 27860 6377 27863
rect 6328 27832 6377 27860
rect 6328 27820 6334 27832
rect 6365 27829 6377 27832
rect 6411 27829 6423 27863
rect 6365 27823 6423 27829
rect 8294 27820 8300 27872
rect 8352 27860 8358 27872
rect 8846 27860 8852 27872
rect 8352 27832 8852 27860
rect 8352 27820 8358 27832
rect 8846 27820 8852 27832
rect 8904 27820 8910 27872
rect 11517 27863 11575 27869
rect 11517 27829 11529 27863
rect 11563 27860 11575 27863
rect 11790 27860 11796 27872
rect 11563 27832 11796 27860
rect 11563 27829 11575 27832
rect 11517 27823 11575 27829
rect 11790 27820 11796 27832
rect 11848 27820 11854 27872
rect 12526 27820 12532 27872
rect 12584 27860 12590 27872
rect 13078 27860 13084 27872
rect 12584 27832 13084 27860
rect 12584 27820 12590 27832
rect 13078 27820 13084 27832
rect 13136 27820 13142 27872
rect 18046 27820 18052 27872
rect 18104 27820 18110 27872
rect 18138 27820 18144 27872
rect 18196 27820 18202 27872
rect 19702 27820 19708 27872
rect 19760 27820 19766 27872
rect 20622 27820 20628 27872
rect 20680 27820 20686 27872
rect 21453 27863 21511 27869
rect 21453 27829 21465 27863
rect 21499 27860 21511 27863
rect 21634 27860 21640 27872
rect 21499 27832 21640 27860
rect 21499 27829 21511 27832
rect 21453 27823 21511 27829
rect 21634 27820 21640 27832
rect 21692 27820 21698 27872
rect 22094 27820 22100 27872
rect 22152 27860 22158 27872
rect 22833 27863 22891 27869
rect 22833 27860 22845 27863
rect 22152 27832 22845 27860
rect 22152 27820 22158 27832
rect 22833 27829 22845 27832
rect 22879 27829 22891 27863
rect 22833 27823 22891 27829
rect 26418 27820 26424 27872
rect 26476 27820 26482 27872
rect 26510 27820 26516 27872
rect 26568 27820 26574 27872
rect 27430 27820 27436 27872
rect 27488 27860 27494 27872
rect 27525 27863 27583 27869
rect 27525 27860 27537 27863
rect 27488 27832 27537 27860
rect 27488 27820 27494 27832
rect 27525 27829 27537 27832
rect 27571 27829 27583 27863
rect 27525 27823 27583 27829
rect 28721 27863 28779 27869
rect 28721 27829 28733 27863
rect 28767 27860 28779 27863
rect 28994 27860 29000 27872
rect 28767 27832 29000 27860
rect 28767 27829 28779 27832
rect 28721 27823 28779 27829
rect 28994 27820 29000 27832
rect 29052 27820 29058 27872
rect 1104 27770 35328 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 35328 27770
rect 1104 27696 35328 27718
rect 6086 27616 6092 27668
rect 6144 27616 6150 27668
rect 7466 27616 7472 27668
rect 7524 27656 7530 27668
rect 7561 27659 7619 27665
rect 7561 27656 7573 27659
rect 7524 27628 7573 27656
rect 7524 27616 7530 27628
rect 7561 27625 7573 27628
rect 7607 27625 7619 27659
rect 7561 27619 7619 27625
rect 9493 27659 9551 27665
rect 9493 27625 9505 27659
rect 9539 27656 9551 27659
rect 15838 27656 15844 27668
rect 9539 27628 15844 27656
rect 9539 27625 9551 27628
rect 9493 27619 9551 27625
rect 15838 27616 15844 27628
rect 15896 27616 15902 27668
rect 16758 27616 16764 27668
rect 16816 27616 16822 27668
rect 18138 27656 18144 27668
rect 18064 27628 18144 27656
rect 3605 27591 3663 27597
rect 3605 27557 3617 27591
rect 3651 27588 3663 27591
rect 4062 27588 4068 27600
rect 3651 27560 4068 27588
rect 3651 27557 3663 27560
rect 3605 27551 3663 27557
rect 4062 27548 4068 27560
rect 4120 27548 4126 27600
rect 12158 27548 12164 27600
rect 12216 27548 12222 27600
rect 12621 27591 12679 27597
rect 12621 27557 12633 27591
rect 12667 27588 12679 27591
rect 13538 27588 13544 27600
rect 12667 27560 13544 27588
rect 12667 27557 12679 27560
rect 12621 27551 12679 27557
rect 2222 27480 2228 27532
rect 2280 27480 2286 27532
rect 4246 27480 4252 27532
rect 4304 27520 4310 27532
rect 4433 27523 4491 27529
rect 4433 27520 4445 27523
rect 4304 27492 4445 27520
rect 4304 27480 4310 27492
rect 4433 27489 4445 27492
rect 4479 27489 4491 27523
rect 4433 27483 4491 27489
rect 7190 27480 7196 27532
rect 7248 27520 7254 27532
rect 8202 27520 8208 27532
rect 7248 27492 8208 27520
rect 7248 27480 7254 27492
rect 8202 27480 8208 27492
rect 8260 27520 8266 27532
rect 8481 27523 8539 27529
rect 8481 27520 8493 27523
rect 8260 27492 8493 27520
rect 8260 27480 8266 27492
rect 8481 27489 8493 27492
rect 8527 27489 8539 27523
rect 8481 27483 8539 27489
rect 8573 27523 8631 27529
rect 8573 27489 8585 27523
rect 8619 27489 8631 27523
rect 9122 27520 9128 27532
rect 8573 27483 8631 27489
rect 8956 27492 9128 27520
rect 2240 27452 2268 27480
rect 4709 27455 4767 27461
rect 4709 27452 4721 27455
rect 2240 27424 4721 27452
rect 4709 27421 4721 27424
rect 4755 27452 4767 27455
rect 6178 27452 6184 27464
rect 4755 27424 6184 27452
rect 4755 27421 4767 27424
rect 4709 27415 4767 27421
rect 6178 27412 6184 27424
rect 6236 27412 6242 27464
rect 8294 27412 8300 27464
rect 8352 27452 8358 27464
rect 8588 27452 8616 27483
rect 8956 27461 8984 27492
rect 9122 27480 9128 27492
rect 9180 27480 9186 27532
rect 10686 27480 10692 27532
rect 10744 27520 10750 27532
rect 11609 27523 11667 27529
rect 11609 27520 11621 27523
rect 10744 27492 11621 27520
rect 10744 27480 10750 27492
rect 11609 27489 11621 27492
rect 11655 27520 11667 27523
rect 11655 27492 11928 27520
rect 11655 27489 11667 27492
rect 11609 27483 11667 27489
rect 8352 27424 8616 27452
rect 8941 27455 8999 27461
rect 8352 27412 8358 27424
rect 8941 27421 8953 27455
rect 8987 27421 8999 27455
rect 8941 27415 8999 27421
rect 9030 27412 9036 27464
rect 9088 27412 9094 27464
rect 9214 27452 9220 27464
rect 9140 27424 9220 27452
rect 2492 27387 2550 27393
rect 2492 27353 2504 27387
rect 2538 27384 2550 27387
rect 2590 27384 2596 27396
rect 2538 27356 2596 27384
rect 2538 27353 2550 27356
rect 2492 27347 2550 27353
rect 2590 27344 2596 27356
rect 2648 27344 2654 27396
rect 3050 27344 3056 27396
rect 3108 27384 3114 27396
rect 4249 27387 4307 27393
rect 4249 27384 4261 27387
rect 3108 27356 4261 27384
rect 3108 27344 3114 27356
rect 4249 27353 4261 27356
rect 4295 27353 4307 27387
rect 4249 27347 4307 27353
rect 4976 27387 5034 27393
rect 4976 27353 4988 27387
rect 5022 27384 5034 27387
rect 6270 27384 6276 27396
rect 5022 27356 6276 27384
rect 5022 27353 5034 27356
rect 4976 27347 5034 27353
rect 6270 27344 6276 27356
rect 6328 27344 6334 27396
rect 6448 27387 6506 27393
rect 6448 27353 6460 27387
rect 6494 27384 6506 27387
rect 6822 27384 6828 27396
rect 6494 27356 6828 27384
rect 6494 27353 6506 27356
rect 6448 27347 6506 27353
rect 6822 27344 6828 27356
rect 6880 27344 6886 27396
rect 8389 27387 8447 27393
rect 8389 27353 8401 27387
rect 8435 27384 8447 27387
rect 9140 27384 9168 27424
rect 9214 27412 9220 27424
rect 9272 27412 9278 27464
rect 9309 27455 9367 27461
rect 9309 27421 9321 27455
rect 9355 27421 9367 27455
rect 9309 27415 9367 27421
rect 8435 27356 9168 27384
rect 9324 27384 9352 27415
rect 9582 27412 9588 27464
rect 9640 27412 9646 27464
rect 11790 27412 11796 27464
rect 11848 27412 11854 27464
rect 11900 27452 11928 27492
rect 11974 27480 11980 27532
rect 12032 27520 12038 27532
rect 12636 27520 12664 27551
rect 13538 27548 13544 27560
rect 13596 27548 13602 27600
rect 15654 27548 15660 27600
rect 15712 27588 15718 27600
rect 17954 27588 17960 27600
rect 15712 27560 17960 27588
rect 15712 27548 15718 27560
rect 17954 27548 17960 27560
rect 18012 27548 18018 27600
rect 12032 27492 12664 27520
rect 12805 27523 12863 27529
rect 12032 27480 12038 27492
rect 12805 27489 12817 27523
rect 12851 27520 12863 27523
rect 13357 27523 13415 27529
rect 13357 27520 13369 27523
rect 12851 27492 13369 27520
rect 12851 27489 12863 27492
rect 12805 27483 12863 27489
rect 13357 27489 13369 27492
rect 13403 27520 13415 27523
rect 14090 27520 14096 27532
rect 13403 27492 14096 27520
rect 13403 27489 13415 27492
rect 13357 27483 13415 27489
rect 12820 27452 12848 27483
rect 14090 27480 14096 27492
rect 14148 27480 14154 27532
rect 16942 27480 16948 27532
rect 17000 27520 17006 27532
rect 17313 27523 17371 27529
rect 17313 27520 17325 27523
rect 17000 27492 17325 27520
rect 17000 27480 17006 27492
rect 17313 27489 17325 27492
rect 17359 27520 17371 27523
rect 18064 27520 18092 27628
rect 18138 27616 18144 27628
rect 18196 27616 18202 27668
rect 20162 27616 20168 27668
rect 20220 27656 20226 27668
rect 20530 27656 20536 27668
rect 20220 27628 20536 27656
rect 20220 27616 20226 27628
rect 20530 27616 20536 27628
rect 20588 27656 20594 27668
rect 20625 27659 20683 27665
rect 20625 27656 20637 27659
rect 20588 27628 20637 27656
rect 20588 27616 20594 27628
rect 20625 27625 20637 27628
rect 20671 27625 20683 27659
rect 20625 27619 20683 27625
rect 20898 27616 20904 27668
rect 20956 27656 20962 27668
rect 22281 27659 22339 27665
rect 20956 27628 22232 27656
rect 20956 27616 20962 27628
rect 22204 27588 22232 27628
rect 22281 27625 22293 27659
rect 22327 27656 22339 27659
rect 22370 27656 22376 27668
rect 22327 27628 22376 27656
rect 22327 27625 22339 27628
rect 22281 27619 22339 27625
rect 22370 27616 22376 27628
rect 22428 27616 22434 27668
rect 25590 27616 25596 27668
rect 25648 27616 25654 27668
rect 34514 27616 34520 27668
rect 34572 27616 34578 27668
rect 23937 27591 23995 27597
rect 23937 27588 23949 27591
rect 22204 27560 23949 27588
rect 17359 27492 18092 27520
rect 17359 27489 17371 27492
rect 17313 27483 17371 27489
rect 22462 27480 22468 27532
rect 22520 27520 22526 27532
rect 23400 27520 23428 27560
rect 23937 27557 23949 27560
rect 23983 27557 23995 27591
rect 23937 27551 23995 27557
rect 24210 27548 24216 27600
rect 24268 27588 24274 27600
rect 31846 27588 31852 27600
rect 24268 27560 31852 27588
rect 24268 27548 24274 27560
rect 31846 27548 31852 27560
rect 31904 27548 31910 27600
rect 23750 27520 23756 27532
rect 22520 27492 23336 27520
rect 23400 27492 23520 27520
rect 22520 27480 22526 27492
rect 11900 27424 12848 27452
rect 13449 27455 13507 27461
rect 13449 27421 13461 27455
rect 13495 27452 13507 27455
rect 14274 27452 14280 27464
rect 13495 27424 14280 27452
rect 13495 27421 13507 27424
rect 13449 27415 13507 27421
rect 14274 27412 14280 27424
rect 14332 27412 14338 27464
rect 14550 27412 14556 27464
rect 14608 27412 14614 27464
rect 16022 27452 16028 27464
rect 14752 27424 16028 27452
rect 9852 27387 9910 27393
rect 9324 27356 9812 27384
rect 8435 27353 8447 27356
rect 8389 27347 8447 27353
rect 9784 27328 9812 27356
rect 9852 27353 9864 27387
rect 9898 27384 9910 27387
rect 10134 27384 10140 27396
rect 9898 27356 10140 27384
rect 9898 27353 9910 27356
rect 9852 27347 9910 27353
rect 10134 27344 10140 27356
rect 10192 27344 10198 27396
rect 11701 27387 11759 27393
rect 11701 27353 11713 27387
rect 11747 27384 11759 27387
rect 12894 27384 12900 27396
rect 11747 27356 12900 27384
rect 11747 27353 11759 27356
rect 11701 27347 11759 27353
rect 12894 27344 12900 27356
rect 12952 27344 12958 27396
rect 13541 27387 13599 27393
rect 13541 27353 13553 27387
rect 13587 27384 13599 27387
rect 14752 27384 14780 27424
rect 16022 27412 16028 27424
rect 16080 27412 16086 27464
rect 16206 27412 16212 27464
rect 16264 27412 16270 27464
rect 16390 27412 16396 27464
rect 16448 27412 16454 27464
rect 17129 27455 17187 27461
rect 17129 27421 17141 27455
rect 17175 27452 17187 27455
rect 18046 27452 18052 27464
rect 17175 27424 18052 27452
rect 17175 27421 17187 27424
rect 17129 27415 17187 27421
rect 17328 27396 17356 27424
rect 18046 27412 18052 27424
rect 18104 27412 18110 27464
rect 19061 27455 19119 27461
rect 19061 27421 19073 27455
rect 19107 27452 19119 27455
rect 19245 27455 19303 27461
rect 19245 27452 19257 27455
rect 19107 27424 19257 27452
rect 19107 27421 19119 27424
rect 19061 27415 19119 27421
rect 19245 27421 19257 27424
rect 19291 27452 19303 27455
rect 20901 27455 20959 27461
rect 20901 27452 20913 27455
rect 19291 27424 20913 27452
rect 19291 27421 19303 27424
rect 19245 27415 19303 27421
rect 20901 27421 20913 27424
rect 20947 27452 20959 27455
rect 20947 27424 22048 27452
rect 20947 27421 20959 27424
rect 20901 27415 20959 27421
rect 13587 27356 14780 27384
rect 14820 27387 14878 27393
rect 13587 27353 13599 27356
rect 13541 27347 13599 27353
rect 14820 27353 14832 27387
rect 14866 27384 14878 27387
rect 15102 27384 15108 27396
rect 14866 27356 15108 27384
rect 14866 27353 14878 27356
rect 14820 27347 14878 27353
rect 15102 27344 15108 27356
rect 15160 27344 15166 27396
rect 16301 27387 16359 27393
rect 16301 27353 16313 27387
rect 16347 27353 16359 27387
rect 16301 27347 16359 27353
rect 3878 27276 3884 27328
rect 3936 27276 3942 27328
rect 4338 27276 4344 27328
rect 4396 27276 4402 27328
rect 4614 27276 4620 27328
rect 4672 27316 4678 27328
rect 4890 27316 4896 27328
rect 4672 27288 4896 27316
rect 4672 27276 4678 27288
rect 4890 27276 4896 27288
rect 4948 27276 4954 27328
rect 8018 27276 8024 27328
rect 8076 27276 8082 27328
rect 9766 27276 9772 27328
rect 9824 27276 9830 27328
rect 10962 27276 10968 27328
rect 11020 27276 11026 27328
rect 11606 27276 11612 27328
rect 11664 27316 11670 27328
rect 12345 27319 12403 27325
rect 12345 27316 12357 27319
rect 11664 27288 12357 27316
rect 11664 27276 11670 27288
rect 12345 27285 12357 27288
rect 12391 27316 12403 27319
rect 12618 27316 12624 27328
rect 12391 27288 12624 27316
rect 12391 27285 12403 27288
rect 12345 27279 12403 27285
rect 12618 27276 12624 27288
rect 12676 27276 12682 27328
rect 13906 27276 13912 27328
rect 13964 27276 13970 27328
rect 14090 27276 14096 27328
rect 14148 27276 14154 27328
rect 14274 27276 14280 27328
rect 14332 27316 14338 27328
rect 15010 27316 15016 27328
rect 14332 27288 15016 27316
rect 14332 27276 14338 27288
rect 15010 27276 15016 27288
rect 15068 27276 15074 27328
rect 15930 27276 15936 27328
rect 15988 27316 15994 27328
rect 16316 27316 16344 27347
rect 17310 27344 17316 27396
rect 17368 27344 17374 27396
rect 18816 27387 18874 27393
rect 18816 27353 18828 27387
rect 18862 27384 18874 27387
rect 18966 27384 18972 27396
rect 18862 27356 18972 27384
rect 18862 27353 18874 27356
rect 18816 27347 18874 27353
rect 18966 27344 18972 27356
rect 19024 27344 19030 27396
rect 19512 27387 19570 27393
rect 19512 27353 19524 27387
rect 19558 27384 19570 27387
rect 19702 27384 19708 27396
rect 19558 27356 19708 27384
rect 19558 27353 19570 27356
rect 19512 27347 19570 27353
rect 19702 27344 19708 27356
rect 19760 27344 19766 27396
rect 21168 27387 21226 27393
rect 21168 27353 21180 27387
rect 21214 27384 21226 27387
rect 21450 27384 21456 27396
rect 21214 27356 21456 27384
rect 21214 27353 21226 27356
rect 21168 27347 21226 27353
rect 21450 27344 21456 27356
rect 21508 27344 21514 27396
rect 22020 27384 22048 27424
rect 22094 27412 22100 27464
rect 22152 27452 22158 27464
rect 22373 27455 22431 27461
rect 22373 27452 22385 27455
rect 22152 27424 22385 27452
rect 22152 27412 22158 27424
rect 22373 27421 22385 27424
rect 22419 27421 22431 27455
rect 22373 27415 22431 27421
rect 22646 27412 22652 27464
rect 22704 27452 22710 27464
rect 23198 27452 23204 27464
rect 22704 27424 23204 27452
rect 22704 27412 22710 27424
rect 23198 27412 23204 27424
rect 23256 27412 23262 27464
rect 23308 27461 23336 27492
rect 23492 27461 23520 27492
rect 23584 27492 23756 27520
rect 23584 27461 23612 27492
rect 23750 27480 23756 27492
rect 23808 27480 23814 27532
rect 26142 27480 26148 27532
rect 26200 27520 26206 27532
rect 27522 27520 27528 27532
rect 26200 27492 27528 27520
rect 26200 27480 26206 27492
rect 27522 27480 27528 27492
rect 27580 27480 27586 27532
rect 28718 27480 28724 27532
rect 28776 27520 28782 27532
rect 29270 27520 29276 27532
rect 28776 27492 29276 27520
rect 28776 27480 28782 27492
rect 29270 27480 29276 27492
rect 29328 27480 29334 27532
rect 30098 27480 30104 27532
rect 30156 27480 30162 27532
rect 31754 27520 31760 27532
rect 31588 27492 31760 27520
rect 23293 27455 23351 27461
rect 23293 27421 23305 27455
rect 23339 27421 23351 27455
rect 23293 27415 23351 27421
rect 23477 27455 23535 27461
rect 23477 27421 23489 27455
rect 23523 27421 23535 27455
rect 23477 27415 23535 27421
rect 23569 27455 23627 27461
rect 23569 27421 23581 27455
rect 23615 27421 23627 27455
rect 23569 27415 23627 27421
rect 23658 27412 23664 27464
rect 23716 27452 23722 27464
rect 24121 27455 24179 27461
rect 24121 27452 24133 27455
rect 23716 27424 24133 27452
rect 23716 27412 23722 27424
rect 24121 27421 24133 27424
rect 24167 27421 24179 27455
rect 24121 27415 24179 27421
rect 25961 27455 26019 27461
rect 25961 27421 25973 27455
rect 26007 27452 26019 27455
rect 26418 27452 26424 27464
rect 26007 27424 26424 27452
rect 26007 27421 26019 27424
rect 25961 27415 26019 27421
rect 26418 27412 26424 27424
rect 26476 27412 26482 27464
rect 27154 27412 27160 27464
rect 27212 27412 27218 27464
rect 27430 27412 27436 27464
rect 27488 27412 27494 27464
rect 27893 27455 27951 27461
rect 27893 27421 27905 27455
rect 27939 27452 27951 27455
rect 28905 27455 28963 27461
rect 27939 27424 28028 27452
rect 27939 27421 27951 27424
rect 27893 27415 27951 27421
rect 22278 27384 22284 27396
rect 22020 27356 22284 27384
rect 22278 27344 22284 27356
rect 22336 27344 22342 27396
rect 25409 27387 25467 27393
rect 25409 27384 25421 27387
rect 23768 27356 25421 27384
rect 15988 27288 16344 27316
rect 15988 27276 15994 27288
rect 16574 27276 16580 27328
rect 16632 27276 16638 27328
rect 16758 27276 16764 27328
rect 16816 27316 16822 27328
rect 17218 27316 17224 27328
rect 16816 27288 17224 27316
rect 16816 27276 16822 27288
rect 17218 27276 17224 27288
rect 17276 27276 17282 27328
rect 17494 27276 17500 27328
rect 17552 27316 17558 27328
rect 17681 27319 17739 27325
rect 17681 27316 17693 27319
rect 17552 27288 17693 27316
rect 17552 27276 17558 27288
rect 17681 27285 17693 27288
rect 17727 27285 17739 27319
rect 17681 27279 17739 27285
rect 17770 27276 17776 27328
rect 17828 27316 17834 27328
rect 23768 27316 23796 27356
rect 25409 27353 25421 27356
rect 25455 27384 25467 27387
rect 26053 27387 26111 27393
rect 26053 27384 26065 27387
rect 25455 27356 26065 27384
rect 25455 27353 25467 27356
rect 25409 27347 25467 27353
rect 26053 27353 26065 27356
rect 26099 27384 26111 27387
rect 26510 27384 26516 27396
rect 26099 27356 26516 27384
rect 26099 27353 26111 27356
rect 26053 27347 26111 27353
rect 26510 27344 26516 27356
rect 26568 27344 26574 27396
rect 27172 27384 27200 27412
rect 27172 27356 27752 27384
rect 17828 27288 23796 27316
rect 17828 27276 17834 27288
rect 23842 27276 23848 27328
rect 23900 27276 23906 27328
rect 26970 27276 26976 27328
rect 27028 27316 27034 27328
rect 27249 27319 27307 27325
rect 27249 27316 27261 27319
rect 27028 27288 27261 27316
rect 27028 27276 27034 27288
rect 27249 27285 27261 27288
rect 27295 27285 27307 27319
rect 27249 27279 27307 27285
rect 27614 27276 27620 27328
rect 27672 27276 27678 27328
rect 27724 27325 27752 27356
rect 28000 27328 28028 27424
rect 28905 27421 28917 27455
rect 28951 27452 28963 27455
rect 28997 27455 29055 27461
rect 28997 27452 29009 27455
rect 28951 27424 29009 27452
rect 28951 27421 28963 27424
rect 28905 27415 28963 27421
rect 28997 27421 29009 27424
rect 29043 27452 29055 27455
rect 29086 27452 29092 27464
rect 29043 27424 29092 27452
rect 29043 27421 29055 27424
rect 28997 27415 29055 27421
rect 29086 27412 29092 27424
rect 29144 27412 29150 27464
rect 29181 27455 29239 27461
rect 29181 27421 29193 27455
rect 29227 27452 29239 27455
rect 31478 27452 31484 27464
rect 29227 27424 31484 27452
rect 29227 27421 29239 27424
rect 29181 27415 29239 27421
rect 28629 27387 28687 27393
rect 28629 27353 28641 27387
rect 28675 27384 28687 27387
rect 29196 27384 29224 27415
rect 31478 27412 31484 27424
rect 31536 27412 31542 27464
rect 31588 27461 31616 27492
rect 31754 27480 31760 27492
rect 31812 27520 31818 27532
rect 32766 27520 32772 27532
rect 31812 27492 32772 27520
rect 31812 27480 31818 27492
rect 32766 27480 32772 27492
rect 32824 27480 32830 27532
rect 31573 27455 31631 27461
rect 31573 27421 31585 27455
rect 31619 27421 31631 27455
rect 31573 27415 31631 27421
rect 30098 27384 30104 27396
rect 28675 27356 29224 27384
rect 29380 27356 30104 27384
rect 28675 27353 28687 27356
rect 28629 27347 28687 27353
rect 27709 27319 27767 27325
rect 27709 27285 27721 27319
rect 27755 27285 27767 27319
rect 27709 27279 27767 27285
rect 27982 27276 27988 27328
rect 28040 27276 28046 27328
rect 28718 27276 28724 27328
rect 28776 27276 28782 27328
rect 29380 27325 29408 27356
rect 30098 27344 30104 27356
rect 30156 27344 30162 27396
rect 33045 27387 33103 27393
rect 33045 27353 33057 27387
rect 33091 27384 33103 27387
rect 33318 27384 33324 27396
rect 33091 27356 33324 27384
rect 33091 27353 33103 27356
rect 33045 27347 33103 27353
rect 33318 27344 33324 27356
rect 33376 27344 33382 27396
rect 34054 27344 34060 27396
rect 34112 27344 34118 27396
rect 29365 27319 29423 27325
rect 29365 27285 29377 27319
rect 29411 27285 29423 27319
rect 29365 27279 29423 27285
rect 29549 27319 29607 27325
rect 29549 27285 29561 27319
rect 29595 27316 29607 27319
rect 29638 27316 29644 27328
rect 29595 27288 29644 27316
rect 29595 27285 29607 27288
rect 29549 27279 29607 27285
rect 29638 27276 29644 27288
rect 29696 27276 29702 27328
rect 29914 27276 29920 27328
rect 29972 27276 29978 27328
rect 30006 27276 30012 27328
rect 30064 27276 30070 27328
rect 1104 27226 35328 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35328 27226
rect 1104 27152 35328 27174
rect 2590 27072 2596 27124
rect 2648 27072 2654 27124
rect 2961 27115 3019 27121
rect 2961 27081 2973 27115
rect 3007 27112 3019 27115
rect 4154 27112 4160 27124
rect 3007 27084 4160 27112
rect 3007 27081 3019 27084
rect 2961 27075 3019 27081
rect 4154 27072 4160 27084
rect 4212 27072 4218 27124
rect 4338 27072 4344 27124
rect 4396 27112 4402 27124
rect 4706 27112 4712 27124
rect 4396 27084 4712 27112
rect 4396 27072 4402 27084
rect 4706 27072 4712 27084
rect 4764 27112 4770 27124
rect 4801 27115 4859 27121
rect 4801 27112 4813 27115
rect 4764 27084 4813 27112
rect 4764 27072 4770 27084
rect 4801 27081 4813 27084
rect 4847 27081 4859 27115
rect 4801 27075 4859 27081
rect 6822 27072 6828 27124
rect 6880 27072 6886 27124
rect 7193 27115 7251 27121
rect 7193 27081 7205 27115
rect 7239 27112 7251 27115
rect 7466 27112 7472 27124
rect 7239 27084 7472 27112
rect 7239 27081 7251 27084
rect 7193 27075 7251 27081
rect 7466 27072 7472 27084
rect 7524 27072 7530 27124
rect 9214 27072 9220 27124
rect 9272 27112 9278 27124
rect 9309 27115 9367 27121
rect 9309 27112 9321 27115
rect 9272 27084 9321 27112
rect 9272 27072 9278 27084
rect 9309 27081 9321 27084
rect 9355 27081 9367 27115
rect 9309 27075 9367 27081
rect 10134 27072 10140 27124
rect 10192 27072 10198 27124
rect 10505 27115 10563 27121
rect 10505 27081 10517 27115
rect 10551 27112 10563 27115
rect 10962 27112 10968 27124
rect 10551 27084 10968 27112
rect 10551 27081 10563 27084
rect 10505 27075 10563 27081
rect 10962 27072 10968 27084
rect 11020 27112 11026 27124
rect 11020 27084 12112 27112
rect 11020 27072 11026 27084
rect 3688 27047 3746 27053
rect 3688 27013 3700 27047
rect 3734 27044 3746 27047
rect 3878 27044 3884 27056
rect 3734 27016 3884 27044
rect 3734 27013 3746 27016
rect 3688 27007 3746 27013
rect 3878 27004 3884 27016
rect 3936 27004 3942 27056
rect 4246 27004 4252 27056
rect 4304 27044 4310 27056
rect 4982 27044 4988 27056
rect 4304 27016 4988 27044
rect 4304 27004 4310 27016
rect 4982 27004 4988 27016
rect 5040 27004 5046 27056
rect 6178 27004 6184 27056
rect 6236 27044 6242 27056
rect 9582 27044 9588 27056
rect 6236 27016 9588 27044
rect 6236 27004 6242 27016
rect 7190 26936 7196 26988
rect 7248 26976 7254 26988
rect 7285 26979 7343 26985
rect 7285 26976 7297 26979
rect 7248 26948 7297 26976
rect 7248 26936 7254 26948
rect 7285 26945 7297 26948
rect 7331 26945 7343 26979
rect 7285 26939 7343 26945
rect 7374 26936 7380 26988
rect 7432 26976 7438 26988
rect 7944 26985 7972 27016
rect 9582 27004 9588 27016
rect 9640 27004 9646 27056
rect 11606 27044 11612 27056
rect 9968 27016 11612 27044
rect 7929 26979 7987 26985
rect 7432 26948 7512 26976
rect 7432 26936 7438 26948
rect 3050 26868 3056 26920
rect 3108 26868 3114 26920
rect 3237 26911 3295 26917
rect 3237 26877 3249 26911
rect 3283 26908 3295 26911
rect 3283 26880 3372 26908
rect 3283 26877 3295 26880
rect 3237 26871 3295 26877
rect 3344 26772 3372 26880
rect 3418 26868 3424 26920
rect 3476 26868 3482 26920
rect 7484 26917 7512 26948
rect 7929 26945 7941 26979
rect 7975 26945 7987 26979
rect 7929 26939 7987 26945
rect 8018 26936 8024 26988
rect 8076 26976 8082 26988
rect 8185 26979 8243 26985
rect 8185 26976 8197 26979
rect 8076 26948 8197 26976
rect 8076 26936 8082 26948
rect 8185 26945 8197 26948
rect 8231 26945 8243 26979
rect 8185 26939 8243 26945
rect 9030 26936 9036 26988
rect 9088 26976 9094 26988
rect 9968 26976 9996 27016
rect 11606 27004 11612 27016
rect 11664 27044 11670 27056
rect 11664 27016 11744 27044
rect 11664 27004 11670 27016
rect 9088 26948 9996 26976
rect 10045 26979 10103 26985
rect 9088 26936 9094 26948
rect 10045 26945 10057 26979
rect 10091 26976 10103 26979
rect 10594 26976 10600 26988
rect 10091 26948 10600 26976
rect 10091 26945 10103 26948
rect 10045 26939 10103 26945
rect 7469 26911 7527 26917
rect 7469 26877 7481 26911
rect 7515 26877 7527 26911
rect 7469 26871 7527 26877
rect 8938 26868 8944 26920
rect 8996 26908 9002 26920
rect 10060 26908 10088 26939
rect 10594 26936 10600 26948
rect 10652 26936 10658 26988
rect 11716 26985 11744 27016
rect 11790 27004 11796 27056
rect 11848 27004 11854 27056
rect 11885 27047 11943 27053
rect 11885 27013 11897 27047
rect 11931 27044 11943 27047
rect 11974 27044 11980 27056
rect 11931 27016 11980 27044
rect 11931 27013 11943 27016
rect 11885 27007 11943 27013
rect 11974 27004 11980 27016
rect 12032 27004 12038 27056
rect 12084 26985 12112 27084
rect 12342 27072 12348 27124
rect 12400 27072 12406 27124
rect 12618 27072 12624 27124
rect 12676 27112 12682 27124
rect 14737 27115 14795 27121
rect 12676 27084 14044 27112
rect 12676 27072 12682 27084
rect 11701 26979 11759 26985
rect 11701 26945 11713 26979
rect 11747 26945 11759 26979
rect 11701 26939 11759 26945
rect 12069 26979 12127 26985
rect 12069 26945 12081 26979
rect 12115 26945 12127 26979
rect 12360 26976 12388 27072
rect 12802 27004 12808 27056
rect 12860 27044 12866 27056
rect 13265 27047 13323 27053
rect 13265 27044 13277 27047
rect 12860 27016 13277 27044
rect 12860 27004 12866 27016
rect 13265 27013 13277 27016
rect 13311 27044 13323 27047
rect 13446 27044 13452 27056
rect 13311 27016 13452 27044
rect 13311 27013 13323 27016
rect 13265 27007 13323 27013
rect 13446 27004 13452 27016
rect 13504 27004 13510 27056
rect 13624 27047 13682 27053
rect 13624 27013 13636 27047
rect 13670 27044 13682 27047
rect 13906 27044 13912 27056
rect 13670 27016 13912 27044
rect 13670 27013 13682 27016
rect 13624 27007 13682 27013
rect 13906 27004 13912 27016
rect 13964 27004 13970 27056
rect 14016 27044 14044 27084
rect 14737 27081 14749 27115
rect 14783 27112 14795 27115
rect 16022 27112 16028 27124
rect 14783 27084 16028 27112
rect 14783 27081 14795 27084
rect 14737 27075 14795 27081
rect 16022 27072 16028 27084
rect 16080 27072 16086 27124
rect 17034 27072 17040 27124
rect 17092 27072 17098 27124
rect 18601 27115 18659 27121
rect 18601 27112 18613 27115
rect 17512 27084 18613 27112
rect 17512 27056 17540 27084
rect 18601 27081 18613 27084
rect 18647 27081 18659 27115
rect 18601 27075 18659 27081
rect 18966 27072 18972 27124
rect 19024 27072 19030 27124
rect 23474 27072 23480 27124
rect 23532 27112 23538 27124
rect 26605 27115 26663 27121
rect 26605 27112 26617 27115
rect 23532 27084 26617 27112
rect 23532 27072 23538 27084
rect 26605 27081 26617 27084
rect 26651 27112 26663 27115
rect 26694 27112 26700 27124
rect 26651 27084 26700 27112
rect 26651 27081 26663 27084
rect 26605 27075 26663 27081
rect 26694 27072 26700 27084
rect 26752 27072 26758 27124
rect 26970 27072 26976 27124
rect 27028 27072 27034 27124
rect 28537 27115 28595 27121
rect 28537 27081 28549 27115
rect 28583 27112 28595 27115
rect 29178 27112 29184 27124
rect 28583 27084 29184 27112
rect 28583 27081 28595 27084
rect 28537 27075 28595 27081
rect 29178 27072 29184 27084
rect 29236 27112 29242 27124
rect 30006 27112 30012 27124
rect 29236 27084 30012 27112
rect 29236 27072 29242 27084
rect 30006 27072 30012 27084
rect 30064 27072 30070 27124
rect 33318 27072 33324 27124
rect 33376 27112 33382 27124
rect 33781 27115 33839 27121
rect 33781 27112 33793 27115
rect 33376 27084 33793 27112
rect 33376 27072 33382 27084
rect 33781 27081 33793 27084
rect 33827 27081 33839 27115
rect 33781 27075 33839 27081
rect 34149 27115 34207 27121
rect 34149 27081 34161 27115
rect 34195 27112 34207 27115
rect 34514 27112 34520 27124
rect 34195 27084 34520 27112
rect 34195 27081 34207 27084
rect 34149 27075 34207 27081
rect 34514 27072 34520 27084
rect 34572 27072 34578 27124
rect 15933 27047 15991 27053
rect 15933 27044 15945 27047
rect 14016 27016 15945 27044
rect 15933 27013 15945 27016
rect 15979 27044 15991 27047
rect 16206 27044 16212 27056
rect 15979 27016 16212 27044
rect 15979 27013 15991 27016
rect 15933 27007 15991 27013
rect 16206 27004 16212 27016
rect 16264 27004 16270 27056
rect 17494 27004 17500 27056
rect 17552 27004 17558 27056
rect 19996 27016 20944 27044
rect 19996 26988 20024 27016
rect 12575 26979 12633 26985
rect 12575 26976 12587 26979
rect 12360 26948 12587 26976
rect 12069 26939 12127 26945
rect 12575 26945 12587 26948
rect 12621 26945 12633 26979
rect 12575 26939 12633 26945
rect 12710 26936 12716 26988
rect 12768 26936 12774 26988
rect 12986 26936 12992 26988
rect 13044 26936 13050 26988
rect 13078 26936 13084 26988
rect 13136 26936 13142 26988
rect 14550 26936 14556 26988
rect 14608 26976 14614 26988
rect 14826 26976 14832 26988
rect 14608 26948 14832 26976
rect 14608 26936 14614 26948
rect 14826 26936 14832 26948
rect 14884 26936 14890 26988
rect 16574 26936 16580 26988
rect 16632 26976 16638 26988
rect 17310 26985 17316 26988
rect 17129 26979 17187 26985
rect 17129 26976 17141 26979
rect 16632 26948 17141 26976
rect 16632 26936 16638 26948
rect 17129 26945 17141 26948
rect 17175 26945 17187 26979
rect 17129 26939 17187 26945
rect 17277 26979 17316 26985
rect 17277 26945 17289 26979
rect 17277 26939 17316 26945
rect 17310 26936 17316 26939
rect 17368 26936 17374 26988
rect 17402 26936 17408 26988
rect 17460 26936 17466 26988
rect 17594 26979 17652 26985
rect 17594 26976 17606 26979
rect 17512 26948 17606 26976
rect 8996 26880 10088 26908
rect 8996 26868 9002 26880
rect 10410 26868 10416 26920
rect 10468 26908 10474 26920
rect 10689 26911 10747 26917
rect 10689 26908 10701 26911
rect 10468 26880 10701 26908
rect 10468 26868 10474 26880
rect 10689 26877 10701 26880
rect 10735 26877 10747 26911
rect 10689 26871 10747 26877
rect 9122 26800 9128 26852
rect 9180 26840 9186 26852
rect 9180 26812 9904 26840
rect 9180 26800 9186 26812
rect 3694 26772 3700 26784
rect 3344 26744 3700 26772
rect 3694 26732 3700 26744
rect 3752 26732 3758 26784
rect 4522 26732 4528 26784
rect 4580 26772 4586 26784
rect 4706 26772 4712 26784
rect 4580 26744 4712 26772
rect 4580 26732 4586 26744
rect 4706 26732 4712 26744
rect 4764 26732 4770 26784
rect 4982 26732 4988 26784
rect 5040 26732 5046 26784
rect 9677 26775 9735 26781
rect 9677 26741 9689 26775
rect 9723 26772 9735 26775
rect 9766 26772 9772 26784
rect 9723 26744 9772 26772
rect 9723 26741 9735 26744
rect 9677 26735 9735 26741
rect 9766 26732 9772 26744
rect 9824 26732 9830 26784
rect 9876 26781 9904 26812
rect 9861 26775 9919 26781
rect 9861 26741 9873 26775
rect 9907 26772 9919 26775
rect 10502 26772 10508 26784
rect 9907 26744 10508 26772
rect 9907 26741 9919 26744
rect 9861 26735 9919 26741
rect 10502 26732 10508 26744
rect 10560 26732 10566 26784
rect 10704 26772 10732 26871
rect 13354 26868 13360 26920
rect 13412 26868 13418 26920
rect 17034 26868 17040 26920
rect 17092 26908 17098 26920
rect 17512 26908 17540 26948
rect 17594 26945 17606 26948
rect 17640 26945 17652 26979
rect 17594 26939 17652 26945
rect 18046 26936 18052 26988
rect 18104 26976 18110 26988
rect 18141 26979 18199 26985
rect 18141 26976 18153 26979
rect 18104 26948 18153 26976
rect 18104 26936 18110 26948
rect 18141 26945 18153 26948
rect 18187 26976 18199 26979
rect 19794 26976 19800 26988
rect 18187 26948 19800 26976
rect 18187 26945 18199 26948
rect 18141 26939 18199 26945
rect 19794 26936 19800 26948
rect 19852 26936 19858 26988
rect 19978 26936 19984 26988
rect 20036 26936 20042 26988
rect 20162 26936 20168 26988
rect 20220 26936 20226 26988
rect 20530 26936 20536 26988
rect 20588 26936 20594 26988
rect 17092 26880 17540 26908
rect 17092 26868 17098 26880
rect 17954 26868 17960 26920
rect 18012 26908 18018 26920
rect 18325 26911 18383 26917
rect 18325 26908 18337 26911
rect 18012 26880 18337 26908
rect 18012 26868 18018 26880
rect 18325 26877 18337 26880
rect 18371 26877 18383 26911
rect 18325 26871 18383 26877
rect 18509 26911 18567 26917
rect 18509 26877 18521 26911
rect 18555 26877 18567 26911
rect 18509 26871 18567 26877
rect 14734 26800 14740 26852
rect 14792 26840 14798 26852
rect 16025 26843 16083 26849
rect 16025 26840 16037 26843
rect 14792 26812 16037 26840
rect 14792 26800 14798 26812
rect 16025 26809 16037 26812
rect 16071 26840 16083 26843
rect 16390 26840 16396 26852
rect 16071 26812 16396 26840
rect 16071 26809 16083 26812
rect 16025 26803 16083 26809
rect 16390 26800 16396 26812
rect 16448 26800 16454 26852
rect 18524 26840 18552 26871
rect 20254 26868 20260 26920
rect 20312 26868 20318 26920
rect 20916 26917 20944 27016
rect 21818 27004 21824 27056
rect 21876 27004 21882 27056
rect 22388 27016 24072 27044
rect 22005 26979 22063 26985
rect 22005 26945 22017 26979
rect 22051 26945 22063 26979
rect 22005 26939 22063 26945
rect 20349 26911 20407 26917
rect 20349 26877 20361 26911
rect 20395 26877 20407 26911
rect 20349 26871 20407 26877
rect 20901 26911 20959 26917
rect 20901 26877 20913 26911
rect 20947 26908 20959 26911
rect 20990 26908 20996 26920
rect 20947 26880 20996 26908
rect 20947 26877 20959 26880
rect 20901 26871 20959 26877
rect 20364 26840 20392 26871
rect 20990 26868 20996 26880
rect 21048 26868 21054 26920
rect 21085 26843 21143 26849
rect 21085 26840 21097 26843
rect 17628 26812 18552 26840
rect 19306 26812 21097 26840
rect 11057 26775 11115 26781
rect 11057 26772 11069 26775
rect 10704 26744 11069 26772
rect 11057 26741 11069 26744
rect 11103 26772 11115 26775
rect 11146 26772 11152 26784
rect 11103 26744 11152 26772
rect 11103 26741 11115 26744
rect 11057 26735 11115 26741
rect 11146 26732 11152 26744
rect 11204 26732 11210 26784
rect 11514 26732 11520 26784
rect 11572 26732 11578 26784
rect 12342 26732 12348 26784
rect 12400 26772 12406 26784
rect 12437 26775 12495 26781
rect 12437 26772 12449 26775
rect 12400 26744 12449 26772
rect 12400 26732 12406 26744
rect 12437 26741 12449 26744
rect 12483 26741 12495 26775
rect 12437 26735 12495 26741
rect 16758 26732 16764 26784
rect 16816 26772 16822 26784
rect 17628 26772 17656 26812
rect 16816 26744 17656 26772
rect 16816 26732 16822 26744
rect 17770 26732 17776 26784
rect 17828 26732 17834 26784
rect 17862 26732 17868 26784
rect 17920 26772 17926 26784
rect 19306 26772 19334 26812
rect 21085 26809 21097 26812
rect 21131 26809 21143 26843
rect 21085 26803 21143 26809
rect 21818 26800 21824 26852
rect 21876 26840 21882 26852
rect 22020 26840 22048 26939
rect 22278 26868 22284 26920
rect 22336 26908 22342 26920
rect 22388 26908 22416 27016
rect 22548 26979 22606 26985
rect 22548 26945 22560 26979
rect 22594 26976 22606 26979
rect 22830 26976 22836 26988
rect 22594 26948 22836 26976
rect 22594 26945 22606 26948
rect 22548 26939 22606 26945
rect 22830 26936 22836 26948
rect 22888 26936 22894 26988
rect 24044 26985 24072 27016
rect 25498 27004 25504 27056
rect 25556 27004 25562 27056
rect 30098 27044 30104 27056
rect 28368 27016 30104 27044
rect 24029 26979 24087 26985
rect 24029 26945 24041 26979
rect 24075 26976 24087 26979
rect 24118 26976 24124 26988
rect 24075 26948 24124 26976
rect 24075 26945 24087 26948
rect 24029 26939 24087 26945
rect 24118 26936 24124 26948
rect 24176 26936 24182 26988
rect 24296 26979 24354 26985
rect 24296 26945 24308 26979
rect 24342 26976 24354 26979
rect 24578 26976 24584 26988
rect 24342 26948 24584 26976
rect 24342 26945 24354 26948
rect 24296 26939 24354 26945
rect 24578 26936 24584 26948
rect 24636 26936 24642 26988
rect 26326 26936 26332 26988
rect 26384 26976 26390 26988
rect 26697 26979 26755 26985
rect 26697 26976 26709 26979
rect 26384 26948 26709 26976
rect 26384 26936 26390 26948
rect 26697 26945 26709 26948
rect 26743 26945 26755 26979
rect 26697 26939 26755 26945
rect 27338 26936 27344 26988
rect 27396 26976 27402 26988
rect 28368 26985 28396 27016
rect 28086 26979 28144 26985
rect 28086 26976 28098 26979
rect 27396 26948 28098 26976
rect 27396 26936 27402 26948
rect 28086 26945 28098 26948
rect 28132 26945 28144 26979
rect 28086 26939 28144 26945
rect 28353 26979 28411 26985
rect 28353 26945 28365 26979
rect 28399 26945 28411 26979
rect 28353 26939 28411 26945
rect 29638 26936 29644 26988
rect 29696 26985 29702 26988
rect 29932 26985 29960 27016
rect 30098 27004 30104 27016
rect 30156 27044 30162 27056
rect 31754 27044 31760 27056
rect 30156 27016 31760 27044
rect 30156 27004 30162 27016
rect 31754 27004 31760 27016
rect 31812 27004 31818 27056
rect 29696 26976 29708 26985
rect 29917 26979 29975 26985
rect 29696 26948 29741 26976
rect 29696 26939 29708 26948
rect 29917 26945 29929 26979
rect 29963 26945 29975 26979
rect 29917 26939 29975 26945
rect 29696 26936 29702 26939
rect 30374 26936 30380 26988
rect 30432 26976 30438 26988
rect 30929 26979 30987 26985
rect 30929 26976 30941 26979
rect 30432 26948 30941 26976
rect 30432 26936 30438 26948
rect 30929 26945 30941 26948
rect 30975 26976 30987 26979
rect 31021 26979 31079 26985
rect 31021 26976 31033 26979
rect 30975 26948 31033 26976
rect 30975 26945 30987 26948
rect 30929 26939 30987 26945
rect 31021 26945 31033 26948
rect 31067 26945 31079 26979
rect 31021 26939 31079 26945
rect 33962 26936 33968 26988
rect 34020 26936 34026 26988
rect 34238 26936 34244 26988
rect 34296 26936 34302 26988
rect 34514 26936 34520 26988
rect 34572 26936 34578 26988
rect 22336 26880 22416 26908
rect 22336 26868 22342 26880
rect 34790 26868 34796 26920
rect 34848 26868 34854 26920
rect 21876 26812 22048 26840
rect 23584 26812 24073 26840
rect 21876 26800 21882 26812
rect 17920 26744 19334 26772
rect 20717 26775 20775 26781
rect 17920 26732 17926 26744
rect 20717 26741 20729 26775
rect 20763 26772 20775 26775
rect 23584 26772 23612 26812
rect 20763 26744 23612 26772
rect 20763 26741 20775 26744
rect 20717 26735 20775 26741
rect 23658 26732 23664 26784
rect 23716 26732 23722 26784
rect 24045 26772 24073 26812
rect 24210 26772 24216 26784
rect 24045 26744 24216 26772
rect 24210 26732 24216 26744
rect 24268 26732 24274 26784
rect 25406 26732 25412 26784
rect 25464 26732 25470 26784
rect 26326 26732 26332 26784
rect 26384 26732 26390 26784
rect 26602 26732 26608 26784
rect 26660 26772 26666 26784
rect 30282 26772 30288 26784
rect 26660 26744 30288 26772
rect 26660 26732 26666 26744
rect 30282 26732 30288 26744
rect 30340 26732 30346 26784
rect 1104 26682 35328 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 35328 26682
rect 1104 26608 35328 26630
rect 5353 26571 5411 26577
rect 5353 26537 5365 26571
rect 5399 26568 5411 26571
rect 5442 26568 5448 26580
rect 5399 26540 5448 26568
rect 5399 26537 5411 26540
rect 5353 26531 5411 26537
rect 5442 26528 5448 26540
rect 5500 26528 5506 26580
rect 5718 26528 5724 26580
rect 5776 26528 5782 26580
rect 9766 26528 9772 26580
rect 9824 26568 9830 26580
rect 9950 26568 9956 26580
rect 9824 26540 9956 26568
rect 9824 26528 9830 26540
rect 9950 26528 9956 26540
rect 10008 26528 10014 26580
rect 11517 26571 11575 26577
rect 11517 26537 11529 26571
rect 11563 26568 11575 26571
rect 12342 26568 12348 26580
rect 11563 26540 12348 26568
rect 11563 26537 11575 26540
rect 11517 26531 11575 26537
rect 12342 26528 12348 26540
rect 12400 26528 12406 26580
rect 12710 26568 12716 26580
rect 12544 26540 12716 26568
rect 4982 26460 4988 26512
rect 5040 26500 5046 26512
rect 5258 26500 5264 26512
rect 5040 26472 5264 26500
rect 5040 26460 5046 26472
rect 5258 26460 5264 26472
rect 5316 26500 5322 26512
rect 9490 26500 9496 26512
rect 5316 26472 9496 26500
rect 5316 26460 5322 26472
rect 9490 26460 9496 26472
rect 9548 26460 9554 26512
rect 11698 26460 11704 26512
rect 11756 26460 11762 26512
rect 12069 26503 12127 26509
rect 12069 26469 12081 26503
rect 12115 26500 12127 26503
rect 12544 26500 12572 26540
rect 12710 26528 12716 26540
rect 12768 26528 12774 26580
rect 15102 26528 15108 26580
rect 15160 26528 15166 26580
rect 15378 26528 15384 26580
rect 15436 26568 15442 26580
rect 15933 26571 15991 26577
rect 15933 26568 15945 26571
rect 15436 26540 15945 26568
rect 15436 26528 15442 26540
rect 15933 26537 15945 26540
rect 15979 26537 15991 26571
rect 15933 26531 15991 26537
rect 16482 26528 16488 26580
rect 16540 26568 16546 26580
rect 16540 26540 17632 26568
rect 16540 26528 16546 26540
rect 17126 26500 17132 26512
rect 12115 26472 12572 26500
rect 17052 26472 17132 26500
rect 12115 26469 12127 26472
rect 12069 26463 12127 26469
rect 11330 26392 11336 26444
rect 11388 26392 11394 26444
rect 15657 26435 15715 26441
rect 15657 26432 15669 26435
rect 14936 26404 15669 26432
rect 1302 26324 1308 26376
rect 1360 26364 1366 26376
rect 1489 26367 1547 26373
rect 1489 26364 1501 26367
rect 1360 26336 1501 26364
rect 1360 26324 1366 26336
rect 1489 26333 1501 26336
rect 1535 26364 1547 26367
rect 1949 26367 2007 26373
rect 1949 26364 1961 26367
rect 1535 26336 1961 26364
rect 1535 26333 1547 26336
rect 1489 26327 1547 26333
rect 1949 26333 1961 26336
rect 1995 26333 2007 26367
rect 1949 26327 2007 26333
rect 3513 26367 3571 26373
rect 3513 26333 3525 26367
rect 3559 26364 3571 26367
rect 3878 26364 3884 26376
rect 3559 26336 3884 26364
rect 3559 26333 3571 26336
rect 3513 26327 3571 26333
rect 3878 26324 3884 26336
rect 3936 26324 3942 26376
rect 5537 26367 5595 26373
rect 5537 26333 5549 26367
rect 5583 26364 5595 26367
rect 5718 26364 5724 26376
rect 5583 26336 5724 26364
rect 5583 26333 5595 26336
rect 5537 26327 5595 26333
rect 5718 26324 5724 26336
rect 5776 26324 5782 26376
rect 11514 26324 11520 26376
rect 11572 26324 11578 26376
rect 13354 26324 13360 26376
rect 13412 26364 13418 26376
rect 13449 26367 13507 26373
rect 13449 26364 13461 26367
rect 13412 26336 13461 26364
rect 13412 26324 13418 26336
rect 13449 26333 13461 26336
rect 13495 26364 13507 26367
rect 13722 26364 13728 26376
rect 13495 26336 13728 26364
rect 13495 26333 13507 26336
rect 13449 26327 13507 26333
rect 13722 26324 13728 26336
rect 13780 26324 13786 26376
rect 1673 26299 1731 26305
rect 1673 26265 1685 26299
rect 1719 26296 1731 26299
rect 1854 26296 1860 26308
rect 1719 26268 1860 26296
rect 1719 26265 1731 26268
rect 1673 26259 1731 26265
rect 1854 26256 1860 26268
rect 1912 26256 1918 26308
rect 3694 26256 3700 26308
rect 3752 26296 3758 26308
rect 3789 26299 3847 26305
rect 3789 26296 3801 26299
rect 3752 26268 3801 26296
rect 3752 26256 3758 26268
rect 3789 26265 3801 26268
rect 3835 26265 3847 26299
rect 3789 26259 3847 26265
rect 7469 26299 7527 26305
rect 7469 26265 7481 26299
rect 7515 26265 7527 26299
rect 7469 26259 7527 26265
rect 8496 26268 9536 26296
rect 3050 26188 3056 26240
rect 3108 26228 3114 26240
rect 3329 26231 3387 26237
rect 3329 26228 3341 26231
rect 3108 26200 3341 26228
rect 3108 26188 3114 26200
rect 3329 26197 3341 26200
rect 3375 26228 3387 26231
rect 4246 26228 4252 26240
rect 3375 26200 4252 26228
rect 3375 26197 3387 26200
rect 3329 26191 3387 26197
rect 4246 26188 4252 26200
rect 4304 26188 4310 26240
rect 6546 26188 6552 26240
rect 6604 26228 6610 26240
rect 7484 26228 7512 26259
rect 6604 26200 7512 26228
rect 6604 26188 6610 26200
rect 7742 26188 7748 26240
rect 7800 26228 7806 26240
rect 8496 26228 8524 26268
rect 7800 26200 8524 26228
rect 7800 26188 7806 26200
rect 8570 26188 8576 26240
rect 8628 26228 8634 26240
rect 9033 26231 9091 26237
rect 9033 26228 9045 26231
rect 8628 26200 9045 26228
rect 8628 26188 8634 26200
rect 9033 26197 9045 26200
rect 9079 26228 9091 26231
rect 9398 26228 9404 26240
rect 9079 26200 9404 26228
rect 9079 26197 9091 26200
rect 9033 26191 9091 26197
rect 9398 26188 9404 26200
rect 9456 26188 9462 26240
rect 9508 26228 9536 26268
rect 10594 26256 10600 26308
rect 10652 26296 10658 26308
rect 11241 26299 11299 26305
rect 11241 26296 11253 26299
rect 10652 26268 11253 26296
rect 10652 26256 10658 26268
rect 11241 26265 11253 26268
rect 11287 26265 11299 26299
rect 11241 26259 11299 26265
rect 12526 26256 12532 26308
rect 12584 26296 12590 26308
rect 13182 26299 13240 26305
rect 13182 26296 13194 26299
rect 12584 26268 13194 26296
rect 12584 26256 12590 26268
rect 13182 26265 13194 26268
rect 13228 26265 13240 26299
rect 13182 26259 13240 26265
rect 14458 26256 14464 26308
rect 14516 26296 14522 26308
rect 14936 26305 14964 26404
rect 15657 26401 15669 26404
rect 15703 26401 15715 26435
rect 15657 26395 15715 26401
rect 15473 26367 15531 26373
rect 15473 26333 15485 26367
rect 15519 26364 15531 26367
rect 15930 26364 15936 26376
rect 15519 26336 15936 26364
rect 15519 26333 15531 26336
rect 15473 26327 15531 26333
rect 15930 26324 15936 26336
rect 15988 26324 15994 26376
rect 16022 26324 16028 26376
rect 16080 26364 16086 26376
rect 16761 26367 16819 26373
rect 16761 26364 16773 26367
rect 16080 26336 16773 26364
rect 16080 26324 16086 26336
rect 16761 26333 16773 26336
rect 16807 26333 16819 26367
rect 16761 26327 16819 26333
rect 16850 26324 16856 26376
rect 16908 26324 16914 26376
rect 17052 26373 17080 26472
rect 17126 26460 17132 26472
rect 17184 26460 17190 26512
rect 17037 26367 17095 26373
rect 17037 26333 17049 26367
rect 17083 26333 17095 26367
rect 17037 26327 17095 26333
rect 17126 26324 17132 26376
rect 17184 26324 17190 26376
rect 17292 26373 17320 26540
rect 17402 26460 17408 26512
rect 17460 26460 17466 26512
rect 17604 26500 17632 26540
rect 17678 26528 17684 26580
rect 17736 26528 17742 26580
rect 17865 26571 17923 26577
rect 17865 26537 17877 26571
rect 17911 26568 17923 26571
rect 20254 26568 20260 26580
rect 17911 26540 20260 26568
rect 17911 26537 17923 26540
rect 17865 26531 17923 26537
rect 20254 26528 20260 26540
rect 20312 26528 20318 26580
rect 21450 26528 21456 26580
rect 21508 26528 21514 26580
rect 21818 26568 21824 26580
rect 21560 26540 21824 26568
rect 17604 26472 17715 26500
rect 17687 26432 17715 26472
rect 17770 26460 17776 26512
rect 17828 26500 17834 26512
rect 19978 26500 19984 26512
rect 17828 26472 19984 26500
rect 17828 26460 17834 26472
rect 19978 26460 19984 26472
rect 20036 26460 20042 26512
rect 21560 26500 21588 26540
rect 21818 26528 21824 26540
rect 21876 26568 21882 26580
rect 22281 26571 22339 26577
rect 22281 26568 22293 26571
rect 21876 26540 22293 26568
rect 21876 26528 21882 26540
rect 22281 26537 22293 26540
rect 22327 26537 22339 26571
rect 22281 26531 22339 26537
rect 22830 26528 22836 26580
rect 22888 26528 22894 26580
rect 22922 26528 22928 26580
rect 22980 26568 22986 26580
rect 22980 26540 23888 26568
rect 22980 26528 22986 26540
rect 22370 26500 22376 26512
rect 20272 26472 21588 26500
rect 21928 26472 22376 26500
rect 20272 26444 20300 26472
rect 17687 26404 18276 26432
rect 18248 26376 18276 26404
rect 20254 26392 20260 26444
rect 20312 26392 20318 26444
rect 21928 26441 21956 26472
rect 22370 26460 22376 26472
rect 22428 26460 22434 26512
rect 23860 26500 23888 26540
rect 24578 26528 24584 26580
rect 24636 26528 24642 26580
rect 26234 26568 26240 26580
rect 25332 26540 26240 26568
rect 25332 26500 25360 26540
rect 26234 26528 26240 26540
rect 26292 26528 26298 26580
rect 27338 26528 27344 26580
rect 27396 26528 27402 26580
rect 29365 26571 29423 26577
rect 29365 26537 29377 26571
rect 29411 26568 29423 26571
rect 33962 26568 33968 26580
rect 29411 26540 33968 26568
rect 29411 26537 29423 26540
rect 29365 26531 29423 26537
rect 33962 26528 33968 26540
rect 34020 26528 34026 26580
rect 23860 26472 25360 26500
rect 21913 26435 21971 26441
rect 21913 26401 21925 26435
rect 21959 26401 21971 26435
rect 21913 26395 21971 26401
rect 22002 26392 22008 26444
rect 22060 26392 22066 26444
rect 22738 26392 22744 26444
rect 22796 26432 22802 26444
rect 25240 26441 25268 26472
rect 25406 26460 25412 26512
rect 25464 26460 25470 26512
rect 25498 26460 25504 26512
rect 25556 26500 25562 26512
rect 25556 26472 25912 26500
rect 25556 26460 25562 26472
rect 23385 26435 23443 26441
rect 23385 26432 23397 26435
rect 22796 26404 23397 26432
rect 22796 26392 22802 26404
rect 23385 26401 23397 26404
rect 23431 26401 23443 26435
rect 23385 26395 23443 26401
rect 25225 26435 25283 26441
rect 25225 26401 25237 26435
rect 25271 26401 25283 26435
rect 25424 26432 25452 26460
rect 25225 26395 25283 26401
rect 25332 26404 25544 26432
rect 17267 26367 17325 26373
rect 17267 26333 17279 26367
rect 17313 26333 17325 26367
rect 17497 26367 17555 26373
rect 17497 26342 17509 26367
rect 17267 26327 17325 26333
rect 17420 26333 17509 26342
rect 17543 26333 17555 26367
rect 17420 26327 17555 26333
rect 17420 26314 17540 26327
rect 17586 26324 17592 26376
rect 17644 26324 17650 26376
rect 18046 26324 18052 26376
rect 18104 26324 18110 26376
rect 18230 26324 18236 26376
rect 18288 26324 18294 26376
rect 21634 26324 21640 26376
rect 21692 26364 21698 26376
rect 21821 26367 21879 26373
rect 21821 26364 21833 26367
rect 21692 26336 21833 26364
rect 21692 26324 21698 26336
rect 21821 26333 21833 26336
rect 21867 26364 21879 26367
rect 23201 26367 23259 26373
rect 21867 26362 22140 26364
rect 22204 26362 22784 26364
rect 21867 26336 22784 26362
rect 21867 26333 21879 26336
rect 22112 26334 22232 26336
rect 21821 26327 21879 26333
rect 14921 26299 14979 26305
rect 14921 26296 14933 26299
rect 14516 26268 14933 26296
rect 14516 26256 14522 26268
rect 14921 26265 14933 26268
rect 14967 26265 14979 26299
rect 14921 26259 14979 26265
rect 15010 26256 15016 26308
rect 15068 26296 15074 26308
rect 15565 26299 15623 26305
rect 15565 26296 15577 26299
rect 15068 26268 15577 26296
rect 15068 26256 15074 26268
rect 15565 26265 15577 26268
rect 15611 26265 15623 26299
rect 15565 26259 15623 26265
rect 15838 26256 15844 26308
rect 15896 26296 15902 26308
rect 17420 26296 17448 26314
rect 15896 26268 17448 26296
rect 17880 26268 18092 26296
rect 15896 26256 15902 26268
rect 10410 26228 10416 26240
rect 9508 26200 10416 26228
rect 10410 26188 10416 26200
rect 10468 26188 10474 26240
rect 13078 26188 13084 26240
rect 13136 26228 13142 26240
rect 13630 26228 13636 26240
rect 13136 26200 13636 26228
rect 13136 26188 13142 26200
rect 13630 26188 13636 26200
rect 13688 26188 13694 26240
rect 14090 26188 14096 26240
rect 14148 26228 14154 26240
rect 15102 26228 15108 26240
rect 14148 26200 15108 26228
rect 14148 26188 14154 26200
rect 15102 26188 15108 26200
rect 15160 26188 15166 26240
rect 16390 26188 16396 26240
rect 16448 26228 16454 26240
rect 17880 26228 17908 26268
rect 16448 26200 17908 26228
rect 18064 26228 18092 26268
rect 18138 26256 18144 26308
rect 18196 26296 18202 26308
rect 22756 26296 22784 26336
rect 23201 26333 23213 26367
rect 23247 26364 23259 26367
rect 23658 26364 23664 26376
rect 23247 26336 23664 26364
rect 23247 26333 23259 26336
rect 23201 26327 23259 26333
rect 23658 26324 23664 26336
rect 23716 26324 23722 26376
rect 24949 26367 25007 26373
rect 24949 26333 24961 26367
rect 24995 26364 25007 26367
rect 25332 26364 25360 26404
rect 25516 26373 25544 26404
rect 24995 26336 25360 26364
rect 25409 26367 25467 26373
rect 24995 26333 25007 26336
rect 24949 26327 25007 26333
rect 25409 26333 25421 26367
rect 25455 26333 25467 26367
rect 25409 26327 25467 26333
rect 25502 26367 25560 26373
rect 25502 26333 25514 26367
rect 25548 26333 25560 26367
rect 25502 26327 25560 26333
rect 23293 26299 23351 26305
rect 23293 26296 23305 26299
rect 18196 26268 22692 26296
rect 22756 26268 23305 26296
rect 18196 26256 18202 26268
rect 21542 26228 21548 26240
rect 18064 26200 21548 26228
rect 16448 26188 16454 26200
rect 21542 26188 21548 26200
rect 21600 26188 21606 26240
rect 21726 26188 21732 26240
rect 21784 26228 21790 26240
rect 22094 26228 22100 26240
rect 21784 26200 22100 26228
rect 21784 26188 21790 26200
rect 22094 26188 22100 26200
rect 22152 26188 22158 26240
rect 22664 26228 22692 26268
rect 23293 26265 23305 26268
rect 23339 26296 23351 26299
rect 23474 26296 23480 26308
rect 23339 26268 23480 26296
rect 23339 26265 23351 26268
rect 23293 26259 23351 26265
rect 23474 26256 23480 26268
rect 23532 26256 23538 26308
rect 23842 26256 23848 26308
rect 23900 26296 23906 26308
rect 25424 26296 25452 26327
rect 25590 26324 25596 26376
rect 25648 26364 25654 26376
rect 25884 26373 25912 26472
rect 25958 26460 25964 26512
rect 26016 26500 26022 26512
rect 26329 26503 26387 26509
rect 26329 26500 26341 26503
rect 26016 26472 26341 26500
rect 26016 26460 26022 26472
rect 26329 26469 26341 26472
rect 26375 26500 26387 26503
rect 27430 26500 27436 26512
rect 26375 26472 27436 26500
rect 26375 26469 26387 26472
rect 26329 26463 26387 26469
rect 27430 26460 27436 26472
rect 27488 26460 27494 26512
rect 26694 26392 26700 26444
rect 26752 26392 26758 26444
rect 27614 26392 27620 26444
rect 27672 26432 27678 26444
rect 27672 26404 28856 26432
rect 27672 26392 27678 26404
rect 25777 26367 25835 26373
rect 25777 26364 25789 26367
rect 25648 26336 25789 26364
rect 25648 26324 25654 26336
rect 25777 26333 25789 26336
rect 25823 26333 25835 26367
rect 25777 26327 25835 26333
rect 25874 26367 25932 26373
rect 25874 26333 25886 26367
rect 25920 26333 25932 26367
rect 25874 26327 25932 26333
rect 26234 26324 26240 26376
rect 26292 26324 26298 26376
rect 26510 26324 26516 26376
rect 26568 26364 26574 26376
rect 26881 26367 26939 26373
rect 26881 26364 26893 26367
rect 26568 26336 26893 26364
rect 26568 26324 26574 26336
rect 26881 26333 26893 26336
rect 26927 26333 26939 26367
rect 26881 26327 26939 26333
rect 26970 26324 26976 26376
rect 27028 26324 27034 26376
rect 28629 26367 28687 26373
rect 28629 26333 28641 26367
rect 28675 26364 28687 26367
rect 28718 26364 28724 26376
rect 28675 26336 28724 26364
rect 28675 26333 28687 26336
rect 28629 26327 28687 26333
rect 28718 26324 28724 26336
rect 28776 26324 28782 26376
rect 28828 26373 28856 26404
rect 28902 26392 28908 26444
rect 28960 26392 28966 26444
rect 28997 26435 29055 26441
rect 28997 26401 29009 26435
rect 29043 26432 29055 26435
rect 29043 26404 29684 26432
rect 29043 26401 29055 26404
rect 28997 26395 29055 26401
rect 28813 26367 28871 26373
rect 28813 26333 28825 26367
rect 28859 26333 28871 26367
rect 28813 26327 28871 26333
rect 29178 26324 29184 26376
rect 29236 26324 29242 26376
rect 29656 26373 29684 26404
rect 30098 26392 30104 26444
rect 30156 26392 30162 26444
rect 29641 26367 29699 26373
rect 29641 26333 29653 26367
rect 29687 26364 29699 26367
rect 31110 26364 31116 26376
rect 29687 26336 31116 26364
rect 29687 26333 29699 26336
rect 29641 26327 29699 26333
rect 31110 26324 31116 26336
rect 31168 26324 31174 26376
rect 31846 26324 31852 26376
rect 31904 26364 31910 26376
rect 33965 26367 34023 26373
rect 33965 26364 33977 26367
rect 31904 26336 33977 26364
rect 31904 26324 31910 26336
rect 33965 26333 33977 26336
rect 34011 26333 34023 26367
rect 33965 26327 34023 26333
rect 34238 26324 34244 26376
rect 34296 26324 34302 26376
rect 23900 26268 25452 26296
rect 25685 26299 25743 26305
rect 23900 26256 23906 26268
rect 25685 26265 25697 26299
rect 25731 26296 25743 26299
rect 25958 26296 25964 26308
rect 25731 26268 25964 26296
rect 25731 26265 25743 26268
rect 25685 26259 25743 26265
rect 25958 26256 25964 26268
rect 26016 26256 26022 26308
rect 30368 26299 30426 26305
rect 30368 26265 30380 26299
rect 30414 26296 30426 26299
rect 30466 26296 30472 26308
rect 30414 26268 30472 26296
rect 30414 26265 30426 26268
rect 30368 26259 30426 26265
rect 30466 26256 30472 26268
rect 30524 26256 30530 26308
rect 34149 26299 34207 26305
rect 34149 26265 34161 26299
rect 34195 26296 34207 26299
rect 34514 26296 34520 26308
rect 34195 26268 34520 26296
rect 34195 26265 34207 26268
rect 34149 26259 34207 26265
rect 34514 26256 34520 26268
rect 34572 26296 34578 26308
rect 34974 26296 34980 26308
rect 34572 26268 34980 26296
rect 34572 26256 34578 26268
rect 34974 26256 34980 26268
rect 35032 26256 35038 26308
rect 23750 26228 23756 26240
rect 22664 26200 23756 26228
rect 23750 26188 23756 26200
rect 23808 26188 23814 26240
rect 25041 26231 25099 26237
rect 25041 26197 25053 26231
rect 25087 26228 25099 26231
rect 25314 26228 25320 26240
rect 25087 26200 25320 26228
rect 25087 26197 25099 26200
rect 25041 26191 25099 26197
rect 25314 26188 25320 26200
rect 25372 26188 25378 26240
rect 26050 26188 26056 26240
rect 26108 26188 26114 26240
rect 31478 26188 31484 26240
rect 31536 26188 31542 26240
rect 33778 26188 33784 26240
rect 33836 26188 33842 26240
rect 1104 26138 35328 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35328 26138
rect 1104 26064 35328 26086
rect 4525 26027 4583 26033
rect 4525 25993 4537 26027
rect 4571 26024 4583 26027
rect 4706 26024 4712 26036
rect 4571 25996 4712 26024
rect 4571 25993 4583 25996
rect 4525 25987 4583 25993
rect 4706 25984 4712 25996
rect 4764 25984 4770 26036
rect 5445 26027 5503 26033
rect 5445 25993 5457 26027
rect 5491 26024 5503 26027
rect 5491 25996 10180 26024
rect 5491 25993 5503 25996
rect 5445 25987 5503 25993
rect 3973 25959 4031 25965
rect 3973 25925 3985 25959
rect 4019 25956 4031 25959
rect 4062 25956 4068 25968
rect 4019 25928 4068 25956
rect 4019 25925 4031 25928
rect 3973 25919 4031 25925
rect 4062 25916 4068 25928
rect 4120 25956 4126 25968
rect 4120 25928 4936 25956
rect 4120 25916 4126 25928
rect 4798 25848 4804 25900
rect 4856 25848 4862 25900
rect 4908 25897 4936 25928
rect 5534 25916 5540 25968
rect 5592 25956 5598 25968
rect 8021 25959 8079 25965
rect 8021 25956 8033 25959
rect 5592 25928 8033 25956
rect 5592 25916 5598 25928
rect 8021 25925 8033 25928
rect 8067 25956 8079 25959
rect 9217 25959 9275 25965
rect 8067 25928 8708 25956
rect 8067 25925 8079 25928
rect 8021 25919 8079 25925
rect 4894 25891 4952 25897
rect 4894 25857 4906 25891
rect 4940 25857 4952 25891
rect 4894 25851 4952 25857
rect 5077 25891 5135 25897
rect 5077 25857 5089 25891
rect 5123 25857 5135 25891
rect 5077 25851 5135 25857
rect 4065 25823 4123 25829
rect 4065 25789 4077 25823
rect 4111 25789 4123 25823
rect 4065 25783 4123 25789
rect 4157 25823 4215 25829
rect 4157 25789 4169 25823
rect 4203 25820 4215 25823
rect 4706 25820 4712 25832
rect 4203 25792 4712 25820
rect 4203 25789 4215 25792
rect 4157 25783 4215 25789
rect 4080 25752 4108 25783
rect 4706 25780 4712 25792
rect 4764 25780 4770 25832
rect 5092 25820 5120 25851
rect 5166 25848 5172 25900
rect 5224 25848 5230 25900
rect 5307 25891 5365 25897
rect 5307 25857 5319 25891
rect 5353 25888 5365 25891
rect 5442 25888 5448 25900
rect 5353 25860 5448 25888
rect 5353 25857 5365 25860
rect 5307 25851 5365 25857
rect 5442 25848 5448 25860
rect 5500 25848 5506 25900
rect 5721 25891 5779 25897
rect 5721 25857 5733 25891
rect 5767 25888 5779 25891
rect 6825 25891 6883 25897
rect 5767 25860 5948 25888
rect 5767 25857 5779 25860
rect 5721 25851 5779 25857
rect 5810 25820 5816 25832
rect 5092 25792 5816 25820
rect 4246 25752 4252 25764
rect 4080 25724 4252 25752
rect 4246 25712 4252 25724
rect 4304 25752 4310 25764
rect 5442 25752 5448 25764
rect 4304 25724 5448 25752
rect 4304 25712 4310 25724
rect 5442 25712 5448 25724
rect 5500 25712 5506 25764
rect 3602 25644 3608 25696
rect 3660 25644 3666 25696
rect 5537 25687 5595 25693
rect 5537 25653 5549 25687
rect 5583 25684 5595 25687
rect 5626 25684 5632 25696
rect 5583 25656 5632 25684
rect 5583 25653 5595 25656
rect 5537 25647 5595 25653
rect 5626 25644 5632 25656
rect 5684 25644 5690 25696
rect 5736 25684 5764 25792
rect 5810 25780 5816 25792
rect 5868 25780 5874 25832
rect 5920 25761 5948 25860
rect 6825 25857 6837 25891
rect 6871 25888 6883 25891
rect 7282 25888 7288 25900
rect 6871 25860 7288 25888
rect 6871 25857 6883 25860
rect 6825 25851 6883 25857
rect 7282 25848 7288 25860
rect 7340 25848 7346 25900
rect 7929 25891 7987 25897
rect 7929 25857 7941 25891
rect 7975 25888 7987 25891
rect 8202 25888 8208 25900
rect 7975 25860 8208 25888
rect 7975 25857 7987 25860
rect 7929 25851 7987 25857
rect 8202 25848 8208 25860
rect 8260 25848 8266 25900
rect 8481 25891 8539 25897
rect 8481 25857 8493 25891
rect 8527 25888 8539 25891
rect 8570 25888 8576 25900
rect 8527 25860 8576 25888
rect 8527 25857 8539 25860
rect 8481 25851 8539 25857
rect 8570 25848 8576 25860
rect 8628 25848 8634 25900
rect 8680 25888 8708 25928
rect 9217 25925 9229 25959
rect 9263 25956 9275 25959
rect 9674 25956 9680 25968
rect 9263 25928 9680 25956
rect 9263 25925 9275 25928
rect 9217 25919 9275 25925
rect 9674 25916 9680 25928
rect 9732 25956 9738 25968
rect 10152 25956 10180 25996
rect 10594 25984 10600 26036
rect 10652 25984 10658 26036
rect 12526 25984 12532 26036
rect 12584 25984 12590 26036
rect 12710 25984 12716 26036
rect 12768 26024 12774 26036
rect 12989 26027 13047 26033
rect 12989 26024 13001 26027
rect 12768 25996 13001 26024
rect 12768 25984 12774 25996
rect 12989 25993 13001 25996
rect 13035 25993 13047 26027
rect 12989 25987 13047 25993
rect 13262 25984 13268 26036
rect 13320 26024 13326 26036
rect 13357 26027 13415 26033
rect 13357 26024 13369 26027
rect 13320 25996 13369 26024
rect 13320 25984 13326 25996
rect 13357 25993 13369 25996
rect 13403 25993 13415 26027
rect 13357 25987 13415 25993
rect 15378 25984 15384 26036
rect 15436 26024 15442 26036
rect 15654 26024 15660 26036
rect 15436 25996 15660 26024
rect 15436 25984 15442 25996
rect 15654 25984 15660 25996
rect 15712 26024 15718 26036
rect 16117 26027 16175 26033
rect 16117 26024 16129 26027
rect 15712 25996 16129 26024
rect 15712 25984 15718 25996
rect 16117 25993 16129 25996
rect 16163 25993 16175 26027
rect 16117 25987 16175 25993
rect 16390 25984 16396 26036
rect 16448 25984 16454 26036
rect 16669 26027 16727 26033
rect 16669 25993 16681 26027
rect 16715 26024 16727 26027
rect 16850 26024 16856 26036
rect 16715 25996 16856 26024
rect 16715 25993 16727 25996
rect 16669 25987 16727 25993
rect 16850 25984 16856 25996
rect 16908 25984 16914 26036
rect 18785 26027 18843 26033
rect 18785 25993 18797 26027
rect 18831 26024 18843 26027
rect 20070 26024 20076 26036
rect 18831 25996 20076 26024
rect 18831 25993 18843 25996
rect 18785 25987 18843 25993
rect 20070 25984 20076 25996
rect 20128 25984 20134 26036
rect 20162 25984 20168 26036
rect 20220 26024 20226 26036
rect 20257 26027 20315 26033
rect 20257 26024 20269 26027
rect 20220 25996 20269 26024
rect 20220 25984 20226 25996
rect 20257 25993 20269 25996
rect 20303 25993 20315 26027
rect 20257 25987 20315 25993
rect 20438 25984 20444 26036
rect 20496 26024 20502 26036
rect 22738 26024 22744 26036
rect 20496 25996 22744 26024
rect 20496 25984 20502 25996
rect 22738 25984 22744 25996
rect 22796 25984 22802 26036
rect 23198 25984 23204 26036
rect 23256 26024 23262 26036
rect 23256 25996 25452 26024
rect 23256 25984 23262 25996
rect 11330 25956 11336 25968
rect 9732 25928 10088 25956
rect 10152 25928 11336 25956
rect 9732 25916 9738 25928
rect 9309 25891 9367 25897
rect 9309 25888 9321 25891
rect 8680 25860 9321 25888
rect 9309 25857 9321 25860
rect 9355 25857 9367 25891
rect 9309 25851 9367 25857
rect 9490 25848 9496 25900
rect 9548 25888 9554 25900
rect 10060 25897 10088 25928
rect 11330 25916 11336 25928
rect 11388 25916 11394 25968
rect 12894 25916 12900 25968
rect 12952 25916 12958 25968
rect 14826 25956 14832 25968
rect 14108 25928 14832 25956
rect 9953 25891 10011 25897
rect 9953 25888 9965 25891
rect 9548 25860 9965 25888
rect 9548 25848 9554 25860
rect 9953 25857 9965 25860
rect 9999 25857 10011 25891
rect 9953 25851 10011 25857
rect 10046 25891 10104 25897
rect 10046 25857 10058 25891
rect 10092 25857 10104 25891
rect 10046 25851 10104 25857
rect 10134 25848 10140 25900
rect 10192 25888 10198 25900
rect 10229 25891 10287 25897
rect 10229 25888 10241 25891
rect 10192 25860 10241 25888
rect 10192 25848 10198 25860
rect 10229 25857 10241 25860
rect 10275 25857 10287 25891
rect 10229 25851 10287 25857
rect 6546 25780 6552 25832
rect 6604 25780 6610 25832
rect 8113 25823 8171 25829
rect 8113 25789 8125 25823
rect 8159 25820 8171 25823
rect 8294 25820 8300 25832
rect 8159 25792 8300 25820
rect 8159 25789 8171 25792
rect 8113 25783 8171 25789
rect 8294 25780 8300 25792
rect 8352 25780 8358 25832
rect 9401 25823 9459 25829
rect 9401 25789 9413 25823
rect 9447 25820 9459 25823
rect 9766 25820 9772 25832
rect 9447 25792 9772 25820
rect 9447 25789 9459 25792
rect 9401 25783 9459 25789
rect 9766 25780 9772 25792
rect 9824 25780 9830 25832
rect 10244 25820 10272 25851
rect 10318 25848 10324 25900
rect 10376 25848 10382 25900
rect 10410 25848 10416 25900
rect 10468 25897 10474 25900
rect 10468 25891 10517 25897
rect 10468 25857 10471 25891
rect 10505 25888 10517 25891
rect 10505 25860 11008 25888
rect 10505 25857 10517 25860
rect 10468 25851 10517 25857
rect 10468 25848 10474 25851
rect 10980 25832 11008 25860
rect 13722 25848 13728 25900
rect 13780 25888 13786 25900
rect 14108 25897 14136 25928
rect 14826 25916 14832 25928
rect 14884 25956 14890 25968
rect 16482 25956 16488 25968
rect 14884 25928 16488 25956
rect 14884 25916 14890 25928
rect 16482 25916 16488 25928
rect 16540 25916 16546 25968
rect 19889 25959 19947 25965
rect 17052 25928 18460 25956
rect 14093 25891 14151 25897
rect 14093 25888 14105 25891
rect 13780 25860 14105 25888
rect 13780 25848 13786 25860
rect 14093 25857 14105 25860
rect 14139 25857 14151 25891
rect 14093 25851 14151 25857
rect 14360 25891 14418 25897
rect 14360 25857 14372 25891
rect 14406 25888 14418 25891
rect 14642 25888 14648 25900
rect 14406 25860 14648 25888
rect 14406 25857 14418 25860
rect 14360 25851 14418 25857
rect 14642 25848 14648 25860
rect 14700 25848 14706 25900
rect 15841 25891 15899 25897
rect 15841 25857 15853 25891
rect 15887 25888 15899 25891
rect 16390 25888 16396 25900
rect 15887 25860 16396 25888
rect 15887 25857 15899 25860
rect 15841 25851 15899 25857
rect 16390 25848 16396 25860
rect 16448 25848 16454 25900
rect 10689 25823 10747 25829
rect 10689 25820 10701 25823
rect 10244 25792 10701 25820
rect 10689 25789 10701 25792
rect 10735 25789 10747 25823
rect 10689 25783 10747 25789
rect 10962 25780 10968 25832
rect 11020 25780 11026 25832
rect 13173 25823 13231 25829
rect 13173 25789 13185 25823
rect 13219 25820 13231 25823
rect 13262 25820 13268 25832
rect 13219 25792 13268 25820
rect 13219 25789 13231 25792
rect 13173 25783 13231 25789
rect 13262 25780 13268 25792
rect 13320 25780 13326 25832
rect 15102 25780 15108 25832
rect 15160 25820 15166 25832
rect 17052 25820 17080 25928
rect 17218 25848 17224 25900
rect 17276 25888 17282 25900
rect 17782 25891 17840 25897
rect 17782 25888 17794 25891
rect 17276 25860 17794 25888
rect 17276 25848 17282 25860
rect 17782 25857 17794 25860
rect 17828 25857 17840 25891
rect 17782 25851 17840 25857
rect 15160 25792 17080 25820
rect 15160 25780 15166 25792
rect 18046 25780 18052 25832
rect 18104 25780 18110 25832
rect 5905 25755 5963 25761
rect 5905 25721 5917 25755
rect 5951 25752 5963 25755
rect 11698 25752 11704 25764
rect 5951 25724 11704 25752
rect 5951 25721 5963 25724
rect 5905 25715 5963 25721
rect 11698 25712 11704 25724
rect 11756 25712 11762 25764
rect 6089 25687 6147 25693
rect 6089 25684 6101 25687
rect 5736 25656 6101 25684
rect 6089 25653 6101 25656
rect 6135 25684 6147 25687
rect 6178 25684 6184 25696
rect 6135 25656 6184 25684
rect 6135 25653 6147 25656
rect 6089 25647 6147 25653
rect 6178 25644 6184 25656
rect 6236 25644 6242 25696
rect 7558 25644 7564 25696
rect 7616 25644 7622 25696
rect 7650 25644 7656 25696
rect 7708 25684 7714 25696
rect 8754 25684 8760 25696
rect 7708 25656 8760 25684
rect 7708 25644 7714 25656
rect 8754 25644 8760 25656
rect 8812 25644 8818 25696
rect 8846 25644 8852 25696
rect 8904 25644 8910 25696
rect 9122 25644 9128 25696
rect 9180 25684 9186 25696
rect 9769 25687 9827 25693
rect 9769 25684 9781 25687
rect 9180 25656 9781 25684
rect 9180 25644 9186 25656
rect 9769 25653 9781 25656
rect 9815 25684 9827 25687
rect 9858 25684 9864 25696
rect 9815 25656 9864 25684
rect 9815 25653 9827 25656
rect 9769 25647 9827 25653
rect 9858 25644 9864 25656
rect 9916 25684 9922 25696
rect 10502 25684 10508 25696
rect 9916 25656 10508 25684
rect 9916 25644 9922 25656
rect 10502 25644 10508 25656
rect 10560 25644 10566 25696
rect 15473 25687 15531 25693
rect 15473 25653 15485 25687
rect 15519 25684 15531 25687
rect 15562 25684 15568 25696
rect 15519 25656 15568 25684
rect 15519 25653 15531 25656
rect 15473 25647 15531 25653
rect 15562 25644 15568 25656
rect 15620 25644 15626 25696
rect 16025 25687 16083 25693
rect 16025 25653 16037 25687
rect 16071 25684 16083 25687
rect 16114 25684 16120 25696
rect 16071 25656 16120 25684
rect 16071 25653 16083 25656
rect 16025 25647 16083 25653
rect 16114 25644 16120 25656
rect 16172 25644 16178 25696
rect 18322 25644 18328 25696
rect 18380 25644 18386 25696
rect 18432 25684 18460 25928
rect 19076 25928 19748 25956
rect 19076 25900 19104 25928
rect 18693 25891 18751 25897
rect 18693 25857 18705 25891
rect 18739 25888 18751 25891
rect 19058 25888 19064 25900
rect 18739 25860 19064 25888
rect 18739 25857 18751 25860
rect 18693 25851 18751 25857
rect 19058 25848 19064 25860
rect 19116 25848 19122 25900
rect 19610 25848 19616 25900
rect 19668 25848 19674 25900
rect 19720 25897 19748 25928
rect 19889 25925 19901 25959
rect 19935 25956 19947 25959
rect 20622 25956 20628 25968
rect 19935 25928 20628 25956
rect 19935 25925 19947 25928
rect 19889 25919 19947 25925
rect 20622 25916 20628 25928
rect 20680 25916 20686 25968
rect 21836 25928 22977 25956
rect 19706 25891 19764 25897
rect 19706 25857 19718 25891
rect 19752 25857 19764 25891
rect 19706 25851 19764 25857
rect 19978 25848 19984 25900
rect 20036 25848 20042 25900
rect 20119 25891 20177 25897
rect 20119 25857 20131 25891
rect 20165 25888 20177 25891
rect 21836 25888 21864 25928
rect 20165 25860 21864 25888
rect 20165 25857 20177 25860
rect 20119 25851 20177 25857
rect 21910 25848 21916 25900
rect 21968 25848 21974 25900
rect 22949 25888 22977 25928
rect 23014 25916 23020 25968
rect 23072 25956 23078 25968
rect 23072 25928 25351 25956
rect 23072 25916 23078 25928
rect 23566 25888 23572 25900
rect 22949 25860 23572 25888
rect 23566 25848 23572 25860
rect 23624 25848 23630 25900
rect 24118 25848 24124 25900
rect 24176 25888 24182 25900
rect 24305 25891 24363 25897
rect 24305 25888 24317 25891
rect 24176 25860 24317 25888
rect 24176 25848 24182 25860
rect 24305 25857 24317 25860
rect 24351 25857 24363 25891
rect 24305 25851 24363 25857
rect 24572 25891 24630 25897
rect 24572 25857 24584 25891
rect 24618 25888 24630 25891
rect 24854 25888 24860 25900
rect 24618 25860 24860 25888
rect 24618 25857 24630 25860
rect 24572 25851 24630 25857
rect 24854 25848 24860 25860
rect 24912 25848 24918 25900
rect 18874 25780 18880 25832
rect 18932 25820 18938 25832
rect 19153 25823 19211 25829
rect 19153 25820 19165 25823
rect 18932 25792 19165 25820
rect 18932 25780 18938 25792
rect 19153 25789 19165 25792
rect 19199 25789 19211 25823
rect 21726 25820 21732 25832
rect 19153 25783 19211 25789
rect 19352 25792 21732 25820
rect 19352 25684 19380 25792
rect 21726 25780 21732 25792
rect 21784 25780 21790 25832
rect 25323 25820 25351 25928
rect 25424 25888 25452 25996
rect 26510 25984 26516 26036
rect 26568 25984 26574 26036
rect 28166 25984 28172 26036
rect 28224 26024 28230 26036
rect 29825 26027 29883 26033
rect 29825 26024 29837 26027
rect 28224 25996 29837 26024
rect 28224 25984 28230 25996
rect 29825 25993 29837 25996
rect 29871 26024 29883 26027
rect 30285 26027 30343 26033
rect 29871 25996 30236 26024
rect 29871 25993 29883 25996
rect 29825 25987 29883 25993
rect 25961 25891 26019 25897
rect 25961 25888 25973 25891
rect 25424 25860 25973 25888
rect 25961 25857 25973 25860
rect 26007 25888 26019 25891
rect 27246 25888 27252 25900
rect 26007 25860 27252 25888
rect 26007 25857 26019 25860
rect 25961 25851 26019 25857
rect 27246 25848 27252 25860
rect 27304 25848 27310 25900
rect 30208 25888 30236 25996
rect 30285 25993 30297 26027
rect 30331 26024 30343 26027
rect 30466 26024 30472 26036
rect 30331 25996 30472 26024
rect 30331 25993 30343 25996
rect 30285 25987 30343 25993
rect 30466 25984 30472 25996
rect 30524 25984 30530 26036
rect 30653 26027 30711 26033
rect 30653 25993 30665 26027
rect 30699 26024 30711 26027
rect 30742 26024 30748 26036
rect 30699 25996 30748 26024
rect 30699 25993 30711 25996
rect 30653 25987 30711 25993
rect 30742 25984 30748 25996
rect 30800 26024 30806 26036
rect 31478 26024 31484 26036
rect 30800 25996 31484 26024
rect 30800 25984 30806 25996
rect 31478 25984 31484 25996
rect 31536 25984 31542 26036
rect 33594 25984 33600 26036
rect 33652 26024 33658 26036
rect 33652 25996 33916 26024
rect 33652 25984 33658 25996
rect 33505 25959 33563 25965
rect 33505 25925 33517 25959
rect 33551 25956 33563 25959
rect 33778 25956 33784 25968
rect 33551 25928 33784 25956
rect 33551 25925 33563 25928
rect 33505 25919 33563 25925
rect 33778 25916 33784 25928
rect 33836 25916 33842 25968
rect 33888 25956 33916 25996
rect 34974 25984 34980 26036
rect 35032 25984 35038 26036
rect 33962 25956 33968 25968
rect 33888 25928 33968 25956
rect 33962 25916 33968 25928
rect 34020 25916 34026 25968
rect 30208 25860 30880 25888
rect 30098 25820 30104 25832
rect 25323 25792 30104 25820
rect 30098 25780 30104 25792
rect 30156 25780 30162 25832
rect 30650 25780 30656 25832
rect 30708 25820 30714 25832
rect 30852 25829 30880 25860
rect 30745 25823 30803 25829
rect 30745 25820 30757 25823
rect 30708 25792 30757 25820
rect 30708 25780 30714 25792
rect 30745 25789 30757 25792
rect 30791 25789 30803 25823
rect 30745 25783 30803 25789
rect 30837 25823 30895 25829
rect 30837 25789 30849 25823
rect 30883 25789 30895 25823
rect 30837 25783 30895 25789
rect 32766 25780 32772 25832
rect 32824 25820 32830 25832
rect 33229 25823 33287 25829
rect 33229 25820 33241 25823
rect 32824 25792 33241 25820
rect 32824 25780 32830 25792
rect 33229 25789 33241 25792
rect 33275 25789 33287 25823
rect 33229 25783 33287 25789
rect 25314 25712 25320 25764
rect 25372 25752 25378 25764
rect 25777 25755 25835 25761
rect 25777 25752 25789 25755
rect 25372 25724 25789 25752
rect 25372 25712 25378 25724
rect 25777 25721 25789 25724
rect 25823 25721 25835 25755
rect 25777 25715 25835 25721
rect 28994 25712 29000 25764
rect 29052 25752 29058 25764
rect 29052 25724 30144 25752
rect 29052 25712 29058 25724
rect 18432 25656 19380 25684
rect 20441 25687 20499 25693
rect 20441 25653 20453 25687
rect 20487 25684 20499 25687
rect 20622 25684 20628 25696
rect 20487 25656 20628 25684
rect 20487 25653 20499 25656
rect 20441 25647 20499 25653
rect 20622 25644 20628 25656
rect 20680 25644 20686 25696
rect 22094 25644 22100 25696
rect 22152 25684 22158 25696
rect 22281 25687 22339 25693
rect 22281 25684 22293 25687
rect 22152 25656 22293 25684
rect 22152 25644 22158 25656
rect 22281 25653 22293 25656
rect 22327 25653 22339 25687
rect 22281 25647 22339 25653
rect 22462 25644 22468 25696
rect 22520 25644 22526 25696
rect 25222 25644 25228 25696
rect 25280 25684 25286 25696
rect 25590 25684 25596 25696
rect 25280 25656 25596 25684
rect 25280 25644 25286 25656
rect 25590 25644 25596 25656
rect 25648 25684 25654 25696
rect 30116 25693 30144 25724
rect 25685 25687 25743 25693
rect 25685 25684 25697 25687
rect 25648 25656 25697 25684
rect 25648 25644 25654 25656
rect 25685 25653 25697 25656
rect 25731 25653 25743 25687
rect 25685 25647 25743 25653
rect 30101 25687 30159 25693
rect 30101 25653 30113 25687
rect 30147 25684 30159 25687
rect 31018 25684 31024 25696
rect 30147 25656 31024 25684
rect 30147 25653 30159 25656
rect 30101 25647 30159 25653
rect 31018 25644 31024 25656
rect 31076 25644 31082 25696
rect 1104 25594 35328 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 35328 25594
rect 1104 25520 35328 25542
rect 5166 25440 5172 25492
rect 5224 25480 5230 25492
rect 5261 25483 5319 25489
rect 5261 25480 5273 25483
rect 5224 25452 5273 25480
rect 5224 25440 5230 25452
rect 5261 25449 5273 25452
rect 5307 25449 5319 25483
rect 5261 25443 5319 25449
rect 8202 25440 8208 25492
rect 8260 25440 8266 25492
rect 9490 25440 9496 25492
rect 9548 25440 9554 25492
rect 12710 25480 12716 25492
rect 9646 25452 12716 25480
rect 3418 25304 3424 25356
rect 3476 25344 3482 25356
rect 3881 25347 3939 25353
rect 3881 25344 3893 25347
rect 3476 25316 3893 25344
rect 3476 25304 3482 25316
rect 3881 25313 3893 25316
rect 3927 25313 3939 25347
rect 3881 25307 3939 25313
rect 3896 25276 3924 25307
rect 5353 25279 5411 25285
rect 5353 25276 5365 25279
rect 3896 25248 5365 25276
rect 5353 25245 5365 25248
rect 5399 25276 5411 25279
rect 6825 25279 6883 25285
rect 6825 25276 6837 25279
rect 5399 25248 6837 25276
rect 5399 25245 5411 25248
rect 5353 25239 5411 25245
rect 6825 25245 6837 25248
rect 6871 25245 6883 25279
rect 6825 25239 6883 25245
rect 7092 25279 7150 25285
rect 7092 25245 7104 25279
rect 7138 25276 7150 25279
rect 7558 25276 7564 25288
rect 7138 25248 7564 25276
rect 7138 25245 7150 25248
rect 7092 25239 7150 25245
rect 7558 25236 7564 25248
rect 7616 25236 7622 25288
rect 8220 25276 8248 25440
rect 9398 25372 9404 25424
rect 9456 25412 9462 25424
rect 9646 25412 9674 25452
rect 12710 25440 12716 25452
rect 12768 25440 12774 25492
rect 12986 25440 12992 25492
rect 13044 25440 13050 25492
rect 14642 25440 14648 25492
rect 14700 25440 14706 25492
rect 16022 25440 16028 25492
rect 16080 25440 16086 25492
rect 16298 25440 16304 25492
rect 16356 25440 16362 25492
rect 17129 25483 17187 25489
rect 17129 25449 17141 25483
rect 17175 25480 17187 25483
rect 17218 25480 17224 25492
rect 17175 25452 17224 25480
rect 17175 25449 17187 25452
rect 17129 25443 17187 25449
rect 17218 25440 17224 25452
rect 17276 25440 17282 25492
rect 18046 25480 18052 25492
rect 17696 25452 18052 25480
rect 9456 25384 9674 25412
rect 15028 25384 16160 25412
rect 9456 25372 9462 25384
rect 8754 25304 8760 25356
rect 8812 25344 8818 25356
rect 8812 25316 9352 25344
rect 8812 25304 8818 25316
rect 9324 25285 9352 25316
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 8220 25248 8953 25276
rect 8941 25245 8953 25248
rect 8987 25245 8999 25279
rect 9217 25279 9275 25285
rect 9217 25276 9229 25279
rect 8941 25239 8999 25245
rect 9048 25248 9229 25276
rect 4148 25211 4206 25217
rect 4148 25177 4160 25211
rect 4194 25208 4206 25211
rect 4522 25208 4528 25220
rect 4194 25180 4528 25208
rect 4194 25177 4206 25180
rect 4148 25171 4206 25177
rect 4522 25168 4528 25180
rect 4580 25168 4586 25220
rect 5620 25211 5678 25217
rect 5620 25177 5632 25211
rect 5666 25208 5678 25211
rect 6362 25208 6368 25220
rect 5666 25180 6368 25208
rect 5666 25177 5678 25180
rect 5620 25171 5678 25177
rect 6362 25168 6368 25180
rect 6420 25168 6426 25220
rect 9048 25208 9076 25248
rect 9217 25245 9229 25248
rect 9263 25245 9275 25279
rect 9217 25239 9275 25245
rect 9309 25279 9367 25285
rect 9309 25245 9321 25279
rect 9355 25245 9367 25279
rect 9309 25239 9367 25245
rect 9677 25279 9735 25285
rect 9677 25245 9689 25279
rect 9723 25276 9735 25279
rect 9766 25276 9772 25288
rect 9723 25248 9772 25276
rect 9723 25245 9735 25248
rect 9677 25239 9735 25245
rect 9766 25236 9772 25248
rect 9824 25276 9830 25288
rect 11609 25279 11667 25285
rect 11609 25276 11621 25279
rect 9824 25248 11621 25276
rect 9824 25236 9830 25248
rect 11609 25245 11621 25248
rect 11655 25245 11667 25279
rect 11609 25239 11667 25245
rect 11698 25236 11704 25288
rect 11756 25276 11762 25288
rect 13998 25276 14004 25288
rect 11756 25248 14004 25276
rect 11756 25236 11762 25248
rect 13998 25236 14004 25248
rect 14056 25276 14062 25288
rect 15028 25276 15056 25384
rect 15194 25304 15200 25356
rect 15252 25344 15258 25356
rect 15289 25347 15347 25353
rect 15289 25344 15301 25347
rect 15252 25316 15301 25344
rect 15252 25304 15258 25316
rect 15289 25313 15301 25316
rect 15335 25344 15347 25347
rect 16022 25344 16028 25356
rect 15335 25316 16028 25344
rect 15335 25313 15347 25316
rect 15289 25307 15347 25313
rect 16022 25304 16028 25316
rect 16080 25304 16086 25356
rect 14056 25248 15056 25276
rect 14056 25236 14062 25248
rect 15102 25236 15108 25288
rect 15160 25276 15166 25288
rect 15473 25279 15531 25285
rect 15473 25276 15485 25279
rect 15160 25248 15485 25276
rect 15160 25236 15166 25248
rect 15473 25245 15485 25248
rect 15519 25245 15531 25279
rect 15473 25239 15531 25245
rect 15562 25236 15568 25288
rect 15620 25276 15626 25288
rect 15749 25279 15807 25285
rect 15749 25276 15761 25279
rect 15620 25248 15761 25276
rect 15620 25236 15626 25248
rect 15749 25245 15761 25248
rect 15795 25245 15807 25279
rect 15749 25239 15807 25245
rect 15841 25279 15899 25285
rect 15841 25245 15853 25279
rect 15887 25245 15899 25279
rect 15841 25239 15899 25245
rect 6748 25180 9076 25208
rect 6748 25152 6776 25180
rect 9122 25168 9128 25220
rect 9180 25168 9186 25220
rect 9944 25211 10002 25217
rect 9944 25177 9956 25211
rect 9990 25208 10002 25211
rect 10134 25208 10140 25220
rect 9990 25180 10140 25208
rect 9990 25177 10002 25180
rect 9944 25171 10002 25177
rect 10134 25168 10140 25180
rect 10192 25168 10198 25220
rect 10962 25208 10968 25220
rect 10244 25180 10968 25208
rect 6730 25100 6736 25152
rect 6788 25100 6794 25152
rect 8294 25100 8300 25152
rect 8352 25140 8358 25152
rect 8573 25143 8631 25149
rect 8573 25140 8585 25143
rect 8352 25112 8585 25140
rect 8352 25100 8358 25112
rect 8573 25109 8585 25112
rect 8619 25140 8631 25143
rect 10244 25140 10272 25180
rect 10962 25168 10968 25180
rect 11020 25168 11026 25220
rect 11876 25211 11934 25217
rect 11876 25177 11888 25211
rect 11922 25208 11934 25211
rect 12158 25208 12164 25220
rect 11922 25180 12164 25208
rect 11922 25177 11934 25180
rect 11876 25171 11934 25177
rect 12158 25168 12164 25180
rect 12216 25168 12222 25220
rect 15013 25211 15071 25217
rect 15013 25177 15025 25211
rect 15059 25208 15071 25211
rect 15580 25208 15608 25236
rect 15059 25180 15608 25208
rect 15059 25177 15071 25180
rect 15013 25171 15071 25177
rect 15654 25168 15660 25220
rect 15712 25168 15718 25220
rect 8619 25112 10272 25140
rect 8619 25109 8631 25112
rect 8573 25103 8631 25109
rect 10318 25100 10324 25152
rect 10376 25140 10382 25152
rect 11057 25143 11115 25149
rect 11057 25140 11069 25143
rect 10376 25112 11069 25140
rect 10376 25100 10382 25112
rect 11057 25109 11069 25112
rect 11103 25109 11115 25143
rect 11057 25103 11115 25109
rect 14918 25100 14924 25152
rect 14976 25140 14982 25152
rect 15105 25143 15163 25149
rect 15105 25140 15117 25143
rect 14976 25112 15117 25140
rect 14976 25100 14982 25112
rect 15105 25109 15117 25112
rect 15151 25109 15163 25143
rect 15857 25140 15885 25239
rect 16132 25208 16160 25384
rect 16482 25372 16488 25424
rect 16540 25412 16546 25424
rect 17696 25412 17724 25452
rect 18046 25440 18052 25452
rect 18104 25440 18110 25492
rect 19058 25440 19064 25492
rect 19116 25440 19122 25492
rect 19150 25440 19156 25492
rect 19208 25480 19214 25492
rect 19208 25452 24808 25480
rect 19208 25440 19214 25452
rect 16540 25384 17724 25412
rect 16540 25372 16546 25384
rect 16574 25304 16580 25356
rect 16632 25304 16638 25356
rect 16669 25347 16727 25353
rect 16669 25313 16681 25347
rect 16715 25344 16727 25347
rect 16850 25344 16856 25356
rect 16715 25316 16856 25344
rect 16715 25313 16727 25316
rect 16669 25307 16727 25313
rect 16850 25304 16856 25316
rect 16908 25304 16914 25356
rect 17696 25353 17724 25384
rect 22094 25372 22100 25424
rect 22152 25412 22158 25424
rect 22373 25415 22431 25421
rect 22373 25412 22385 25415
rect 22152 25384 22385 25412
rect 22152 25372 22158 25384
rect 22373 25381 22385 25384
rect 22419 25381 22431 25415
rect 24780 25412 24808 25452
rect 24854 25440 24860 25492
rect 24912 25440 24918 25492
rect 25774 25440 25780 25492
rect 25832 25480 25838 25492
rect 25869 25483 25927 25489
rect 25869 25480 25881 25483
rect 25832 25452 25881 25480
rect 25832 25440 25838 25452
rect 25869 25449 25881 25452
rect 25915 25449 25927 25483
rect 25869 25443 25927 25449
rect 27246 25440 27252 25492
rect 27304 25480 27310 25492
rect 30650 25480 30656 25492
rect 27304 25452 29500 25480
rect 27304 25440 27310 25452
rect 29365 25415 29423 25421
rect 24780 25384 26372 25412
rect 22373 25375 22431 25381
rect 17681 25347 17739 25353
rect 17681 25313 17693 25347
rect 17727 25313 17739 25347
rect 17681 25307 17739 25313
rect 22186 25304 22192 25356
rect 22244 25344 22250 25356
rect 22462 25344 22468 25356
rect 22244 25316 22468 25344
rect 22244 25304 22250 25316
rect 22462 25304 22468 25316
rect 22520 25304 22526 25356
rect 25409 25347 25467 25353
rect 25409 25344 25421 25347
rect 24688 25316 25421 25344
rect 16758 25236 16764 25288
rect 16816 25236 16822 25288
rect 17948 25279 18006 25285
rect 17948 25245 17960 25279
rect 17994 25276 18006 25279
rect 18322 25276 18328 25288
rect 17994 25248 18328 25276
rect 17994 25245 18006 25248
rect 17948 25239 18006 25245
rect 18322 25236 18328 25248
rect 18380 25236 18386 25288
rect 18966 25236 18972 25288
rect 19024 25276 19030 25288
rect 19337 25279 19395 25285
rect 19337 25276 19349 25279
rect 19024 25248 19349 25276
rect 19024 25236 19030 25248
rect 19337 25245 19349 25248
rect 19383 25245 19395 25279
rect 20438 25276 20444 25288
rect 19337 25239 19395 25245
rect 19444 25248 20444 25276
rect 19444 25208 19472 25248
rect 20438 25236 20444 25248
rect 20496 25236 20502 25288
rect 20901 25279 20959 25285
rect 20901 25245 20913 25279
rect 20947 25276 20959 25279
rect 22278 25276 22284 25288
rect 20947 25248 22284 25276
rect 20947 25245 20959 25248
rect 20901 25239 20959 25245
rect 22278 25236 22284 25248
rect 22336 25276 22342 25288
rect 22554 25276 22560 25288
rect 22336 25248 22560 25276
rect 22336 25236 22342 25248
rect 22554 25236 22560 25248
rect 22612 25236 22618 25288
rect 16132 25180 19472 25208
rect 19604 25211 19662 25217
rect 19604 25177 19616 25211
rect 19650 25208 19662 25211
rect 19702 25208 19708 25220
rect 19650 25180 19708 25208
rect 19650 25177 19662 25180
rect 19604 25171 19662 25177
rect 19702 25168 19708 25180
rect 19760 25168 19766 25220
rect 21168 25211 21226 25217
rect 21168 25177 21180 25211
rect 21214 25208 21226 25211
rect 21818 25208 21824 25220
rect 21214 25180 21824 25208
rect 21214 25177 21226 25180
rect 21168 25171 21226 25177
rect 21818 25168 21824 25180
rect 21876 25168 21882 25220
rect 22824 25211 22882 25217
rect 22824 25177 22836 25211
rect 22870 25208 22882 25211
rect 23106 25208 23112 25220
rect 22870 25180 23112 25208
rect 22870 25177 22882 25180
rect 22824 25171 22882 25177
rect 23106 25168 23112 25180
rect 23164 25168 23170 25220
rect 23750 25168 23756 25220
rect 23808 25208 23814 25220
rect 24029 25211 24087 25217
rect 24029 25208 24041 25211
rect 23808 25180 24041 25208
rect 23808 25168 23814 25180
rect 24029 25177 24041 25180
rect 24075 25177 24087 25211
rect 24029 25171 24087 25177
rect 16298 25140 16304 25152
rect 15857 25112 16304 25140
rect 15105 25103 15163 25109
rect 16298 25100 16304 25112
rect 16356 25100 16362 25152
rect 16574 25100 16580 25152
rect 16632 25140 16638 25152
rect 17313 25143 17371 25149
rect 17313 25140 17325 25143
rect 16632 25112 17325 25140
rect 16632 25100 16638 25112
rect 17313 25109 17325 25112
rect 17359 25140 17371 25143
rect 17494 25140 17500 25152
rect 17359 25112 17500 25140
rect 17359 25109 17371 25112
rect 17313 25103 17371 25109
rect 17494 25100 17500 25112
rect 17552 25100 17558 25152
rect 19978 25100 19984 25152
rect 20036 25140 20042 25152
rect 20717 25143 20775 25149
rect 20717 25140 20729 25143
rect 20036 25112 20729 25140
rect 20036 25100 20042 25112
rect 20717 25109 20729 25112
rect 20763 25109 20775 25143
rect 20717 25103 20775 25109
rect 22278 25100 22284 25152
rect 22336 25100 22342 25152
rect 23934 25100 23940 25152
rect 23992 25100 23998 25152
rect 24578 25100 24584 25152
rect 24636 25140 24642 25152
rect 24688 25149 24716 25316
rect 25409 25313 25421 25316
rect 25455 25313 25467 25347
rect 26344 25344 26372 25384
rect 29365 25381 29377 25415
rect 29411 25381 29423 25415
rect 29365 25375 29423 25381
rect 26344 25316 26464 25344
rect 25409 25307 25467 25313
rect 24946 25236 24952 25288
rect 25004 25276 25010 25288
rect 26329 25279 26387 25285
rect 26329 25276 26341 25279
rect 25004 25248 26341 25276
rect 25004 25236 25010 25248
rect 26329 25245 26341 25248
rect 26375 25245 26387 25279
rect 26436 25276 26464 25316
rect 26436 25248 27936 25276
rect 26329 25239 26387 25245
rect 25222 25168 25228 25220
rect 25280 25168 25286 25220
rect 26596 25211 26654 25217
rect 26596 25177 26608 25211
rect 26642 25208 26654 25211
rect 26970 25208 26976 25220
rect 26642 25180 26976 25208
rect 26642 25177 26654 25180
rect 26596 25171 26654 25177
rect 26970 25168 26976 25180
rect 27028 25168 27034 25220
rect 27908 25208 27936 25248
rect 27982 25236 27988 25288
rect 28040 25236 28046 25288
rect 29380 25276 29408 25375
rect 29472 25344 29500 25452
rect 30024 25452 30656 25480
rect 30024 25353 30052 25452
rect 30650 25440 30656 25452
rect 30708 25480 30714 25492
rect 30926 25480 30932 25492
rect 30708 25452 30932 25480
rect 30708 25440 30714 25452
rect 30926 25440 30932 25452
rect 30984 25440 30990 25492
rect 31294 25412 31300 25424
rect 30300 25384 31300 25412
rect 30009 25347 30067 25353
rect 30009 25344 30021 25347
rect 29472 25316 30021 25344
rect 30009 25313 30021 25316
rect 30055 25313 30067 25347
rect 30009 25307 30067 25313
rect 30190 25304 30196 25356
rect 30248 25344 30254 25356
rect 30300 25344 30328 25384
rect 31294 25372 31300 25384
rect 31352 25372 31358 25424
rect 30558 25344 30564 25356
rect 30248 25316 30328 25344
rect 30392 25316 30564 25344
rect 30248 25304 30254 25316
rect 30392 25285 30420 25316
rect 30558 25304 30564 25316
rect 30616 25304 30622 25356
rect 29917 25279 29975 25285
rect 29917 25276 29929 25279
rect 29380 25248 29929 25276
rect 29917 25245 29929 25248
rect 29963 25245 29975 25279
rect 29917 25239 29975 25245
rect 30377 25279 30435 25285
rect 30377 25245 30389 25279
rect 30423 25245 30435 25279
rect 30377 25239 30435 25245
rect 30470 25279 30528 25285
rect 30470 25245 30482 25279
rect 30516 25245 30528 25279
rect 30470 25239 30528 25245
rect 28074 25208 28080 25220
rect 27908 25180 28080 25208
rect 28074 25168 28080 25180
rect 28132 25168 28138 25220
rect 28252 25211 28310 25217
rect 28252 25177 28264 25211
rect 28298 25208 28310 25211
rect 29932 25208 29960 25239
rect 30484 25208 30512 25239
rect 30742 25236 30748 25288
rect 30800 25236 30806 25288
rect 30883 25279 30941 25285
rect 30883 25245 30895 25279
rect 30929 25276 30941 25279
rect 31018 25276 31024 25288
rect 30929 25248 31024 25276
rect 30929 25245 30941 25248
rect 30883 25239 30941 25245
rect 31018 25236 31024 25248
rect 31076 25236 31082 25288
rect 28298 25180 29592 25208
rect 29932 25180 30512 25208
rect 30653 25211 30711 25217
rect 28298 25177 28310 25180
rect 28252 25171 28310 25177
rect 24673 25143 24731 25149
rect 24673 25140 24685 25143
rect 24636 25112 24685 25140
rect 24636 25100 24642 25112
rect 24673 25109 24685 25112
rect 24719 25109 24731 25143
rect 24673 25103 24731 25109
rect 25314 25100 25320 25152
rect 25372 25100 25378 25152
rect 25682 25100 25688 25152
rect 25740 25100 25746 25152
rect 26234 25100 26240 25152
rect 26292 25100 26298 25152
rect 27338 25100 27344 25152
rect 27396 25140 27402 25152
rect 29564 25149 29592 25180
rect 30653 25177 30665 25211
rect 30699 25208 30711 25211
rect 31113 25211 31171 25217
rect 31113 25208 31125 25211
rect 30699 25180 31125 25208
rect 30699 25177 30711 25180
rect 30653 25171 30711 25177
rect 31113 25177 31125 25180
rect 31159 25177 31171 25211
rect 31113 25171 31171 25177
rect 27709 25143 27767 25149
rect 27709 25140 27721 25143
rect 27396 25112 27721 25140
rect 27396 25100 27402 25112
rect 27709 25109 27721 25112
rect 27755 25109 27767 25143
rect 27709 25103 27767 25109
rect 29549 25143 29607 25149
rect 29549 25109 29561 25143
rect 29595 25109 29607 25143
rect 29549 25103 29607 25109
rect 30098 25100 30104 25152
rect 30156 25140 30162 25152
rect 30668 25140 30696 25171
rect 30156 25112 30696 25140
rect 30156 25100 30162 25112
rect 30834 25100 30840 25152
rect 30892 25140 30898 25152
rect 31021 25143 31079 25149
rect 31021 25140 31033 25143
rect 30892 25112 31033 25140
rect 30892 25100 30898 25112
rect 31021 25109 31033 25112
rect 31067 25109 31079 25143
rect 31021 25103 31079 25109
rect 31294 25100 31300 25152
rect 31352 25100 31358 25152
rect 1104 25050 35328 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35328 25050
rect 1104 24976 35328 24998
rect 4154 24896 4160 24948
rect 4212 24936 4218 24948
rect 4249 24939 4307 24945
rect 4249 24936 4261 24939
rect 4212 24908 4261 24936
rect 4212 24896 4218 24908
rect 4249 24905 4261 24908
rect 4295 24905 4307 24939
rect 4249 24899 4307 24905
rect 4522 24896 4528 24948
rect 4580 24896 4586 24948
rect 4893 24939 4951 24945
rect 4893 24905 4905 24939
rect 4939 24936 4951 24939
rect 5258 24936 5264 24948
rect 4939 24908 5264 24936
rect 4939 24905 4951 24908
rect 4893 24899 4951 24905
rect 5258 24896 5264 24908
rect 5316 24896 5322 24948
rect 6362 24896 6368 24948
rect 6420 24896 6426 24948
rect 6730 24896 6736 24948
rect 6788 24896 6794 24948
rect 9674 24896 9680 24948
rect 9732 24896 9738 24948
rect 10134 24896 10140 24948
rect 10192 24896 10198 24948
rect 10318 24896 10324 24948
rect 10376 24936 10382 24948
rect 10505 24939 10563 24945
rect 10505 24936 10517 24939
rect 10376 24908 10517 24936
rect 10376 24896 10382 24908
rect 10505 24905 10517 24908
rect 10551 24905 10563 24939
rect 10505 24899 10563 24905
rect 11054 24896 11060 24948
rect 11112 24936 11118 24948
rect 14918 24936 14924 24948
rect 11112 24908 14924 24936
rect 11112 24896 11118 24908
rect 14918 24896 14924 24908
rect 14976 24896 14982 24948
rect 15102 24896 15108 24948
rect 15160 24936 15166 24948
rect 15565 24939 15623 24945
rect 15565 24936 15577 24939
rect 15160 24908 15577 24936
rect 15160 24896 15166 24908
rect 15565 24905 15577 24908
rect 15611 24905 15623 24939
rect 15565 24899 15623 24905
rect 16114 24896 16120 24948
rect 16172 24936 16178 24948
rect 19518 24936 19524 24948
rect 16172 24908 19524 24936
rect 16172 24896 16178 24908
rect 19518 24896 19524 24908
rect 19576 24896 19582 24948
rect 19702 24896 19708 24948
rect 19760 24896 19766 24948
rect 19978 24896 19984 24948
rect 20036 24936 20042 24948
rect 20073 24939 20131 24945
rect 20073 24936 20085 24939
rect 20036 24908 20085 24936
rect 20036 24896 20042 24908
rect 20073 24905 20085 24908
rect 20119 24905 20131 24939
rect 20073 24899 20131 24905
rect 21818 24896 21824 24948
rect 21876 24896 21882 24948
rect 22189 24939 22247 24945
rect 22189 24905 22201 24939
rect 22235 24936 22247 24939
rect 22278 24936 22284 24948
rect 22235 24908 22284 24936
rect 22235 24905 22247 24908
rect 22189 24899 22247 24905
rect 22278 24896 22284 24908
rect 22336 24896 22342 24948
rect 23106 24896 23112 24948
rect 23164 24896 23170 24948
rect 23658 24936 23664 24948
rect 23400 24908 23664 24936
rect 3418 24868 3424 24880
rect 2884 24840 3424 24868
rect 2884 24809 2912 24840
rect 3418 24828 3424 24840
rect 3476 24828 3482 24880
rect 8564 24871 8622 24877
rect 8564 24837 8576 24871
rect 8610 24868 8622 24871
rect 8846 24868 8852 24880
rect 8610 24840 8852 24868
rect 8610 24837 8622 24840
rect 8564 24831 8622 24837
rect 8846 24828 8852 24840
rect 8904 24828 8910 24880
rect 10597 24871 10655 24877
rect 10597 24837 10609 24871
rect 10643 24868 10655 24871
rect 10643 24840 10916 24868
rect 10643 24837 10655 24840
rect 10597 24831 10655 24837
rect 2869 24803 2927 24809
rect 2869 24769 2881 24803
rect 2915 24769 2927 24803
rect 2869 24763 2927 24769
rect 3136 24803 3194 24809
rect 3136 24769 3148 24803
rect 3182 24800 3194 24803
rect 3602 24800 3608 24812
rect 3182 24772 3608 24800
rect 3182 24769 3194 24772
rect 3136 24763 3194 24769
rect 3602 24760 3608 24772
rect 3660 24760 3666 24812
rect 4985 24803 5043 24809
rect 4985 24769 4997 24803
rect 5031 24800 5043 24803
rect 5442 24800 5448 24812
rect 5031 24772 5448 24800
rect 5031 24769 5043 24772
rect 4985 24763 5043 24769
rect 5442 24760 5448 24772
rect 5500 24760 5506 24812
rect 6825 24803 6883 24809
rect 6825 24769 6837 24803
rect 6871 24800 6883 24803
rect 6871 24772 9352 24800
rect 6871 24769 6883 24772
rect 6825 24763 6883 24769
rect 5169 24735 5227 24741
rect 5169 24701 5181 24735
rect 5215 24732 5227 24735
rect 5626 24732 5632 24744
rect 5215 24704 5632 24732
rect 5215 24701 5227 24704
rect 5169 24695 5227 24701
rect 5626 24692 5632 24704
rect 5684 24692 5690 24744
rect 3878 24624 3884 24676
rect 3936 24664 3942 24676
rect 6840 24664 6868 24763
rect 7009 24735 7067 24741
rect 7009 24701 7021 24735
rect 7055 24732 7067 24735
rect 7282 24732 7288 24744
rect 7055 24704 7288 24732
rect 7055 24701 7067 24704
rect 7009 24695 7067 24701
rect 7282 24692 7288 24704
rect 7340 24692 7346 24744
rect 8297 24735 8355 24741
rect 8297 24701 8309 24735
rect 8343 24701 8355 24735
rect 9324 24732 9352 24772
rect 10612 24732 10640 24831
rect 10888 24800 10916 24840
rect 10962 24828 10968 24880
rect 11020 24868 11026 24880
rect 13262 24868 13268 24880
rect 11020 24840 13268 24868
rect 11020 24828 11026 24840
rect 13262 24828 13268 24840
rect 13320 24828 13326 24880
rect 15010 24828 15016 24880
rect 15068 24868 15074 24880
rect 15068 24840 15332 24868
rect 15068 24828 15074 24840
rect 12526 24800 12532 24812
rect 10888 24772 12532 24800
rect 12526 24760 12532 24772
rect 12584 24800 12590 24812
rect 12894 24800 12900 24812
rect 12584 24772 12900 24800
rect 12584 24760 12590 24772
rect 12894 24760 12900 24772
rect 12952 24760 12958 24812
rect 13630 24760 13636 24812
rect 13688 24760 13694 24812
rect 13722 24760 13728 24812
rect 13780 24760 13786 24812
rect 13992 24803 14050 24809
rect 13992 24769 14004 24803
rect 14038 24800 14050 24803
rect 15304 24800 15332 24840
rect 16960 24840 17264 24868
rect 15657 24803 15715 24809
rect 15657 24800 15669 24803
rect 14038 24772 15240 24800
rect 15304 24772 15669 24800
rect 14038 24769 14050 24772
rect 13992 24763 14050 24769
rect 9324 24704 10640 24732
rect 10781 24735 10839 24741
rect 8297 24695 8355 24701
rect 10781 24701 10793 24735
rect 10827 24732 10839 24735
rect 11054 24732 11060 24744
rect 10827 24704 11060 24732
rect 10827 24701 10839 24704
rect 10781 24695 10839 24701
rect 3936 24636 6868 24664
rect 3936 24624 3942 24636
rect 8312 24596 8340 24695
rect 11054 24692 11060 24704
rect 11112 24692 11118 24744
rect 10042 24624 10048 24676
rect 10100 24664 10106 24676
rect 15212 24673 15240 24772
rect 15657 24769 15669 24772
rect 15703 24800 15715 24803
rect 16960 24800 16988 24840
rect 15703 24772 16988 24800
rect 17037 24803 17095 24809
rect 15703 24769 15715 24772
rect 15657 24763 15715 24769
rect 17037 24769 17049 24803
rect 17083 24769 17095 24803
rect 17037 24763 17095 24769
rect 15749 24735 15807 24741
rect 15749 24701 15761 24735
rect 15795 24732 15807 24735
rect 16025 24735 16083 24741
rect 16025 24732 16037 24735
rect 15795 24704 16037 24732
rect 15795 24701 15807 24704
rect 15749 24695 15807 24701
rect 16025 24701 16037 24704
rect 16071 24701 16083 24735
rect 16025 24695 16083 24701
rect 15197 24667 15255 24673
rect 10100 24636 12388 24664
rect 10100 24624 10106 24636
rect 9766 24596 9772 24608
rect 8312 24568 9772 24596
rect 9766 24556 9772 24568
rect 9824 24556 9830 24608
rect 10226 24556 10232 24608
rect 10284 24596 10290 24608
rect 11698 24596 11704 24608
rect 10284 24568 11704 24596
rect 10284 24556 10290 24568
rect 11698 24556 11704 24568
rect 11756 24556 11762 24608
rect 12360 24605 12388 24636
rect 15197 24633 15209 24667
rect 15243 24633 15255 24667
rect 15197 24627 15255 24633
rect 12345 24599 12403 24605
rect 12345 24565 12357 24599
rect 12391 24596 12403 24599
rect 14090 24596 14096 24608
rect 12391 24568 14096 24596
rect 12391 24565 12403 24568
rect 12345 24559 12403 24565
rect 14090 24556 14096 24568
rect 14148 24556 14154 24608
rect 14366 24556 14372 24608
rect 14424 24596 14430 24608
rect 15470 24596 15476 24608
rect 14424 24568 15476 24596
rect 14424 24556 14430 24568
rect 15470 24556 15476 24568
rect 15528 24596 15534 24608
rect 15764 24596 15792 24695
rect 15528 24568 15792 24596
rect 15528 24556 15534 24568
rect 16666 24556 16672 24608
rect 16724 24556 16730 24608
rect 17052 24596 17080 24763
rect 17126 24760 17132 24812
rect 17184 24760 17190 24812
rect 17236 24800 17264 24840
rect 19794 24828 19800 24880
rect 19852 24868 19858 24880
rect 23400 24868 23428 24908
rect 23658 24896 23664 24908
rect 23716 24936 23722 24948
rect 25225 24939 25283 24945
rect 25225 24936 25237 24939
rect 23716 24908 25237 24936
rect 23716 24896 23722 24908
rect 24228 24877 24256 24908
rect 25225 24905 25237 24908
rect 25271 24905 25283 24939
rect 25225 24899 25283 24905
rect 25774 24896 25780 24948
rect 25832 24896 25838 24948
rect 26970 24896 26976 24948
rect 27028 24896 27034 24948
rect 27338 24896 27344 24948
rect 27396 24896 27402 24948
rect 27801 24939 27859 24945
rect 27801 24936 27813 24939
rect 27448 24908 27813 24936
rect 19852 24840 23428 24868
rect 23477 24871 23535 24877
rect 19852 24828 19858 24840
rect 23477 24837 23489 24871
rect 23523 24868 23535 24871
rect 24213 24871 24271 24877
rect 23523 24840 24072 24868
rect 23523 24837 23535 24840
rect 23477 24831 23535 24837
rect 24044 24812 24072 24840
rect 24213 24837 24225 24871
rect 24259 24837 24271 24871
rect 25590 24868 25596 24880
rect 24213 24831 24271 24837
rect 24688 24840 25596 24868
rect 17497 24803 17555 24809
rect 17497 24800 17509 24803
rect 17236 24772 17509 24800
rect 17497 24769 17509 24772
rect 17543 24769 17555 24803
rect 17497 24763 17555 24769
rect 20070 24760 20076 24812
rect 20128 24800 20134 24812
rect 20165 24803 20223 24809
rect 20165 24800 20177 24803
rect 20128 24772 20177 24800
rect 20128 24760 20134 24772
rect 20165 24769 20177 24772
rect 20211 24769 20223 24803
rect 20165 24763 20223 24769
rect 21634 24760 21640 24812
rect 21692 24800 21698 24812
rect 22281 24803 22339 24809
rect 22281 24800 22293 24803
rect 21692 24772 22293 24800
rect 21692 24760 21698 24772
rect 22281 24769 22293 24772
rect 22327 24769 22339 24803
rect 22281 24763 22339 24769
rect 22922 24760 22928 24812
rect 22980 24760 22986 24812
rect 23014 24760 23020 24812
rect 23072 24800 23078 24812
rect 23937 24803 23995 24809
rect 23937 24800 23949 24803
rect 23072 24772 23949 24800
rect 23072 24760 23078 24772
rect 23937 24769 23949 24772
rect 23983 24769 23995 24803
rect 23937 24763 23995 24769
rect 24026 24760 24032 24812
rect 24084 24800 24090 24812
rect 24084 24772 24129 24800
rect 24084 24760 24090 24772
rect 24302 24760 24308 24812
rect 24360 24760 24366 24812
rect 24688 24809 24716 24840
rect 25590 24828 25596 24840
rect 25648 24868 25654 24880
rect 25792 24868 25820 24896
rect 25648 24840 25820 24868
rect 25648 24828 25654 24840
rect 26234 24828 26240 24880
rect 26292 24868 26298 24880
rect 27448 24868 27476 24908
rect 27801 24905 27813 24908
rect 27847 24905 27859 24939
rect 27801 24899 27859 24905
rect 28074 24896 28080 24948
rect 28132 24936 28138 24948
rect 28442 24936 28448 24948
rect 28132 24908 28448 24936
rect 28132 24896 28138 24908
rect 28442 24896 28448 24908
rect 28500 24936 28506 24948
rect 29178 24936 29184 24948
rect 28500 24908 29184 24936
rect 28500 24896 28506 24908
rect 29178 24896 29184 24908
rect 29236 24896 29242 24948
rect 30098 24896 30104 24948
rect 30156 24936 30162 24948
rect 30377 24939 30435 24945
rect 30377 24936 30389 24939
rect 30156 24908 30389 24936
rect 30156 24896 30162 24908
rect 30377 24905 30389 24908
rect 30423 24905 30435 24939
rect 30377 24899 30435 24905
rect 27614 24868 27620 24880
rect 26292 24840 27476 24868
rect 27540 24840 27620 24868
rect 26292 24828 26298 24840
rect 24402 24803 24460 24809
rect 24402 24769 24414 24803
rect 24448 24769 24460 24803
rect 24402 24763 24460 24769
rect 24673 24803 24731 24809
rect 24673 24769 24685 24803
rect 24719 24769 24731 24803
rect 24673 24763 24731 24769
rect 17218 24692 17224 24744
rect 17276 24692 17282 24744
rect 17310 24692 17316 24744
rect 17368 24732 17374 24744
rect 17368 24704 20208 24732
rect 17368 24692 17374 24704
rect 17681 24667 17739 24673
rect 17681 24664 17693 24667
rect 17420 24636 17693 24664
rect 17420 24596 17448 24636
rect 17681 24633 17693 24636
rect 17727 24664 17739 24667
rect 18322 24664 18328 24676
rect 17727 24636 18328 24664
rect 17727 24633 17739 24636
rect 17681 24627 17739 24633
rect 18322 24624 18328 24636
rect 18380 24664 18386 24676
rect 20070 24664 20076 24676
rect 18380 24636 20076 24664
rect 18380 24624 18386 24636
rect 20070 24624 20076 24636
rect 20128 24624 20134 24676
rect 20180 24664 20208 24704
rect 20346 24692 20352 24744
rect 20404 24692 20410 24744
rect 22094 24692 22100 24744
rect 22152 24732 22158 24744
rect 22373 24735 22431 24741
rect 22373 24732 22385 24735
rect 22152 24704 22385 24732
rect 22152 24692 22158 24704
rect 22373 24701 22385 24704
rect 22419 24701 22431 24735
rect 22373 24695 22431 24701
rect 22462 24692 22468 24744
rect 22520 24732 22526 24744
rect 22520 24704 23520 24732
rect 22520 24692 22526 24704
rect 20180 24636 22508 24664
rect 17052 24568 17448 24596
rect 17586 24556 17592 24608
rect 17644 24596 17650 24608
rect 17773 24599 17831 24605
rect 17773 24596 17785 24599
rect 17644 24568 17785 24596
rect 17644 24556 17650 24568
rect 17773 24565 17785 24568
rect 17819 24596 17831 24599
rect 19978 24596 19984 24608
rect 17819 24568 19984 24596
rect 17819 24565 17831 24568
rect 17773 24559 17831 24565
rect 19978 24556 19984 24568
rect 20036 24556 20042 24608
rect 20162 24556 20168 24608
rect 20220 24596 20226 24608
rect 22370 24596 22376 24608
rect 20220 24568 22376 24596
rect 20220 24556 20226 24568
rect 22370 24556 22376 24568
rect 22428 24556 22434 24608
rect 22480 24596 22508 24636
rect 22922 24624 22928 24676
rect 22980 24664 22986 24676
rect 23492 24664 23520 24704
rect 23566 24692 23572 24744
rect 23624 24692 23630 24744
rect 23750 24692 23756 24744
rect 23808 24692 23814 24744
rect 24412 24664 24440 24763
rect 24762 24760 24768 24812
rect 24820 24800 24826 24812
rect 25041 24803 25099 24809
rect 25041 24800 25053 24803
rect 24820 24772 25053 24800
rect 24820 24760 24826 24772
rect 25041 24769 25053 24772
rect 25087 24769 25099 24803
rect 25041 24763 25099 24769
rect 25774 24760 25780 24812
rect 25832 24800 25838 24812
rect 26053 24803 26111 24809
rect 26053 24800 26065 24803
rect 25832 24772 26065 24800
rect 25832 24760 25838 24772
rect 26053 24769 26065 24772
rect 26099 24769 26111 24803
rect 26053 24763 26111 24769
rect 26421 24803 26479 24809
rect 26421 24769 26433 24803
rect 26467 24769 26479 24803
rect 26421 24763 26479 24769
rect 26436 24732 26464 24763
rect 27246 24760 27252 24812
rect 27304 24800 27310 24812
rect 27433 24803 27491 24809
rect 27433 24800 27445 24803
rect 27304 24772 27445 24800
rect 27304 24760 27310 24772
rect 27433 24769 27445 24772
rect 27479 24769 27491 24803
rect 27433 24763 27491 24769
rect 24596 24704 26464 24732
rect 26513 24735 26571 24741
rect 24596 24673 24624 24704
rect 26513 24701 26525 24735
rect 26559 24732 26571 24735
rect 26878 24732 26884 24744
rect 26559 24704 26884 24732
rect 26559 24701 26571 24704
rect 26513 24695 26571 24701
rect 26878 24692 26884 24704
rect 26936 24692 26942 24744
rect 26970 24692 26976 24744
rect 27028 24732 27034 24744
rect 27540 24741 27568 24840
rect 27614 24828 27620 24840
rect 27672 24868 27678 24880
rect 28629 24871 28687 24877
rect 28629 24868 28641 24871
rect 27672 24840 28641 24868
rect 27672 24828 27678 24840
rect 28629 24837 28641 24840
rect 28675 24837 28687 24871
rect 28629 24831 28687 24837
rect 28534 24760 28540 24812
rect 28592 24800 28598 24812
rect 28997 24803 29055 24809
rect 28997 24800 29009 24803
rect 28592 24772 29009 24800
rect 28592 24760 28598 24772
rect 28997 24769 29009 24772
rect 29043 24800 29055 24803
rect 29273 24803 29331 24809
rect 29273 24800 29285 24803
rect 29043 24772 29285 24800
rect 29043 24769 29055 24772
rect 28997 24763 29055 24769
rect 29273 24769 29285 24772
rect 29319 24769 29331 24803
rect 29273 24763 29331 24769
rect 29730 24760 29736 24812
rect 29788 24800 29794 24812
rect 29917 24803 29975 24809
rect 29917 24800 29929 24803
rect 29788 24772 29929 24800
rect 29788 24760 29794 24772
rect 29917 24769 29929 24772
rect 29963 24769 29975 24803
rect 29917 24763 29975 24769
rect 30006 24760 30012 24812
rect 30064 24800 30070 24812
rect 30282 24800 30288 24812
rect 30064 24772 30288 24800
rect 30064 24760 30070 24772
rect 30282 24760 30288 24772
rect 30340 24800 30346 24812
rect 30469 24803 30527 24809
rect 30469 24800 30481 24803
rect 30340 24772 30481 24800
rect 30340 24760 30346 24772
rect 30469 24769 30481 24772
rect 30515 24800 30527 24803
rect 30653 24803 30711 24809
rect 30653 24800 30665 24803
rect 30515 24772 30665 24800
rect 30515 24769 30527 24772
rect 30469 24763 30527 24769
rect 30653 24769 30665 24772
rect 30699 24769 30711 24803
rect 30653 24763 30711 24769
rect 30834 24760 30840 24812
rect 30892 24760 30898 24812
rect 31205 24803 31263 24809
rect 31205 24769 31217 24803
rect 31251 24800 31263 24803
rect 31754 24800 31760 24812
rect 31251 24772 31760 24800
rect 31251 24769 31263 24772
rect 31205 24763 31263 24769
rect 31754 24760 31760 24772
rect 31812 24760 31818 24812
rect 27525 24735 27583 24741
rect 27525 24732 27537 24735
rect 27028 24704 27537 24732
rect 27028 24692 27034 24704
rect 27525 24701 27537 24704
rect 27571 24701 27583 24735
rect 27525 24695 27583 24701
rect 27614 24692 27620 24744
rect 27672 24732 27678 24744
rect 28718 24732 28724 24744
rect 27672 24704 28724 24732
rect 27672 24692 27678 24704
rect 28718 24692 28724 24704
rect 28776 24692 28782 24744
rect 28902 24692 28908 24744
rect 28960 24732 28966 24744
rect 29089 24735 29147 24741
rect 29089 24732 29101 24735
rect 28960 24704 29101 24732
rect 28960 24692 28966 24704
rect 29089 24701 29101 24704
rect 29135 24701 29147 24735
rect 29089 24695 29147 24701
rect 30929 24735 30987 24741
rect 30929 24701 30941 24735
rect 30975 24701 30987 24735
rect 30929 24695 30987 24701
rect 31021 24735 31079 24741
rect 31021 24701 31033 24735
rect 31067 24732 31079 24735
rect 31110 24732 31116 24744
rect 31067 24704 31116 24732
rect 31067 24701 31079 24704
rect 31021 24695 31079 24701
rect 22980 24636 23336 24664
rect 23492 24636 24440 24664
rect 22980 24624 22986 24636
rect 22646 24596 22652 24608
rect 22480 24568 22652 24596
rect 22646 24556 22652 24568
rect 22704 24596 22710 24608
rect 22741 24599 22799 24605
rect 22741 24596 22753 24599
rect 22704 24568 22753 24596
rect 22704 24556 22710 24568
rect 22741 24565 22753 24568
rect 22787 24596 22799 24599
rect 23198 24596 23204 24608
rect 22787 24568 23204 24596
rect 22787 24565 22799 24568
rect 22741 24559 22799 24565
rect 23198 24556 23204 24568
rect 23256 24556 23262 24608
rect 23308 24596 23336 24636
rect 24026 24596 24032 24608
rect 23308 24568 24032 24596
rect 24026 24556 24032 24568
rect 24084 24556 24090 24608
rect 24412 24596 24440 24636
rect 24581 24667 24639 24673
rect 24581 24633 24593 24667
rect 24627 24633 24639 24667
rect 24581 24627 24639 24633
rect 26050 24624 26056 24676
rect 26108 24664 26114 24676
rect 26789 24667 26847 24673
rect 26108 24636 26464 24664
rect 26108 24624 26114 24636
rect 24857 24599 24915 24605
rect 24857 24596 24869 24599
rect 24412 24568 24869 24596
rect 24857 24565 24869 24568
rect 24903 24596 24915 24599
rect 25409 24599 25467 24605
rect 25409 24596 25421 24599
rect 24903 24568 25421 24596
rect 24903 24565 24915 24568
rect 24857 24559 24915 24565
rect 25409 24565 25421 24568
rect 25455 24596 25467 24599
rect 25593 24599 25651 24605
rect 25593 24596 25605 24599
rect 25455 24568 25605 24596
rect 25455 24565 25467 24568
rect 25409 24559 25467 24565
rect 25593 24565 25605 24568
rect 25639 24565 25651 24599
rect 25593 24559 25651 24565
rect 25869 24599 25927 24605
rect 25869 24565 25881 24599
rect 25915 24596 25927 24599
rect 26142 24596 26148 24608
rect 25915 24568 26148 24596
rect 25915 24565 25927 24568
rect 25869 24559 25927 24565
rect 26142 24556 26148 24568
rect 26200 24556 26206 24608
rect 26234 24556 26240 24608
rect 26292 24556 26298 24608
rect 26436 24605 26464 24636
rect 26789 24633 26801 24667
rect 26835 24664 26847 24667
rect 30944 24664 30972 24695
rect 31110 24692 31116 24704
rect 31168 24732 31174 24744
rect 31168 24704 31524 24732
rect 31168 24692 31174 24704
rect 26835 24636 30972 24664
rect 26835 24633 26847 24636
rect 26789 24627 26847 24633
rect 31496 24608 31524 24704
rect 26421 24599 26479 24605
rect 26421 24565 26433 24599
rect 26467 24565 26479 24599
rect 26421 24559 26479 24565
rect 27062 24556 27068 24608
rect 27120 24596 27126 24608
rect 27985 24599 28043 24605
rect 27985 24596 27997 24599
rect 27120 24568 27997 24596
rect 27120 24556 27126 24568
rect 27985 24565 27997 24568
rect 28031 24596 28043 24599
rect 28074 24596 28080 24608
rect 28031 24568 28080 24596
rect 28031 24565 28043 24568
rect 27985 24559 28043 24565
rect 28074 24556 28080 24568
rect 28132 24556 28138 24608
rect 28166 24556 28172 24608
rect 28224 24556 28230 24608
rect 28350 24556 28356 24608
rect 28408 24556 28414 24608
rect 28810 24556 28816 24608
rect 28868 24556 28874 24608
rect 29730 24556 29736 24608
rect 29788 24556 29794 24608
rect 31386 24556 31392 24608
rect 31444 24556 31450 24608
rect 31478 24556 31484 24608
rect 31536 24556 31542 24608
rect 1104 24506 35328 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 35328 24506
rect 1104 24432 35328 24454
rect 10042 24352 10048 24404
rect 10100 24352 10106 24404
rect 12158 24352 12164 24404
rect 12216 24352 12222 24404
rect 14182 24352 14188 24404
rect 14240 24352 14246 24404
rect 16574 24392 16580 24404
rect 14660 24364 16580 24392
rect 3973 24327 4031 24333
rect 3973 24293 3985 24327
rect 4019 24324 4031 24327
rect 5442 24324 5448 24336
rect 4019 24296 5448 24324
rect 4019 24293 4031 24296
rect 3973 24287 4031 24293
rect 5442 24284 5448 24296
rect 5500 24284 5506 24336
rect 7009 24327 7067 24333
rect 7009 24324 7021 24327
rect 6748 24296 7021 24324
rect 6748 24265 6776 24296
rect 7009 24293 7021 24296
rect 7055 24324 7067 24327
rect 11146 24324 11152 24336
rect 7055 24296 11152 24324
rect 7055 24293 7067 24296
rect 7009 24287 7067 24293
rect 11146 24284 11152 24296
rect 11204 24324 11210 24336
rect 12250 24324 12256 24336
rect 11204 24296 12256 24324
rect 11204 24284 11210 24296
rect 12250 24284 12256 24296
rect 12308 24284 12314 24336
rect 13081 24327 13139 24333
rect 13081 24324 13093 24327
rect 12820 24296 13093 24324
rect 6733 24259 6791 24265
rect 2746 24228 4752 24256
rect 1210 24148 1216 24200
rect 1268 24188 1274 24200
rect 1397 24191 1455 24197
rect 1397 24188 1409 24191
rect 1268 24160 1409 24188
rect 1268 24148 1274 24160
rect 1397 24157 1409 24160
rect 1443 24188 1455 24191
rect 1673 24191 1731 24197
rect 1673 24188 1685 24191
rect 1443 24160 1685 24188
rect 1443 24157 1455 24160
rect 1397 24151 1455 24157
rect 1673 24157 1685 24160
rect 1719 24157 1731 24191
rect 1673 24151 1731 24157
rect 2746 24120 2774 24228
rect 4724 24197 4752 24228
rect 6733 24225 6745 24259
rect 6779 24225 6791 24259
rect 6733 24219 6791 24225
rect 9674 24216 9680 24268
rect 9732 24256 9738 24268
rect 11054 24256 11060 24268
rect 9732 24228 11060 24256
rect 9732 24216 9738 24228
rect 11054 24216 11060 24228
rect 11112 24216 11118 24268
rect 12710 24216 12716 24268
rect 12768 24256 12774 24268
rect 12820 24265 12848 24296
rect 13081 24293 13093 24296
rect 13127 24324 13139 24327
rect 13170 24324 13176 24336
rect 13127 24296 13176 24324
rect 13127 24293 13139 24296
rect 13081 24287 13139 24293
rect 13170 24284 13176 24296
rect 13228 24324 13234 24336
rect 14660 24324 14688 24364
rect 16574 24352 16580 24364
rect 16632 24352 16638 24404
rect 17126 24352 17132 24404
rect 17184 24392 17190 24404
rect 17313 24395 17371 24401
rect 17313 24392 17325 24395
rect 17184 24364 17325 24392
rect 17184 24352 17190 24364
rect 17313 24361 17325 24364
rect 17359 24361 17371 24395
rect 17313 24355 17371 24361
rect 19610 24352 19616 24404
rect 19668 24392 19674 24404
rect 19797 24395 19855 24401
rect 19797 24392 19809 24395
rect 19668 24364 19809 24392
rect 19668 24352 19674 24364
rect 19797 24361 19809 24364
rect 19843 24361 19855 24395
rect 19797 24355 19855 24361
rect 19886 24352 19892 24404
rect 19944 24352 19950 24404
rect 19978 24352 19984 24404
rect 20036 24392 20042 24404
rect 20036 24364 22416 24392
rect 20036 24352 20042 24364
rect 13228 24296 14688 24324
rect 13228 24284 13234 24296
rect 19518 24284 19524 24336
rect 19576 24324 19582 24336
rect 21726 24324 21732 24336
rect 19576 24296 21732 24324
rect 19576 24284 19582 24296
rect 21726 24284 21732 24296
rect 21784 24284 21790 24336
rect 12805 24259 12863 24265
rect 12805 24256 12817 24259
rect 12768 24228 12817 24256
rect 12768 24216 12774 24228
rect 12805 24225 12817 24228
rect 12851 24225 12863 24259
rect 12805 24219 12863 24225
rect 12894 24216 12900 24268
rect 12952 24256 12958 24268
rect 13538 24256 13544 24268
rect 12952 24228 13544 24256
rect 12952 24216 12958 24228
rect 13538 24216 13544 24228
rect 13596 24256 13602 24268
rect 13596 24228 16059 24256
rect 13596 24216 13602 24228
rect 3789 24191 3847 24197
rect 3789 24157 3801 24191
rect 3835 24188 3847 24191
rect 4709 24191 4767 24197
rect 3835 24160 4660 24188
rect 3835 24157 3847 24160
rect 3789 24151 3847 24157
rect 1596 24092 2774 24120
rect 1596 24061 1624 24092
rect 3418 24080 3424 24132
rect 3476 24120 3482 24132
rect 3878 24120 3884 24132
rect 3476 24092 3884 24120
rect 3476 24080 3482 24092
rect 3878 24080 3884 24092
rect 3936 24120 3942 24132
rect 4249 24123 4307 24129
rect 4249 24120 4261 24123
rect 3936 24092 4261 24120
rect 3936 24080 3942 24092
rect 4249 24089 4261 24092
rect 4295 24089 4307 24123
rect 4249 24083 4307 24089
rect 1581 24055 1639 24061
rect 1581 24021 1593 24055
rect 1627 24021 1639 24055
rect 4632 24052 4660 24160
rect 4709 24157 4721 24191
rect 4755 24157 4767 24191
rect 4709 24151 4767 24157
rect 9125 24191 9183 24197
rect 9125 24157 9137 24191
rect 9171 24188 9183 24191
rect 9766 24188 9772 24200
rect 9171 24160 9772 24188
rect 9171 24157 9183 24160
rect 9125 24151 9183 24157
rect 9766 24148 9772 24160
rect 9824 24148 9830 24200
rect 11609 24191 11667 24197
rect 11609 24188 11621 24191
rect 9876 24160 11621 24188
rect 8294 24120 8300 24132
rect 4908 24092 8300 24120
rect 4908 24061 4936 24092
rect 8294 24080 8300 24092
rect 8352 24120 8358 24132
rect 9876 24120 9904 24160
rect 11609 24157 11621 24160
rect 11655 24188 11667 24191
rect 11655 24160 12434 24188
rect 11655 24157 11667 24160
rect 11609 24151 11667 24157
rect 12406 24120 12434 24160
rect 12526 24148 12532 24200
rect 12584 24148 12590 24200
rect 12621 24191 12679 24197
rect 12621 24157 12633 24191
rect 12667 24188 12679 24191
rect 12986 24188 12992 24200
rect 12667 24160 12992 24188
rect 12667 24157 12679 24160
rect 12621 24151 12679 24157
rect 12986 24148 12992 24160
rect 13044 24148 13050 24200
rect 15930 24148 15936 24200
rect 15988 24148 15994 24200
rect 16031 24188 16059 24228
rect 17494 24216 17500 24268
rect 17552 24256 17558 24268
rect 22002 24256 22008 24268
rect 17552 24228 22008 24256
rect 17552 24216 17558 24228
rect 22002 24216 22008 24228
rect 22060 24216 22066 24268
rect 22278 24216 22284 24268
rect 22336 24216 22342 24268
rect 22388 24256 22416 24364
rect 22462 24352 22468 24404
rect 22520 24392 22526 24404
rect 22741 24395 22799 24401
rect 22741 24392 22753 24395
rect 22520 24364 22753 24392
rect 22520 24352 22526 24364
rect 22741 24361 22753 24364
rect 22787 24361 22799 24395
rect 22741 24355 22799 24361
rect 23750 24352 23756 24404
rect 23808 24392 23814 24404
rect 24486 24392 24492 24404
rect 23808 24364 24492 24392
rect 23808 24352 23814 24364
rect 24486 24352 24492 24364
rect 24544 24352 24550 24404
rect 25682 24352 25688 24404
rect 25740 24392 25746 24404
rect 26697 24395 26755 24401
rect 26697 24392 26709 24395
rect 25740 24364 26709 24392
rect 25740 24352 25746 24364
rect 26697 24361 26709 24364
rect 26743 24361 26755 24395
rect 26697 24355 26755 24361
rect 22649 24327 22707 24333
rect 22649 24293 22661 24327
rect 22695 24324 22707 24327
rect 23014 24324 23020 24336
rect 22695 24296 23020 24324
rect 22695 24293 22707 24296
rect 22649 24287 22707 24293
rect 23014 24284 23020 24296
rect 23072 24284 23078 24336
rect 23198 24284 23204 24336
rect 23256 24324 23262 24336
rect 23845 24327 23903 24333
rect 23845 24324 23857 24327
rect 23256 24296 23857 24324
rect 23256 24284 23262 24296
rect 23845 24293 23857 24296
rect 23891 24293 23903 24327
rect 26234 24324 26240 24336
rect 23845 24287 23903 24293
rect 25792 24296 26240 24324
rect 25409 24259 25467 24265
rect 25409 24256 25421 24259
rect 22388 24228 25421 24256
rect 25409 24225 25421 24228
rect 25455 24256 25467 24259
rect 25682 24256 25688 24268
rect 25455 24228 25688 24256
rect 25455 24225 25467 24228
rect 25409 24219 25467 24225
rect 25682 24216 25688 24228
rect 25740 24216 25746 24268
rect 16031 24160 16804 24188
rect 13446 24120 13452 24132
rect 8352 24092 9904 24120
rect 11440 24092 12296 24120
rect 12406 24092 13452 24120
rect 8352 24080 8358 24092
rect 4893 24055 4951 24061
rect 4893 24052 4905 24055
rect 4632 24024 4905 24052
rect 1581 24015 1639 24021
rect 4893 24021 4905 24024
rect 4939 24021 4951 24055
rect 4893 24015 4951 24021
rect 6086 24012 6092 24064
rect 6144 24012 6150 24064
rect 6454 24012 6460 24064
rect 6512 24012 6518 24064
rect 6549 24055 6607 24061
rect 6549 24021 6561 24055
rect 6595 24052 6607 24055
rect 6638 24052 6644 24064
rect 6595 24024 6644 24052
rect 6595 24021 6607 24024
rect 6549 24015 6607 24021
rect 6638 24012 6644 24024
rect 6696 24012 6702 24064
rect 11440 24061 11468 24092
rect 11425 24055 11483 24061
rect 11425 24021 11437 24055
rect 11471 24021 11483 24055
rect 12268 24052 12296 24092
rect 13446 24080 13452 24092
rect 13504 24080 13510 24132
rect 16200 24123 16258 24129
rect 16200 24089 16212 24123
rect 16246 24120 16258 24123
rect 16666 24120 16672 24132
rect 16246 24092 16672 24120
rect 16246 24089 16258 24092
rect 16200 24083 16258 24089
rect 16666 24080 16672 24092
rect 16724 24080 16730 24132
rect 16776 24120 16804 24160
rect 19242 24148 19248 24200
rect 19300 24148 19306 24200
rect 19613 24191 19671 24197
rect 19613 24188 19625 24191
rect 19352 24160 19625 24188
rect 19352 24120 19380 24160
rect 19613 24157 19625 24160
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 16776 24092 19380 24120
rect 19429 24123 19487 24129
rect 19429 24089 19441 24123
rect 19475 24089 19487 24123
rect 19429 24083 19487 24089
rect 12434 24052 12440 24064
rect 12268 24024 12440 24052
rect 11425 24015 11483 24021
rect 12434 24012 12440 24024
rect 12492 24012 12498 24064
rect 13630 24012 13636 24064
rect 13688 24052 13694 24064
rect 13725 24055 13783 24061
rect 13725 24052 13737 24055
rect 13688 24024 13737 24052
rect 13688 24012 13694 24024
rect 13725 24021 13737 24024
rect 13771 24021 13783 24055
rect 19444 24052 19472 24083
rect 19518 24080 19524 24132
rect 19576 24080 19582 24132
rect 19628 24120 19656 24151
rect 20070 24148 20076 24200
rect 20128 24148 20134 24200
rect 21913 24191 21971 24197
rect 21913 24157 21925 24191
rect 21959 24157 21971 24191
rect 21913 24151 21971 24157
rect 20162 24120 20168 24132
rect 19628 24092 20168 24120
rect 20162 24080 20168 24092
rect 20220 24080 20226 24132
rect 19886 24052 19892 24064
rect 19444 24024 19892 24052
rect 13725 24015 13783 24021
rect 19886 24012 19892 24024
rect 19944 24012 19950 24064
rect 21928 24052 21956 24151
rect 22094 24148 22100 24200
rect 22152 24148 22158 24200
rect 22296 24188 22324 24216
rect 22373 24191 22431 24197
rect 22373 24188 22385 24191
rect 22296 24160 22385 24188
rect 22373 24157 22385 24160
rect 22419 24157 22431 24191
rect 22373 24151 22431 24157
rect 22465 24191 22523 24197
rect 22465 24157 22477 24191
rect 22511 24188 22523 24191
rect 22922 24188 22928 24200
rect 22511 24160 22928 24188
rect 22511 24157 22523 24160
rect 22465 24151 22523 24157
rect 22922 24148 22928 24160
rect 22980 24188 22986 24200
rect 23106 24188 23112 24200
rect 22980 24160 23112 24188
rect 22980 24148 22986 24160
rect 23106 24148 23112 24160
rect 23164 24148 23170 24200
rect 23290 24148 23296 24200
rect 23348 24148 23354 24200
rect 23474 24148 23480 24200
rect 23532 24188 23538 24200
rect 23750 24188 23756 24200
rect 23532 24160 23756 24188
rect 23532 24148 23538 24160
rect 23750 24148 23756 24160
rect 23808 24148 23814 24200
rect 23842 24148 23848 24200
rect 23900 24188 23906 24200
rect 25225 24191 25283 24197
rect 23900 24160 25176 24188
rect 23900 24148 23906 24160
rect 22281 24123 22339 24129
rect 22281 24089 22293 24123
rect 22327 24120 22339 24123
rect 22646 24120 22652 24132
rect 22327 24092 22652 24120
rect 22327 24089 22339 24092
rect 22281 24083 22339 24089
rect 22646 24080 22652 24092
rect 22704 24080 22710 24132
rect 24397 24123 24455 24129
rect 24397 24120 24409 24123
rect 23676 24092 24409 24120
rect 22925 24055 22983 24061
rect 22925 24052 22937 24055
rect 21928 24024 22937 24052
rect 22925 24021 22937 24024
rect 22971 24052 22983 24055
rect 23198 24052 23204 24064
rect 22971 24024 23204 24052
rect 22971 24021 22983 24024
rect 22925 24015 22983 24021
rect 23198 24012 23204 24024
rect 23256 24012 23262 24064
rect 23566 24012 23572 24064
rect 23624 24052 23630 24064
rect 23676 24061 23704 24092
rect 24397 24089 24409 24092
rect 24443 24089 24455 24123
rect 25148 24120 25176 24160
rect 25225 24157 25237 24191
rect 25271 24188 25283 24191
rect 25314 24188 25320 24200
rect 25271 24160 25320 24188
rect 25271 24157 25283 24160
rect 25225 24151 25283 24157
rect 25314 24148 25320 24160
rect 25372 24148 25378 24200
rect 25792 24197 25820 24296
rect 26234 24284 26240 24296
rect 26292 24284 26298 24336
rect 26421 24327 26479 24333
rect 26421 24293 26433 24327
rect 26467 24293 26479 24327
rect 26712 24324 26740 24355
rect 26878 24352 26884 24404
rect 26936 24352 26942 24404
rect 27246 24352 27252 24404
rect 27304 24392 27310 24404
rect 27304 24364 27844 24392
rect 27304 24352 27310 24364
rect 27816 24324 27844 24364
rect 28074 24352 28080 24404
rect 28132 24392 28138 24404
rect 28442 24392 28448 24404
rect 28132 24364 28448 24392
rect 28132 24352 28138 24364
rect 28442 24352 28448 24364
rect 28500 24352 28506 24404
rect 28534 24352 28540 24404
rect 28592 24352 28598 24404
rect 28718 24352 28724 24404
rect 28776 24352 28782 24404
rect 29270 24392 29276 24404
rect 29012 24364 29276 24392
rect 29012 24336 29040 24364
rect 29270 24352 29276 24364
rect 29328 24352 29334 24404
rect 29917 24395 29975 24401
rect 29917 24361 29929 24395
rect 29963 24392 29975 24395
rect 30558 24392 30564 24404
rect 29963 24364 30564 24392
rect 29963 24361 29975 24364
rect 29917 24355 29975 24361
rect 30558 24352 30564 24364
rect 30616 24352 30622 24404
rect 31754 24352 31760 24404
rect 31812 24352 31818 24404
rect 28994 24324 29000 24336
rect 26712 24296 27752 24324
rect 27816 24296 29000 24324
rect 26421 24287 26479 24293
rect 26142 24256 26148 24268
rect 26068 24228 26148 24256
rect 25958 24197 25964 24200
rect 25777 24191 25835 24197
rect 25777 24157 25789 24191
rect 25823 24157 25835 24191
rect 25777 24151 25835 24157
rect 25925 24191 25964 24197
rect 25925 24157 25937 24191
rect 25925 24151 25964 24157
rect 25792 24120 25820 24151
rect 25958 24148 25964 24151
rect 26016 24148 26022 24200
rect 26068 24197 26096 24228
rect 26142 24216 26148 24228
rect 26200 24216 26206 24268
rect 26436 24256 26464 24287
rect 27724 24256 27752 24296
rect 28994 24284 29000 24296
rect 29052 24284 29058 24336
rect 28166 24256 28172 24268
rect 26436 24228 27568 24256
rect 27724 24228 28172 24256
rect 26053 24191 26111 24197
rect 26053 24157 26065 24191
rect 26099 24157 26111 24191
rect 26053 24151 26111 24157
rect 26234 24148 26240 24200
rect 26292 24197 26298 24200
rect 26292 24188 26300 24197
rect 26292 24160 26337 24188
rect 26292 24151 26300 24160
rect 26292 24148 26298 24151
rect 26510 24148 26516 24200
rect 26568 24148 26574 24200
rect 27062 24197 27068 24200
rect 27060 24188 27068 24197
rect 27023 24160 27068 24188
rect 27060 24151 27068 24160
rect 27062 24148 27068 24151
rect 27120 24148 27126 24200
rect 27246 24148 27252 24200
rect 27304 24148 27310 24200
rect 27338 24148 27344 24200
rect 27396 24197 27402 24200
rect 27540 24197 27568 24228
rect 28166 24216 28172 24228
rect 28224 24216 28230 24268
rect 27396 24191 27435 24197
rect 27423 24157 27435 24191
rect 27396 24151 27435 24157
rect 27525 24191 27583 24197
rect 27525 24157 27537 24191
rect 27571 24157 27583 24191
rect 27525 24151 27583 24157
rect 27396 24148 27402 24151
rect 27614 24148 27620 24200
rect 27672 24148 27678 24200
rect 27798 24148 27804 24200
rect 27856 24188 27862 24200
rect 27985 24191 28043 24197
rect 27985 24188 27997 24191
rect 27856 24160 27997 24188
rect 27856 24148 27862 24160
rect 27985 24157 27997 24160
rect 28031 24157 28043 24191
rect 27985 24151 28043 24157
rect 28074 24148 28080 24200
rect 28132 24188 28138 24200
rect 28353 24191 28411 24197
rect 28353 24188 28365 24191
rect 28132 24160 28365 24188
rect 28132 24148 28138 24160
rect 28353 24157 28365 24160
rect 28399 24157 28411 24191
rect 28353 24151 28411 24157
rect 28718 24148 28724 24200
rect 28776 24188 28782 24200
rect 28902 24188 28908 24200
rect 28776 24160 28908 24188
rect 28776 24148 28782 24160
rect 28902 24148 28908 24160
rect 28960 24148 28966 24200
rect 29638 24148 29644 24200
rect 29696 24148 29702 24200
rect 29733 24191 29791 24197
rect 29733 24157 29745 24191
rect 29779 24157 29791 24191
rect 29733 24151 29791 24157
rect 30377 24191 30435 24197
rect 30377 24157 30389 24191
rect 30423 24188 30435 24191
rect 32766 24188 32772 24200
rect 30423 24160 32772 24188
rect 30423 24157 30435 24160
rect 30377 24151 30435 24157
rect 25148 24092 25820 24120
rect 26145 24123 26203 24129
rect 24397 24083 24455 24089
rect 26145 24089 26157 24123
rect 26191 24089 26203 24123
rect 26145 24083 26203 24089
rect 23661 24055 23719 24061
rect 23661 24052 23673 24055
rect 23624 24024 23673 24052
rect 23624 24012 23630 24024
rect 23661 24021 23673 24024
rect 23707 24021 23719 24055
rect 23661 24015 23719 24021
rect 24026 24012 24032 24064
rect 24084 24012 24090 24064
rect 24673 24055 24731 24061
rect 24673 24021 24685 24055
rect 24719 24052 24731 24055
rect 24762 24052 24768 24064
rect 24719 24024 24768 24052
rect 24719 24021 24731 24024
rect 24673 24015 24731 24021
rect 24762 24012 24768 24024
rect 24820 24012 24826 24064
rect 24854 24012 24860 24064
rect 24912 24012 24918 24064
rect 25317 24055 25375 24061
rect 25317 24021 25329 24055
rect 25363 24052 25375 24055
rect 25774 24052 25780 24064
rect 25363 24024 25780 24052
rect 25363 24021 25375 24024
rect 25317 24015 25375 24021
rect 25774 24012 25780 24024
rect 25832 24052 25838 24064
rect 26160 24052 26188 24083
rect 27154 24080 27160 24132
rect 27212 24080 27218 24132
rect 28810 24120 28816 24132
rect 27347 24092 28816 24120
rect 25832 24024 26188 24052
rect 25832 24012 25838 24024
rect 26234 24012 26240 24064
rect 26292 24052 26298 24064
rect 27347 24052 27375 24092
rect 26292 24024 27375 24052
rect 26292 24012 26298 24024
rect 27798 24012 27804 24064
rect 27856 24012 27862 24064
rect 28184 24061 28212 24092
rect 28810 24080 28816 24092
rect 28868 24080 28874 24132
rect 28994 24080 29000 24132
rect 29052 24080 29058 24132
rect 29270 24080 29276 24132
rect 29328 24120 29334 24132
rect 29748 24120 29776 24151
rect 32766 24148 32772 24160
rect 32824 24148 32830 24200
rect 30650 24129 30656 24132
rect 30009 24123 30067 24129
rect 30009 24120 30021 24123
rect 29328 24092 30021 24120
rect 29328 24080 29334 24092
rect 30009 24089 30021 24092
rect 30055 24089 30067 24123
rect 30009 24083 30067 24089
rect 30644 24083 30656 24129
rect 30650 24080 30656 24083
rect 30708 24080 30714 24132
rect 33042 24080 33048 24132
rect 33100 24080 33106 24132
rect 33502 24080 33508 24132
rect 33560 24080 33566 24132
rect 28169 24055 28227 24061
rect 28169 24021 28181 24055
rect 28215 24021 28227 24055
rect 28169 24015 28227 24021
rect 28350 24012 28356 24064
rect 28408 24052 28414 24064
rect 29181 24055 29239 24061
rect 29181 24052 29193 24055
rect 28408 24024 29193 24052
rect 28408 24012 28414 24024
rect 29181 24021 29193 24024
rect 29227 24021 29239 24055
rect 29181 24015 29239 24021
rect 34514 24012 34520 24064
rect 34572 24012 34578 24064
rect 1104 23962 35328 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35328 23962
rect 1104 23888 35328 23910
rect 5353 23851 5411 23857
rect 5353 23817 5365 23851
rect 5399 23817 5411 23851
rect 5353 23811 5411 23817
rect 4148 23783 4206 23789
rect 2424 23752 3924 23780
rect 2424 23721 2452 23752
rect 3896 23724 3924 23752
rect 4148 23749 4160 23783
rect 4194 23780 4206 23783
rect 5368 23780 5396 23811
rect 5442 23808 5448 23860
rect 5500 23848 5506 23860
rect 5813 23851 5871 23857
rect 5813 23848 5825 23851
rect 5500 23820 5825 23848
rect 5500 23808 5506 23820
rect 5813 23817 5825 23820
rect 5859 23848 5871 23851
rect 6638 23848 6644 23860
rect 5859 23820 6644 23848
rect 5859 23817 5871 23820
rect 5813 23811 5871 23817
rect 6638 23808 6644 23820
rect 6696 23808 6702 23860
rect 10134 23848 10140 23860
rect 6748 23820 10140 23848
rect 4194 23752 5396 23780
rect 6457 23783 6515 23789
rect 4194 23749 4206 23752
rect 4148 23743 4206 23749
rect 6457 23749 6469 23783
rect 6503 23780 6515 23783
rect 6748 23780 6776 23820
rect 10134 23808 10140 23820
rect 10192 23808 10198 23860
rect 11517 23851 11575 23857
rect 11517 23817 11529 23851
rect 11563 23817 11575 23851
rect 11517 23811 11575 23817
rect 12437 23851 12495 23857
rect 12437 23817 12449 23851
rect 12483 23848 12495 23851
rect 12710 23848 12716 23860
rect 12483 23820 12716 23848
rect 12483 23817 12495 23820
rect 12437 23811 12495 23817
rect 10220 23783 10278 23789
rect 6503 23752 6776 23780
rect 6840 23752 9812 23780
rect 6503 23749 6515 23752
rect 6457 23743 6515 23749
rect 2409 23715 2467 23721
rect 2409 23681 2421 23715
rect 2455 23681 2467 23715
rect 2409 23675 2467 23681
rect 2676 23715 2734 23721
rect 2676 23681 2688 23715
rect 2722 23712 2734 23715
rect 3786 23712 3792 23724
rect 2722 23684 3792 23712
rect 2722 23681 2734 23684
rect 2676 23675 2734 23681
rect 3786 23672 3792 23684
rect 3844 23672 3850 23724
rect 3878 23672 3884 23724
rect 3936 23672 3942 23724
rect 5258 23672 5264 23724
rect 5316 23712 5322 23724
rect 5721 23715 5779 23721
rect 5721 23712 5733 23715
rect 5316 23684 5733 23712
rect 5316 23672 5322 23684
rect 5721 23681 5733 23684
rect 5767 23681 5779 23715
rect 5721 23675 5779 23681
rect 5997 23647 6055 23653
rect 5997 23613 6009 23647
rect 6043 23644 6055 23647
rect 6472 23644 6500 23743
rect 6641 23715 6699 23721
rect 6641 23681 6653 23715
rect 6687 23712 6699 23715
rect 6840 23712 6868 23752
rect 6687 23684 6868 23712
rect 6908 23715 6966 23721
rect 6687 23681 6699 23684
rect 6641 23675 6699 23681
rect 6908 23681 6920 23715
rect 6954 23712 6966 23715
rect 7190 23712 7196 23724
rect 6954 23684 7196 23712
rect 6954 23681 6966 23684
rect 6908 23675 6966 23681
rect 7190 23672 7196 23684
rect 7248 23672 7254 23724
rect 8294 23672 8300 23724
rect 8352 23672 8358 23724
rect 8496 23721 8524 23752
rect 9784 23724 9812 23752
rect 10220 23749 10232 23783
rect 10266 23780 10278 23783
rect 11532 23780 11560 23811
rect 12710 23808 12716 23820
rect 12768 23808 12774 23860
rect 13262 23808 13268 23860
rect 13320 23848 13326 23860
rect 13541 23851 13599 23857
rect 13541 23848 13553 23851
rect 13320 23820 13553 23848
rect 13320 23808 13326 23820
rect 13541 23817 13553 23820
rect 13587 23817 13599 23851
rect 13541 23811 13599 23817
rect 13817 23851 13875 23857
rect 13817 23817 13829 23851
rect 13863 23848 13875 23851
rect 19150 23848 19156 23860
rect 13863 23820 19156 23848
rect 13863 23817 13875 23820
rect 13817 23811 13875 23817
rect 10266 23752 11560 23780
rect 10266 23749 10278 23752
rect 10220 23743 10278 23749
rect 8481 23715 8539 23721
rect 8481 23681 8493 23715
rect 8527 23681 8539 23715
rect 8481 23675 8539 23681
rect 8748 23715 8806 23721
rect 8748 23681 8760 23715
rect 8794 23712 8806 23715
rect 9030 23712 9036 23724
rect 8794 23684 9036 23712
rect 8794 23681 8806 23684
rect 8748 23675 8806 23681
rect 9030 23672 9036 23684
rect 9088 23672 9094 23724
rect 9766 23672 9772 23724
rect 9824 23712 9830 23724
rect 9953 23715 10011 23721
rect 9953 23712 9965 23715
rect 9824 23684 9965 23712
rect 9824 23672 9830 23684
rect 9953 23681 9965 23684
rect 9999 23681 10011 23715
rect 9953 23675 10011 23681
rect 11885 23715 11943 23721
rect 11885 23681 11897 23715
rect 11931 23712 11943 23715
rect 12434 23712 12440 23724
rect 11931 23684 12440 23712
rect 11931 23681 11943 23684
rect 11885 23675 11943 23681
rect 12434 23672 12440 23684
rect 12492 23712 12498 23724
rect 13170 23712 13176 23724
rect 12492 23684 13176 23712
rect 12492 23672 12498 23684
rect 13170 23672 13176 23684
rect 13228 23672 13234 23724
rect 13449 23715 13507 23721
rect 13449 23681 13461 23715
rect 13495 23712 13507 23715
rect 13832 23712 13860 23811
rect 19150 23808 19156 23820
rect 19208 23808 19214 23860
rect 19518 23808 19524 23860
rect 19576 23848 19582 23860
rect 20349 23851 20407 23857
rect 20349 23848 20361 23851
rect 19576 23820 20361 23848
rect 19576 23808 19582 23820
rect 20349 23817 20361 23820
rect 20395 23817 20407 23851
rect 20349 23811 20407 23817
rect 20456 23820 21956 23848
rect 15657 23783 15715 23789
rect 15657 23749 15669 23783
rect 15703 23780 15715 23783
rect 15746 23780 15752 23792
rect 15703 23752 15752 23780
rect 15703 23749 15715 23752
rect 15657 23743 15715 23749
rect 15746 23740 15752 23752
rect 15804 23740 15810 23792
rect 19236 23783 19294 23789
rect 17420 23752 19012 23780
rect 13495 23684 13860 23712
rect 15473 23715 15531 23721
rect 13495 23681 13507 23684
rect 13449 23675 13507 23681
rect 15473 23681 15485 23715
rect 15519 23681 15531 23715
rect 15473 23675 15531 23681
rect 11977 23647 12035 23653
rect 11977 23644 11989 23647
rect 6043 23616 6500 23644
rect 11348 23616 11989 23644
rect 6043 23613 6055 23616
rect 5997 23607 6055 23613
rect 11348 23588 11376 23616
rect 11977 23613 11989 23616
rect 12023 23613 12035 23647
rect 11977 23607 12035 23613
rect 12161 23647 12219 23653
rect 12161 23613 12173 23647
rect 12207 23644 12219 23647
rect 12710 23644 12716 23656
rect 12207 23616 12716 23644
rect 12207 23613 12219 23616
rect 12161 23607 12219 23613
rect 12710 23604 12716 23616
rect 12768 23604 12774 23656
rect 15488 23644 15516 23675
rect 15930 23672 15936 23724
rect 15988 23712 15994 23724
rect 17420 23721 17448 23752
rect 18984 23724 19012 23752
rect 19236 23749 19248 23783
rect 19282 23780 19294 23783
rect 19334 23780 19340 23792
rect 19282 23752 19340 23780
rect 19282 23749 19294 23752
rect 19236 23743 19294 23749
rect 19334 23740 19340 23752
rect 19392 23740 19398 23792
rect 17405 23715 17463 23721
rect 17405 23712 17417 23715
rect 15988 23684 17417 23712
rect 15988 23672 15994 23684
rect 17405 23681 17417 23684
rect 17451 23681 17463 23715
rect 17405 23675 17463 23681
rect 17672 23715 17730 23721
rect 17672 23681 17684 23715
rect 17718 23712 17730 23715
rect 18046 23712 18052 23724
rect 17718 23684 18052 23712
rect 17718 23681 17730 23684
rect 17672 23675 17730 23681
rect 18046 23672 18052 23684
rect 18104 23672 18110 23724
rect 18966 23672 18972 23724
rect 19024 23672 19030 23724
rect 19058 23672 19064 23724
rect 19116 23712 19122 23724
rect 20456 23712 20484 23820
rect 21726 23780 21732 23792
rect 21183 23752 21732 23780
rect 21183 23712 21211 23752
rect 21726 23740 21732 23752
rect 21784 23780 21790 23792
rect 21821 23783 21879 23789
rect 21821 23780 21833 23783
rect 21784 23752 21833 23780
rect 21784 23740 21790 23752
rect 21821 23749 21833 23752
rect 21867 23749 21879 23783
rect 21928 23780 21956 23820
rect 22002 23808 22008 23860
rect 22060 23848 22066 23860
rect 22462 23848 22468 23860
rect 22060 23820 22468 23848
rect 22060 23808 22066 23820
rect 22462 23808 22468 23820
rect 22520 23808 22526 23860
rect 23842 23848 23848 23860
rect 22572 23820 23848 23848
rect 22572 23780 22600 23820
rect 23842 23808 23848 23820
rect 23900 23808 23906 23860
rect 23937 23851 23995 23857
rect 23937 23817 23949 23851
rect 23983 23848 23995 23851
rect 24302 23848 24308 23860
rect 23983 23820 24308 23848
rect 23983 23817 23995 23820
rect 23937 23811 23995 23817
rect 24302 23808 24308 23820
rect 24360 23808 24366 23860
rect 24670 23808 24676 23860
rect 24728 23848 24734 23860
rect 25961 23851 26019 23857
rect 25961 23848 25973 23851
rect 24728 23820 25973 23848
rect 24728 23808 24734 23820
rect 25961 23817 25973 23820
rect 26007 23848 26019 23851
rect 26510 23848 26516 23860
rect 26007 23820 26516 23848
rect 26007 23817 26019 23820
rect 25961 23811 26019 23817
rect 26510 23808 26516 23820
rect 26568 23808 26574 23860
rect 28445 23851 28503 23857
rect 28445 23848 28457 23851
rect 26712 23820 28457 23848
rect 24688 23780 24716 23808
rect 21928 23752 22600 23780
rect 24504 23752 24716 23780
rect 21821 23743 21879 23749
rect 19116 23684 20484 23712
rect 21100 23684 21211 23712
rect 21269 23715 21327 23721
rect 19116 23672 19122 23684
rect 15838 23644 15844 23656
rect 15488 23616 15844 23644
rect 15838 23604 15844 23616
rect 15896 23604 15902 23656
rect 21100 23653 21128 23684
rect 21269 23681 21281 23715
rect 21315 23712 21327 23715
rect 22094 23712 22100 23724
rect 21315 23684 22100 23712
rect 21315 23681 21327 23684
rect 21269 23675 21327 23681
rect 22094 23672 22100 23684
rect 22152 23712 22158 23724
rect 22278 23712 22284 23724
rect 22152 23684 22284 23712
rect 22152 23672 22158 23684
rect 22278 23672 22284 23684
rect 22336 23672 22342 23724
rect 22554 23672 22560 23724
rect 22612 23672 22618 23724
rect 22830 23721 22836 23724
rect 22824 23675 22836 23721
rect 22830 23672 22836 23675
rect 22888 23672 22894 23724
rect 23198 23672 23204 23724
rect 23256 23712 23262 23724
rect 24504 23721 24532 23752
rect 24489 23715 24547 23721
rect 23256 23684 24440 23712
rect 23256 23672 23262 23684
rect 21085 23647 21143 23653
rect 21085 23613 21097 23647
rect 21131 23613 21143 23647
rect 21085 23607 21143 23613
rect 21177 23647 21235 23653
rect 21177 23613 21189 23647
rect 21223 23644 21235 23647
rect 21634 23644 21640 23656
rect 21223 23616 21640 23644
rect 21223 23613 21235 23616
rect 21177 23607 21235 23613
rect 21634 23604 21640 23616
rect 21692 23604 21698 23656
rect 24412 23644 24440 23684
rect 24489 23681 24501 23715
rect 24535 23681 24547 23715
rect 24489 23675 24547 23681
rect 24673 23715 24731 23721
rect 24673 23681 24685 23715
rect 24719 23712 24731 23715
rect 24762 23712 24768 23724
rect 24719 23684 24768 23712
rect 24719 23681 24731 23684
rect 24673 23675 24731 23681
rect 24762 23672 24768 23684
rect 24820 23672 24826 23724
rect 26326 23672 26332 23724
rect 26384 23712 26390 23724
rect 26513 23715 26571 23721
rect 26513 23712 26525 23715
rect 26384 23684 26525 23712
rect 26384 23672 26390 23684
rect 26513 23681 26525 23684
rect 26559 23681 26571 23715
rect 26513 23675 26571 23681
rect 26602 23644 26608 23656
rect 24412 23616 26608 23644
rect 26602 23604 26608 23616
rect 26660 23604 26666 23656
rect 7650 23536 7656 23588
rect 7708 23576 7714 23588
rect 8113 23579 8171 23585
rect 8113 23576 8125 23579
rect 7708 23548 8125 23576
rect 7708 23536 7714 23548
rect 8113 23545 8125 23548
rect 8159 23576 8171 23579
rect 8202 23576 8208 23588
rect 8159 23548 8208 23576
rect 8159 23545 8171 23548
rect 8113 23539 8171 23545
rect 8202 23536 8208 23548
rect 8260 23536 8266 23588
rect 11330 23536 11336 23588
rect 11388 23536 11394 23588
rect 3789 23511 3847 23517
rect 3789 23477 3801 23511
rect 3835 23508 3847 23511
rect 4614 23508 4620 23520
rect 3835 23480 4620 23508
rect 3835 23477 3847 23480
rect 3789 23471 3847 23477
rect 4614 23468 4620 23480
rect 4672 23468 4678 23520
rect 5258 23468 5264 23520
rect 5316 23468 5322 23520
rect 8018 23468 8024 23520
rect 8076 23468 8082 23520
rect 9861 23511 9919 23517
rect 9861 23477 9873 23511
rect 9907 23508 9919 23511
rect 10226 23508 10232 23520
rect 9907 23480 10232 23508
rect 9907 23477 9919 23480
rect 9861 23471 9919 23477
rect 10226 23468 10232 23480
rect 10284 23468 10290 23520
rect 15289 23511 15347 23517
rect 15289 23477 15301 23511
rect 15335 23508 15347 23511
rect 15746 23508 15752 23520
rect 15335 23480 15752 23508
rect 15335 23477 15347 23480
rect 15289 23471 15347 23477
rect 15746 23468 15752 23480
rect 15804 23468 15810 23520
rect 18414 23468 18420 23520
rect 18472 23508 18478 23520
rect 18785 23511 18843 23517
rect 18785 23508 18797 23511
rect 18472 23480 18797 23508
rect 18472 23468 18478 23480
rect 18785 23477 18797 23480
rect 18831 23508 18843 23511
rect 19242 23508 19248 23520
rect 18831 23480 19248 23508
rect 18831 23477 18843 23480
rect 18785 23471 18843 23477
rect 19242 23468 19248 23480
rect 19300 23468 19306 23520
rect 21637 23511 21695 23517
rect 21637 23477 21649 23511
rect 21683 23508 21695 23511
rect 21726 23508 21732 23520
rect 21683 23480 21732 23508
rect 21683 23477 21695 23480
rect 21637 23471 21695 23477
rect 21726 23468 21732 23480
rect 21784 23468 21790 23520
rect 22462 23468 22468 23520
rect 22520 23508 22526 23520
rect 26142 23508 26148 23520
rect 22520 23480 26148 23508
rect 22520 23468 22526 23480
rect 26142 23468 26148 23480
rect 26200 23508 26206 23520
rect 26712 23517 26740 23820
rect 28445 23817 28457 23820
rect 28491 23817 28503 23851
rect 28445 23811 28503 23817
rect 29638 23808 29644 23860
rect 29696 23848 29702 23860
rect 29914 23848 29920 23860
rect 29696 23820 29920 23848
rect 29696 23808 29702 23820
rect 29914 23808 29920 23820
rect 29972 23848 29978 23860
rect 30009 23851 30067 23857
rect 30009 23848 30021 23851
rect 29972 23820 30021 23848
rect 29972 23808 29978 23820
rect 30009 23817 30021 23820
rect 30055 23817 30067 23851
rect 30009 23811 30067 23817
rect 30650 23808 30656 23860
rect 30708 23808 30714 23860
rect 30926 23808 30932 23860
rect 30984 23848 30990 23860
rect 31021 23851 31079 23857
rect 31021 23848 31033 23851
rect 30984 23820 31033 23848
rect 30984 23808 30990 23820
rect 31021 23817 31033 23820
rect 31067 23817 31079 23851
rect 31021 23811 31079 23817
rect 31113 23851 31171 23857
rect 31113 23817 31125 23851
rect 31159 23848 31171 23851
rect 31754 23848 31760 23860
rect 31159 23820 31760 23848
rect 31159 23817 31171 23820
rect 31113 23811 31171 23817
rect 31754 23808 31760 23820
rect 31812 23808 31818 23860
rect 33042 23808 33048 23860
rect 33100 23848 33106 23860
rect 33965 23851 34023 23857
rect 33965 23848 33977 23851
rect 33100 23820 33977 23848
rect 33100 23808 33106 23820
rect 33965 23817 33977 23820
rect 34011 23817 34023 23851
rect 33965 23811 34023 23817
rect 27982 23780 27988 23792
rect 26988 23752 27988 23780
rect 26988 23721 27016 23752
rect 27982 23740 27988 23752
rect 28040 23780 28046 23792
rect 34333 23783 34391 23789
rect 28040 23752 28672 23780
rect 28040 23740 28046 23752
rect 27246 23721 27252 23724
rect 26973 23715 27031 23721
rect 26973 23681 26985 23715
rect 27019 23681 27031 23715
rect 26973 23675 27031 23681
rect 27240 23675 27252 23721
rect 27246 23672 27252 23675
rect 27304 23672 27310 23724
rect 28644 23653 28672 23752
rect 34333 23749 34345 23783
rect 34379 23780 34391 23783
rect 34379 23752 34560 23780
rect 34379 23749 34391 23752
rect 34333 23743 34391 23749
rect 34532 23724 34560 23752
rect 34790 23740 34796 23792
rect 34848 23740 34854 23792
rect 28902 23721 28908 23724
rect 28896 23675 28908 23721
rect 28902 23672 28908 23675
rect 28960 23672 28966 23724
rect 30650 23672 30656 23724
rect 30708 23712 30714 23724
rect 31294 23712 31300 23724
rect 30708 23684 31300 23712
rect 30708 23672 30714 23684
rect 31294 23672 31300 23684
rect 31352 23672 31358 23724
rect 31386 23672 31392 23724
rect 31444 23712 31450 23724
rect 34149 23715 34207 23721
rect 34149 23712 34161 23715
rect 31444 23684 34161 23712
rect 31444 23672 31450 23684
rect 34149 23681 34161 23684
rect 34195 23681 34207 23715
rect 34149 23675 34207 23681
rect 34238 23672 34244 23724
rect 34296 23712 34302 23724
rect 34425 23715 34483 23721
rect 34425 23712 34437 23715
rect 34296 23684 34437 23712
rect 34296 23672 34302 23684
rect 34425 23681 34437 23684
rect 34471 23681 34483 23715
rect 34425 23675 34483 23681
rect 34514 23672 34520 23724
rect 34572 23672 34578 23724
rect 28629 23647 28687 23653
rect 28629 23613 28641 23647
rect 28675 23613 28687 23647
rect 28629 23607 28687 23613
rect 26697 23511 26755 23517
rect 26697 23508 26709 23511
rect 26200 23480 26709 23508
rect 26200 23468 26206 23480
rect 26697 23477 26709 23480
rect 26743 23477 26755 23511
rect 26697 23471 26755 23477
rect 27154 23468 27160 23520
rect 27212 23508 27218 23520
rect 28353 23511 28411 23517
rect 28353 23508 28365 23511
rect 27212 23480 28365 23508
rect 27212 23468 27218 23480
rect 28353 23477 28365 23480
rect 28399 23477 28411 23511
rect 28644 23508 28672 23607
rect 30926 23604 30932 23656
rect 30984 23644 30990 23656
rect 31205 23647 31263 23653
rect 31205 23644 31217 23647
rect 30984 23616 31217 23644
rect 30984 23604 30990 23616
rect 31205 23613 31217 23616
rect 31251 23644 31263 23647
rect 31481 23647 31539 23653
rect 31481 23644 31493 23647
rect 31251 23616 31493 23644
rect 31251 23613 31263 23616
rect 31205 23607 31263 23613
rect 31481 23613 31493 23616
rect 31527 23613 31539 23647
rect 31481 23607 31539 23613
rect 29638 23508 29644 23520
rect 28644 23480 29644 23508
rect 28353 23471 28411 23477
rect 29638 23468 29644 23480
rect 29696 23468 29702 23520
rect 1104 23418 35328 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 35328 23418
rect 1104 23344 35328 23366
rect 5261 23307 5319 23313
rect 5261 23273 5273 23307
rect 5307 23304 5319 23307
rect 5307 23276 8984 23304
rect 5307 23273 5319 23276
rect 5261 23267 5319 23273
rect 4154 23128 4160 23180
rect 4212 23168 4218 23180
rect 4249 23171 4307 23177
rect 4249 23168 4261 23171
rect 4212 23140 4261 23168
rect 4212 23128 4218 23140
rect 4249 23137 4261 23140
rect 4295 23137 4307 23171
rect 4249 23131 4307 23137
rect 4264 23032 4292 23131
rect 5077 23103 5135 23109
rect 5077 23069 5089 23103
rect 5123 23100 5135 23103
rect 5276 23100 5304 23267
rect 6454 23196 6460 23248
rect 6512 23236 6518 23248
rect 6825 23239 6883 23245
rect 6825 23236 6837 23239
rect 6512 23208 6837 23236
rect 6512 23196 6518 23208
rect 6825 23205 6837 23208
rect 6871 23205 6883 23239
rect 6825 23199 6883 23205
rect 5123 23072 5304 23100
rect 5445 23103 5503 23109
rect 5123 23069 5135 23072
rect 5077 23063 5135 23069
rect 5445 23069 5457 23103
rect 5491 23069 5503 23103
rect 5445 23063 5503 23069
rect 5712 23103 5770 23109
rect 5712 23069 5724 23103
rect 5758 23100 5770 23103
rect 6086 23100 6092 23112
rect 5758 23072 6092 23100
rect 5758 23069 5770 23072
rect 5712 23063 5770 23069
rect 4614 23032 4620 23044
rect 4264 23004 4620 23032
rect 4614 22992 4620 23004
rect 4672 23032 4678 23044
rect 5460 23032 5488 23063
rect 6086 23060 6092 23072
rect 6144 23060 6150 23112
rect 4672 23004 5488 23032
rect 6840 23032 6868 23199
rect 7190 23196 7196 23248
rect 7248 23196 7254 23248
rect 8018 23236 8024 23248
rect 7576 23208 8024 23236
rect 7576 23109 7604 23208
rect 8018 23196 8024 23208
rect 8076 23196 8082 23248
rect 8110 23196 8116 23248
rect 8168 23236 8174 23248
rect 8665 23239 8723 23245
rect 8665 23236 8677 23239
rect 8168 23208 8677 23236
rect 8168 23196 8174 23208
rect 8665 23205 8677 23208
rect 8711 23205 8723 23239
rect 8665 23199 8723 23205
rect 7650 23128 7656 23180
rect 7708 23128 7714 23180
rect 7742 23128 7748 23180
rect 7800 23128 7806 23180
rect 8036 23168 8064 23196
rect 8036 23140 8432 23168
rect 7561 23103 7619 23109
rect 7561 23069 7573 23103
rect 7607 23069 7619 23103
rect 7561 23063 7619 23069
rect 7834 23060 7840 23112
rect 7892 23100 7898 23112
rect 8404 23109 8432 23140
rect 8021 23103 8079 23109
rect 8021 23100 8033 23103
rect 7892 23072 8033 23100
rect 7892 23060 7898 23072
rect 8021 23069 8033 23072
rect 8067 23069 8079 23103
rect 8021 23063 8079 23069
rect 8114 23103 8172 23109
rect 8114 23069 8126 23103
rect 8160 23069 8172 23103
rect 8114 23063 8172 23069
rect 8389 23103 8447 23109
rect 8389 23069 8401 23103
rect 8435 23069 8447 23103
rect 8389 23063 8447 23069
rect 8527 23103 8585 23109
rect 8527 23069 8539 23103
rect 8573 23100 8585 23103
rect 8846 23100 8852 23112
rect 8573 23072 8852 23100
rect 8573 23069 8585 23072
rect 8527 23063 8585 23069
rect 8128 23032 8156 23063
rect 8846 23060 8852 23072
rect 8904 23060 8910 23112
rect 8956 23109 8984 23276
rect 10410 23264 10416 23316
rect 10468 23304 10474 23316
rect 10597 23307 10655 23313
rect 10597 23304 10609 23307
rect 10468 23276 10609 23304
rect 10468 23264 10474 23276
rect 10597 23273 10609 23276
rect 10643 23273 10655 23307
rect 10597 23267 10655 23273
rect 10870 23264 10876 23316
rect 10928 23264 10934 23316
rect 11790 23264 11796 23316
rect 11848 23264 11854 23316
rect 11977 23307 12035 23313
rect 11977 23273 11989 23307
rect 12023 23304 12035 23307
rect 12802 23304 12808 23316
rect 12023 23276 12808 23304
rect 12023 23273 12035 23276
rect 11977 23267 12035 23273
rect 10428 23236 10456 23264
rect 10152 23208 10456 23236
rect 9766 23128 9772 23180
rect 9824 23128 9830 23180
rect 8941 23103 8999 23109
rect 8941 23069 8953 23103
rect 8987 23100 8999 23103
rect 10042 23100 10048 23112
rect 8987 23072 10048 23100
rect 8987 23069 8999 23072
rect 8941 23063 8999 23069
rect 10042 23060 10048 23072
rect 10100 23060 10106 23112
rect 10152 23109 10180 23208
rect 10686 23168 10692 23180
rect 10336 23140 10692 23168
rect 10137 23103 10195 23109
rect 10137 23069 10149 23103
rect 10183 23069 10195 23103
rect 10137 23063 10195 23069
rect 10226 23060 10232 23112
rect 10284 23060 10290 23112
rect 6840 23004 8156 23032
rect 8297 23035 8355 23041
rect 4672 22992 4678 23004
rect 8297 23001 8309 23035
rect 8343 23001 8355 23035
rect 8297 22995 8355 23001
rect 8312 22964 8340 22995
rect 8754 22992 8760 23044
rect 8812 23032 8818 23044
rect 10336 23032 10364 23140
rect 10686 23128 10692 23140
rect 10744 23128 10750 23180
rect 10962 23128 10968 23180
rect 11020 23168 11026 23180
rect 11808 23168 11836 23264
rect 11020 23140 11836 23168
rect 11020 23128 11026 23140
rect 10413 23103 10471 23109
rect 10413 23069 10425 23103
rect 10459 23069 10471 23103
rect 10413 23063 10471 23069
rect 10505 23103 10563 23109
rect 10505 23069 10517 23103
rect 10551 23100 10563 23103
rect 10870 23100 10876 23112
rect 10551 23072 10876 23100
rect 10551 23069 10563 23072
rect 10505 23063 10563 23069
rect 8812 23004 10364 23032
rect 10428 23032 10456 23063
rect 10870 23060 10876 23072
rect 10928 23060 10934 23112
rect 11057 23103 11115 23109
rect 11057 23069 11069 23103
rect 11103 23100 11115 23103
rect 11146 23100 11152 23112
rect 11103 23072 11152 23100
rect 11103 23069 11115 23072
rect 11057 23063 11115 23069
rect 11146 23060 11152 23072
rect 11204 23060 11210 23112
rect 11256 23109 11284 23140
rect 11241 23103 11299 23109
rect 11241 23069 11253 23103
rect 11287 23069 11299 23103
rect 11241 23063 11299 23069
rect 11330 23060 11336 23112
rect 11388 23060 11394 23112
rect 11425 23103 11483 23109
rect 11425 23069 11437 23103
rect 11471 23100 11483 23103
rect 11992 23100 12020 23267
rect 12802 23264 12808 23276
rect 12860 23264 12866 23316
rect 14090 23264 14096 23316
rect 14148 23304 14154 23316
rect 17957 23307 18015 23313
rect 17957 23304 17969 23307
rect 14148 23276 17969 23304
rect 14148 23264 14154 23276
rect 17957 23273 17969 23276
rect 18003 23273 18015 23307
rect 17957 23267 18015 23273
rect 16390 23196 16396 23248
rect 16448 23236 16454 23248
rect 16761 23239 16819 23245
rect 16761 23236 16773 23239
rect 16448 23208 16773 23236
rect 16448 23196 16454 23208
rect 16761 23205 16773 23208
rect 16807 23205 16819 23239
rect 16761 23199 16819 23205
rect 17034 23196 17040 23248
rect 17092 23236 17098 23248
rect 17129 23239 17187 23245
rect 17129 23236 17141 23239
rect 17092 23208 17141 23236
rect 17092 23196 17098 23208
rect 17129 23205 17141 23208
rect 17175 23205 17187 23239
rect 17129 23199 17187 23205
rect 16022 23128 16028 23180
rect 16080 23168 16086 23180
rect 16080 23140 17172 23168
rect 16080 23128 16086 23140
rect 12158 23100 12164 23112
rect 11471 23072 12020 23100
rect 12119 23072 12164 23100
rect 11471 23069 11483 23072
rect 11425 23063 11483 23069
rect 12158 23060 12164 23072
rect 12216 23100 12222 23112
rect 14277 23103 14335 23109
rect 14277 23100 14289 23103
rect 12216 23072 14289 23100
rect 12216 23060 12222 23072
rect 14277 23069 14289 23072
rect 14323 23069 14335 23103
rect 14277 23063 14335 23069
rect 14366 23060 14372 23112
rect 14424 23100 14430 23112
rect 15749 23103 15807 23109
rect 15749 23100 15761 23103
rect 14424 23072 15761 23100
rect 14424 23060 14430 23072
rect 15749 23069 15761 23072
rect 15795 23069 15807 23103
rect 15749 23063 15807 23069
rect 15842 23103 15900 23109
rect 15842 23069 15854 23103
rect 15888 23069 15900 23103
rect 15842 23063 15900 23069
rect 12428 23035 12486 23041
rect 10428 23004 10916 23032
rect 8812 22992 8818 23004
rect 8938 22964 8944 22976
rect 8312 22936 8944 22964
rect 8938 22924 8944 22936
rect 8996 22924 9002 22976
rect 9950 22924 9956 22976
rect 10008 22924 10014 22976
rect 10888 22964 10916 23004
rect 12428 23001 12440 23035
rect 12474 23032 12486 23035
rect 12710 23032 12716 23044
rect 12474 23004 12716 23032
rect 12474 23001 12486 23004
rect 12428 22995 12486 23001
rect 12710 22992 12716 23004
rect 12768 22992 12774 23044
rect 14544 23035 14602 23041
rect 14544 23001 14556 23035
rect 14590 23032 14602 23035
rect 14826 23032 14832 23044
rect 14590 23004 14832 23032
rect 14590 23001 14602 23004
rect 14544 22995 14602 23001
rect 14826 22992 14832 23004
rect 14884 22992 14890 23044
rect 15856 23032 15884 23063
rect 16206 23060 16212 23112
rect 16264 23109 16270 23112
rect 16264 23100 16272 23109
rect 16577 23103 16635 23109
rect 16577 23100 16589 23103
rect 16264 23072 16589 23100
rect 16264 23063 16272 23072
rect 16577 23069 16589 23072
rect 16623 23100 16635 23103
rect 16945 23103 17003 23109
rect 16945 23100 16957 23103
rect 16623 23072 16957 23100
rect 16623 23069 16635 23072
rect 16577 23063 16635 23069
rect 16945 23069 16957 23072
rect 16991 23069 17003 23103
rect 16945 23063 17003 23069
rect 16264 23060 16270 23063
rect 15672 23004 15884 23032
rect 16025 23035 16083 23041
rect 15672 22976 15700 23004
rect 16025 23001 16037 23035
rect 16071 23001 16083 23035
rect 16025 22995 16083 23001
rect 11609 22967 11667 22973
rect 11609 22964 11621 22967
rect 10888 22936 11621 22964
rect 11609 22933 11621 22936
rect 11655 22933 11667 22967
rect 11609 22927 11667 22933
rect 13538 22924 13544 22976
rect 13596 22924 13602 22976
rect 15654 22924 15660 22976
rect 15712 22924 15718 22976
rect 16040 22964 16068 22995
rect 16114 22992 16120 23044
rect 16172 22992 16178 23044
rect 17034 23032 17040 23044
rect 16215 23004 17040 23032
rect 16215 22964 16243 23004
rect 17034 22992 17040 23004
rect 17092 22992 17098 23044
rect 17144 23032 17172 23140
rect 17972 23100 18000 23267
rect 22830 23264 22836 23316
rect 22888 23304 22894 23316
rect 23017 23307 23075 23313
rect 23017 23304 23029 23307
rect 22888 23276 23029 23304
rect 22888 23264 22894 23276
rect 23017 23273 23029 23276
rect 23063 23273 23075 23307
rect 23017 23267 23075 23273
rect 23308 23276 25728 23304
rect 22738 23196 22744 23248
rect 22796 23236 22802 23248
rect 23308 23236 23336 23276
rect 22796 23208 23336 23236
rect 22796 23196 22802 23208
rect 23382 23196 23388 23248
rect 23440 23196 23446 23248
rect 25700 23236 25728 23276
rect 25774 23264 25780 23316
rect 25832 23264 25838 23316
rect 26418 23264 26424 23316
rect 26476 23264 26482 23316
rect 26510 23264 26516 23316
rect 26568 23264 26574 23316
rect 27157 23307 27215 23313
rect 27157 23273 27169 23307
rect 27203 23304 27215 23307
rect 27246 23304 27252 23316
rect 27203 23276 27252 23304
rect 27203 23273 27215 23276
rect 27157 23267 27215 23273
rect 27246 23264 27252 23276
rect 27304 23264 27310 23316
rect 27706 23264 27712 23316
rect 27764 23304 27770 23316
rect 28166 23304 28172 23316
rect 27764 23276 28172 23304
rect 27764 23264 27770 23276
rect 28166 23264 28172 23276
rect 28224 23264 28230 23316
rect 28902 23264 28908 23316
rect 28960 23304 28966 23316
rect 29549 23307 29607 23313
rect 29549 23304 29561 23307
rect 28960 23276 29561 23304
rect 28960 23264 28966 23276
rect 29549 23273 29561 23276
rect 29595 23273 29607 23307
rect 29549 23267 29607 23273
rect 26973 23239 27031 23245
rect 26973 23236 26985 23239
rect 25700 23208 26985 23236
rect 26973 23205 26985 23208
rect 27019 23205 27031 23239
rect 26973 23199 27031 23205
rect 18966 23128 18972 23180
rect 19024 23168 19030 23180
rect 23400 23168 23428 23196
rect 23477 23171 23535 23177
rect 23477 23168 23489 23171
rect 19024 23140 19288 23168
rect 23400 23140 23489 23168
rect 19024 23128 19030 23140
rect 19260 23109 19288 23140
rect 23477 23137 23489 23140
rect 23523 23137 23535 23171
rect 23477 23131 23535 23137
rect 23566 23128 23572 23180
rect 23624 23168 23630 23180
rect 23845 23171 23903 23177
rect 23845 23168 23857 23171
rect 23624 23140 23857 23168
rect 23624 23128 23630 23140
rect 23845 23137 23857 23140
rect 23891 23137 23903 23171
rect 23845 23131 23903 23137
rect 21726 23109 21732 23112
rect 18141 23103 18199 23109
rect 18141 23100 18153 23103
rect 17972 23072 18153 23100
rect 18141 23069 18153 23072
rect 18187 23069 18199 23103
rect 18141 23063 18199 23069
rect 19245 23103 19303 23109
rect 19245 23069 19257 23103
rect 19291 23100 19303 23103
rect 21453 23103 21511 23109
rect 21453 23100 21465 23103
rect 19291 23072 21465 23100
rect 19291 23069 19303 23072
rect 19245 23063 19303 23069
rect 21453 23069 21465 23072
rect 21499 23069 21511 23103
rect 21720 23100 21732 23109
rect 21687 23072 21732 23100
rect 21453 23063 21511 23069
rect 21720 23063 21732 23072
rect 21726 23060 21732 23063
rect 21784 23060 21790 23112
rect 23385 23103 23443 23109
rect 23385 23069 23397 23103
rect 23431 23100 23443 23103
rect 24302 23100 24308 23112
rect 23431 23072 24308 23100
rect 23431 23069 23443 23072
rect 23385 23063 23443 23069
rect 24302 23060 24308 23072
rect 24360 23060 24366 23112
rect 24397 23103 24455 23109
rect 24397 23069 24409 23103
rect 24443 23100 24455 23103
rect 24946 23100 24952 23112
rect 24443 23072 24952 23100
rect 24443 23069 24455 23072
rect 24397 23063 24455 23069
rect 24946 23060 24952 23072
rect 25004 23060 25010 23112
rect 18230 23032 18236 23044
rect 17144 23004 18236 23032
rect 18230 22992 18236 23004
rect 18288 23032 18294 23044
rect 24664 23035 24722 23041
rect 18288 23004 24624 23032
rect 18288 22992 18294 23004
rect 16040 22936 16243 22964
rect 16393 22967 16451 22973
rect 16393 22933 16405 22967
rect 16439 22964 16451 22967
rect 16758 22964 16764 22976
rect 16439 22936 16764 22964
rect 16439 22933 16451 22936
rect 16393 22927 16451 22933
rect 16758 22924 16764 22936
rect 16816 22924 16822 22976
rect 22278 22924 22284 22976
rect 22336 22964 22342 22976
rect 22833 22967 22891 22973
rect 22833 22964 22845 22967
rect 22336 22936 22845 22964
rect 22336 22924 22342 22936
rect 22833 22933 22845 22936
rect 22879 22933 22891 22967
rect 22833 22927 22891 22933
rect 23474 22924 23480 22976
rect 23532 22964 23538 22976
rect 23934 22964 23940 22976
rect 23532 22936 23940 22964
rect 23532 22924 23538 22936
rect 23934 22924 23940 22936
rect 23992 22964 23998 22976
rect 24029 22967 24087 22973
rect 24029 22964 24041 22967
rect 23992 22936 24041 22964
rect 23992 22924 23998 22936
rect 24029 22933 24041 22936
rect 24075 22933 24087 22967
rect 24596 22964 24624 23004
rect 24664 23001 24676 23035
rect 24710 23032 24722 23035
rect 24854 23032 24860 23044
rect 24710 23004 24860 23032
rect 24710 23001 24722 23004
rect 24664 22995 24722 23001
rect 24854 22992 24860 23004
rect 24912 22992 24918 23044
rect 26988 23032 27016 23199
rect 27522 23196 27528 23248
rect 27580 23196 27586 23248
rect 27540 23168 27568 23196
rect 27709 23171 27767 23177
rect 27709 23168 27721 23171
rect 27540 23140 27721 23168
rect 27709 23137 27721 23140
rect 27755 23137 27767 23171
rect 27709 23131 27767 23137
rect 29454 23128 29460 23180
rect 29512 23168 29518 23180
rect 30101 23171 30159 23177
rect 30101 23168 30113 23171
rect 29512 23140 30113 23168
rect 29512 23128 29518 23140
rect 30101 23137 30113 23140
rect 30147 23168 30159 23171
rect 30377 23171 30435 23177
rect 30377 23168 30389 23171
rect 30147 23140 30389 23168
rect 30147 23137 30159 23140
rect 30101 23131 30159 23137
rect 30377 23137 30389 23140
rect 30423 23168 30435 23171
rect 30742 23168 30748 23180
rect 30423 23140 30748 23168
rect 30423 23137 30435 23140
rect 30377 23131 30435 23137
rect 30742 23128 30748 23140
rect 30800 23128 30806 23180
rect 27154 23060 27160 23112
rect 27212 23100 27218 23112
rect 27525 23103 27583 23109
rect 27525 23100 27537 23103
rect 27212 23072 27537 23100
rect 27212 23060 27218 23072
rect 27525 23069 27537 23072
rect 27571 23069 27583 23103
rect 27525 23063 27583 23069
rect 29365 23103 29423 23109
rect 29365 23069 29377 23103
rect 29411 23100 29423 23103
rect 29546 23100 29552 23112
rect 29411 23072 29552 23100
rect 29411 23069 29423 23072
rect 29365 23063 29423 23069
rect 29546 23060 29552 23072
rect 29604 23060 29610 23112
rect 29914 23060 29920 23112
rect 29972 23060 29978 23112
rect 27617 23035 27675 23041
rect 27617 23032 27629 23035
rect 26988 23004 27629 23032
rect 27617 23001 27629 23004
rect 27663 23032 27675 23035
rect 28997 23035 29055 23041
rect 28997 23032 29009 23035
rect 27663 23004 29009 23032
rect 27663 23001 27675 23004
rect 27617 22995 27675 23001
rect 28997 23001 29009 23004
rect 29043 23032 29055 23035
rect 30009 23035 30067 23041
rect 30009 23032 30021 23035
rect 29043 23004 30021 23032
rect 29043 23001 29055 23004
rect 28997 22995 29055 23001
rect 30009 23001 30021 23004
rect 30055 23001 30067 23035
rect 30009 22995 30067 23001
rect 26234 22964 26240 22976
rect 24596 22936 26240 22964
rect 24029 22927 24087 22933
rect 26234 22924 26240 22936
rect 26292 22964 26298 22976
rect 26697 22967 26755 22973
rect 26697 22964 26709 22967
rect 26292 22936 26709 22964
rect 26292 22924 26298 22936
rect 26697 22933 26709 22936
rect 26743 22933 26755 22967
rect 26697 22927 26755 22933
rect 29181 22967 29239 22973
rect 29181 22933 29193 22967
rect 29227 22964 29239 22967
rect 29270 22964 29276 22976
rect 29227 22936 29276 22964
rect 29227 22933 29239 22936
rect 29181 22927 29239 22933
rect 29270 22924 29276 22936
rect 29328 22924 29334 22976
rect 1104 22874 35328 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35328 22874
rect 1104 22800 35328 22822
rect 3786 22720 3792 22772
rect 3844 22720 3850 22772
rect 4249 22763 4307 22769
rect 4249 22729 4261 22763
rect 4295 22760 4307 22763
rect 4522 22760 4528 22772
rect 4295 22732 4528 22760
rect 4295 22729 4307 22732
rect 4249 22723 4307 22729
rect 4522 22720 4528 22732
rect 4580 22720 4586 22772
rect 4706 22720 4712 22772
rect 4764 22760 4770 22772
rect 5445 22763 5503 22769
rect 5445 22760 5457 22763
rect 4764 22732 5457 22760
rect 4764 22720 4770 22732
rect 1302 22584 1308 22636
rect 1360 22624 1366 22636
rect 1489 22627 1547 22633
rect 1489 22624 1501 22627
rect 1360 22596 1501 22624
rect 1360 22584 1366 22596
rect 1489 22593 1501 22596
rect 1535 22624 1547 22627
rect 1949 22627 2007 22633
rect 1949 22624 1961 22627
rect 1535 22596 1961 22624
rect 1535 22593 1547 22596
rect 1489 22587 1547 22593
rect 1949 22593 1961 22596
rect 1995 22593 2007 22627
rect 1949 22587 2007 22593
rect 4157 22627 4215 22633
rect 4157 22593 4169 22627
rect 4203 22624 4215 22627
rect 4540 22624 4568 22720
rect 5000 22701 5028 22732
rect 5445 22729 5457 22732
rect 5491 22729 5503 22763
rect 5445 22723 5503 22729
rect 7742 22720 7748 22772
rect 7800 22760 7806 22772
rect 8573 22763 8631 22769
rect 8573 22760 8585 22763
rect 7800 22732 8585 22760
rect 7800 22720 7806 22732
rect 8573 22729 8585 22732
rect 8619 22760 8631 22763
rect 8754 22760 8760 22772
rect 8619 22732 8760 22760
rect 8619 22729 8631 22732
rect 8573 22723 8631 22729
rect 8754 22720 8760 22732
rect 8812 22720 8818 22772
rect 8846 22720 8852 22772
rect 8904 22720 8910 22772
rect 9030 22720 9036 22772
rect 9088 22720 9094 22772
rect 9401 22763 9459 22769
rect 9401 22729 9413 22763
rect 9447 22760 9459 22763
rect 10226 22760 10232 22772
rect 9447 22732 10232 22760
rect 9447 22729 9459 22732
rect 9401 22723 9459 22729
rect 10226 22720 10232 22732
rect 10284 22720 10290 22772
rect 12710 22720 12716 22772
rect 12768 22720 12774 22772
rect 14093 22763 14151 22769
rect 14093 22729 14105 22763
rect 14139 22760 14151 22763
rect 14366 22760 14372 22772
rect 14139 22732 14372 22760
rect 14139 22729 14151 22732
rect 14093 22723 14151 22729
rect 14366 22720 14372 22732
rect 14424 22720 14430 22772
rect 14826 22720 14832 22772
rect 14884 22720 14890 22772
rect 15197 22763 15255 22769
rect 15197 22729 15209 22763
rect 15243 22760 15255 22763
rect 15654 22760 15660 22772
rect 15243 22732 15660 22760
rect 15243 22729 15255 22732
rect 15197 22723 15255 22729
rect 15654 22720 15660 22732
rect 15712 22720 15718 22772
rect 17497 22763 17555 22769
rect 17497 22760 17509 22763
rect 16684 22732 17509 22760
rect 4985 22695 5043 22701
rect 4985 22661 4997 22695
rect 5031 22661 5043 22695
rect 4985 22655 5043 22661
rect 5077 22695 5135 22701
rect 5077 22661 5089 22695
rect 5123 22692 5135 22695
rect 5258 22692 5264 22704
rect 5123 22664 5264 22692
rect 5123 22661 5135 22664
rect 5077 22655 5135 22661
rect 5258 22652 5264 22664
rect 5316 22652 5322 22704
rect 7929 22695 7987 22701
rect 7929 22661 7941 22695
rect 7975 22692 7987 22695
rect 9950 22692 9956 22704
rect 7975 22664 9956 22692
rect 7975 22661 7987 22664
rect 7929 22655 7987 22661
rect 9950 22652 9956 22664
rect 10008 22652 10014 22704
rect 10502 22652 10508 22704
rect 10560 22692 10566 22704
rect 13725 22695 13783 22701
rect 13725 22692 13737 22695
rect 10560 22664 13737 22692
rect 10560 22652 10566 22664
rect 13725 22661 13737 22664
rect 13771 22692 13783 22695
rect 14185 22695 14243 22701
rect 14185 22692 14197 22695
rect 13771 22664 14197 22692
rect 13771 22661 13783 22664
rect 13725 22655 13783 22661
rect 14185 22661 14197 22664
rect 14231 22661 14243 22695
rect 14185 22655 14243 22661
rect 4801 22627 4859 22633
rect 4801 22624 4813 22627
rect 4203 22596 4476 22624
rect 4540 22596 4813 22624
rect 4203 22593 4215 22596
rect 4157 22587 4215 22593
rect 4341 22559 4399 22565
rect 4341 22525 4353 22559
rect 4387 22525 4399 22559
rect 4448 22556 4476 22596
rect 4801 22593 4813 22596
rect 4847 22593 4859 22627
rect 4801 22587 4859 22593
rect 5169 22627 5227 22633
rect 5169 22593 5181 22627
rect 5215 22624 5227 22627
rect 5718 22624 5724 22636
rect 5215 22596 5724 22624
rect 5215 22593 5227 22596
rect 5169 22587 5227 22593
rect 5718 22584 5724 22596
rect 5776 22584 5782 22636
rect 8110 22584 8116 22636
rect 8168 22624 8174 22636
rect 8205 22627 8263 22633
rect 8205 22624 8217 22627
rect 8168 22596 8217 22624
rect 8168 22584 8174 22596
rect 8205 22593 8217 22596
rect 8251 22593 8263 22627
rect 8205 22587 8263 22593
rect 8294 22584 8300 22636
rect 8352 22624 8358 22636
rect 9493 22627 9551 22633
rect 9493 22624 9505 22627
rect 8352 22596 9505 22624
rect 8352 22584 8358 22596
rect 9493 22593 9505 22596
rect 9539 22593 9551 22627
rect 9493 22587 9551 22593
rect 9766 22584 9772 22636
rect 9824 22624 9830 22636
rect 9861 22627 9919 22633
rect 9861 22624 9873 22627
rect 9824 22596 9873 22624
rect 9824 22584 9830 22596
rect 9861 22593 9873 22596
rect 9907 22593 9919 22627
rect 9861 22587 9919 22593
rect 10128 22627 10186 22633
rect 10128 22593 10140 22627
rect 10174 22624 10186 22627
rect 10410 22624 10416 22636
rect 10174 22596 10416 22624
rect 10174 22593 10186 22596
rect 10128 22587 10186 22593
rect 10410 22584 10416 22596
rect 10468 22584 10474 22636
rect 13081 22627 13139 22633
rect 13081 22593 13093 22627
rect 13127 22624 13139 22627
rect 13538 22624 13544 22636
rect 13127 22596 13544 22624
rect 13127 22593 13139 22596
rect 13081 22587 13139 22593
rect 13538 22584 13544 22596
rect 13596 22584 13602 22636
rect 13814 22584 13820 22636
rect 13872 22584 13878 22636
rect 13909 22627 13967 22633
rect 13909 22593 13921 22627
rect 13955 22624 13967 22627
rect 14369 22627 14427 22633
rect 14369 22624 14381 22627
rect 13955 22596 14381 22624
rect 13955 22593 13967 22596
rect 13909 22587 13967 22593
rect 14369 22593 14381 22596
rect 14415 22624 14427 22627
rect 16022 22624 16028 22636
rect 14415 22596 16028 22624
rect 14415 22593 14427 22596
rect 14369 22587 14427 22593
rect 16022 22584 16028 22596
rect 16080 22584 16086 22636
rect 16482 22584 16488 22636
rect 16540 22584 16546 22636
rect 16684 22633 16712 22732
rect 17497 22729 17509 22732
rect 17543 22760 17555 22763
rect 17770 22760 17776 22772
rect 17543 22732 17776 22760
rect 17543 22729 17555 22732
rect 17497 22723 17555 22729
rect 17770 22720 17776 22732
rect 17828 22720 17834 22772
rect 17957 22763 18015 22769
rect 17957 22729 17969 22763
rect 18003 22760 18015 22763
rect 18046 22760 18052 22772
rect 18003 22732 18052 22760
rect 18003 22729 18015 22732
rect 17957 22723 18015 22729
rect 18046 22720 18052 22732
rect 18104 22720 18110 22772
rect 18322 22720 18328 22772
rect 18380 22720 18386 22772
rect 18414 22720 18420 22772
rect 18472 22720 18478 22772
rect 19334 22720 19340 22772
rect 19392 22720 19398 22772
rect 19518 22720 19524 22772
rect 19576 22760 19582 22772
rect 19705 22763 19763 22769
rect 19705 22760 19717 22763
rect 19576 22732 19717 22760
rect 19576 22720 19582 22732
rect 19705 22729 19717 22732
rect 19751 22729 19763 22763
rect 21910 22760 21916 22772
rect 19705 22723 19763 22729
rect 20548 22732 21916 22760
rect 16758 22652 16764 22704
rect 16816 22692 16822 22704
rect 18340 22692 18368 22720
rect 19797 22695 19855 22701
rect 19797 22692 19809 22695
rect 16816 22664 16896 22692
rect 18340 22664 19809 22692
rect 16816 22652 16822 22664
rect 16868 22633 16896 22664
rect 19797 22661 19809 22664
rect 19843 22661 19855 22695
rect 19797 22655 19855 22661
rect 16669 22627 16727 22633
rect 16669 22593 16681 22627
rect 16715 22593 16727 22627
rect 16669 22587 16727 22593
rect 16853 22627 16911 22633
rect 16853 22593 16865 22627
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 17218 22584 17224 22636
rect 17276 22584 17282 22636
rect 20548 22624 20576 22732
rect 21910 22720 21916 22732
rect 21968 22720 21974 22772
rect 25958 22720 25964 22772
rect 26016 22760 26022 22772
rect 26329 22763 26387 22769
rect 26329 22760 26341 22763
rect 26016 22732 26341 22760
rect 26016 22720 26022 22732
rect 26329 22729 26341 22732
rect 26375 22729 26387 22763
rect 26329 22723 26387 22729
rect 26602 22720 26608 22772
rect 26660 22760 26666 22772
rect 27246 22760 27252 22772
rect 26660 22732 27252 22760
rect 26660 22720 26666 22732
rect 27246 22720 27252 22732
rect 27304 22760 27310 22772
rect 27801 22763 27859 22769
rect 27801 22760 27813 22763
rect 27304 22732 27813 22760
rect 27304 22720 27310 22732
rect 27801 22729 27813 22732
rect 27847 22729 27859 22763
rect 27801 22723 27859 22729
rect 29089 22763 29147 22769
rect 29089 22729 29101 22763
rect 29135 22760 29147 22763
rect 29270 22760 29276 22772
rect 29135 22732 29276 22760
rect 29135 22729 29147 22732
rect 29089 22723 29147 22729
rect 20993 22695 21051 22701
rect 20993 22692 21005 22695
rect 20640 22664 21005 22692
rect 20640 22633 20668 22664
rect 20993 22661 21005 22664
rect 21039 22692 21051 22695
rect 21039 22664 27752 22692
rect 21039 22661 21051 22664
rect 20993 22655 21051 22661
rect 18616 22596 20576 22624
rect 20625 22627 20683 22633
rect 4706 22556 4712 22568
rect 4448 22528 4712 22556
rect 4341 22519 4399 22525
rect 1673 22491 1731 22497
rect 1673 22457 1685 22491
rect 1719 22488 1731 22491
rect 1854 22488 1860 22500
rect 1719 22460 1860 22488
rect 1719 22457 1731 22460
rect 1673 22451 1731 22457
rect 1854 22448 1860 22460
rect 1912 22448 1918 22500
rect 4356 22420 4384 22519
rect 4706 22516 4712 22528
rect 4764 22556 4770 22568
rect 5442 22556 5448 22568
rect 4764 22528 5448 22556
rect 4764 22516 4770 22528
rect 5442 22516 5448 22528
rect 5500 22516 5506 22568
rect 5534 22516 5540 22568
rect 5592 22556 5598 22568
rect 8021 22559 8079 22565
rect 8021 22556 8033 22559
rect 5592 22528 8033 22556
rect 5592 22516 5598 22528
rect 8021 22525 8033 22528
rect 8067 22525 8079 22559
rect 8021 22519 8079 22525
rect 9585 22559 9643 22565
rect 9585 22525 9597 22559
rect 9631 22556 9643 22559
rect 9674 22556 9680 22568
rect 9631 22528 9680 22556
rect 9631 22525 9643 22528
rect 9585 22519 9643 22525
rect 9674 22516 9680 22528
rect 9732 22516 9738 22568
rect 13170 22516 13176 22568
rect 13228 22516 13234 22568
rect 13262 22516 13268 22568
rect 13320 22516 13326 22568
rect 13446 22516 13452 22568
rect 13504 22556 13510 22568
rect 15289 22559 15347 22565
rect 15289 22556 15301 22559
rect 13504 22528 15301 22556
rect 13504 22516 13510 22528
rect 15289 22525 15301 22528
rect 15335 22525 15347 22559
rect 15289 22519 15347 22525
rect 15473 22559 15531 22565
rect 15473 22525 15485 22559
rect 15519 22556 15531 22559
rect 15746 22556 15752 22568
rect 15519 22528 15752 22556
rect 15519 22525 15531 22528
rect 15473 22519 15531 22525
rect 15746 22516 15752 22528
rect 15804 22516 15810 22568
rect 16206 22516 16212 22568
rect 16264 22516 16270 22568
rect 16500 22556 16528 22584
rect 16758 22556 16764 22568
rect 16500 22528 16764 22556
rect 16758 22516 16764 22528
rect 16816 22516 16822 22568
rect 16945 22559 17003 22565
rect 16945 22525 16957 22559
rect 16991 22525 17003 22559
rect 16945 22519 17003 22525
rect 17037 22559 17095 22565
rect 17037 22525 17049 22559
rect 17083 22556 17095 22559
rect 17681 22559 17739 22565
rect 17681 22556 17693 22559
rect 17083 22528 17693 22556
rect 17083 22525 17095 22528
rect 17037 22519 17095 22525
rect 17681 22525 17693 22528
rect 17727 22556 17739 22559
rect 17862 22556 17868 22568
rect 17727 22528 17868 22556
rect 17727 22525 17739 22528
rect 17681 22519 17739 22525
rect 5353 22491 5411 22497
rect 5353 22457 5365 22491
rect 5399 22488 5411 22491
rect 8389 22491 8447 22497
rect 5399 22460 7972 22488
rect 5399 22457 5411 22460
rect 5353 22451 5411 22457
rect 4709 22423 4767 22429
rect 4709 22420 4721 22423
rect 4356 22392 4721 22420
rect 4709 22389 4721 22392
rect 4755 22420 4767 22423
rect 4798 22420 4804 22432
rect 4755 22392 4804 22420
rect 4755 22389 4767 22392
rect 4709 22383 4767 22389
rect 4798 22380 4804 22392
rect 4856 22420 4862 22432
rect 5258 22420 5264 22432
rect 4856 22392 5264 22420
rect 4856 22380 4862 22392
rect 5258 22380 5264 22392
rect 5316 22380 5322 22432
rect 5718 22380 5724 22432
rect 5776 22380 5782 22432
rect 7944 22429 7972 22460
rect 8389 22457 8401 22491
rect 8435 22488 8447 22491
rect 16960 22488 16988 22519
rect 17862 22516 17868 22528
rect 17920 22516 17926 22568
rect 18616 22565 18644 22596
rect 20625 22593 20637 22627
rect 20671 22593 20683 22627
rect 20625 22587 20683 22593
rect 21821 22627 21879 22633
rect 21821 22593 21833 22627
rect 21867 22624 21879 22627
rect 23750 22624 23756 22636
rect 21867 22596 23756 22624
rect 21867 22593 21879 22596
rect 21821 22587 21879 22593
rect 18601 22559 18659 22565
rect 18601 22525 18613 22559
rect 18647 22525 18659 22559
rect 18601 22519 18659 22525
rect 19889 22559 19947 22565
rect 19889 22525 19901 22559
rect 19935 22525 19947 22559
rect 19889 22519 19947 22525
rect 19904 22488 19932 22519
rect 20438 22516 20444 22568
rect 20496 22556 20502 22568
rect 21836 22556 21864 22587
rect 23750 22584 23756 22596
rect 23808 22584 23814 22636
rect 24765 22627 24823 22633
rect 24765 22593 24777 22627
rect 24811 22624 24823 22627
rect 24946 22624 24952 22636
rect 24811 22596 24952 22624
rect 24811 22593 24823 22596
rect 24765 22587 24823 22593
rect 24946 22584 24952 22596
rect 25004 22584 25010 22636
rect 25216 22627 25274 22633
rect 25216 22593 25228 22627
rect 25262 22624 25274 22627
rect 25498 22624 25504 22636
rect 25262 22596 25504 22624
rect 25262 22593 25274 22596
rect 25216 22587 25274 22593
rect 25498 22584 25504 22596
rect 25556 22584 25562 22636
rect 26326 22584 26332 22636
rect 26384 22624 26390 22636
rect 27065 22627 27123 22633
rect 27065 22624 27077 22627
rect 26384 22596 27077 22624
rect 26384 22584 26390 22596
rect 27065 22593 27077 22596
rect 27111 22624 27123 22627
rect 27154 22624 27160 22636
rect 27111 22596 27160 22624
rect 27111 22593 27123 22596
rect 27065 22587 27123 22593
rect 27154 22584 27160 22596
rect 27212 22584 27218 22636
rect 20496 22528 21864 22556
rect 20496 22516 20502 22528
rect 22186 22516 22192 22568
rect 22244 22556 22250 22568
rect 22830 22556 22836 22568
rect 22244 22528 22836 22556
rect 22244 22516 22250 22528
rect 22830 22516 22836 22528
rect 22888 22516 22894 22568
rect 27724 22556 27752 22664
rect 27816 22624 27844 22723
rect 29270 22720 29276 22732
rect 29328 22720 29334 22772
rect 29178 22652 29184 22704
rect 29236 22692 29242 22704
rect 34333 22695 34391 22701
rect 29236 22664 34192 22692
rect 29236 22652 29242 22664
rect 27985 22627 28043 22633
rect 27985 22624 27997 22627
rect 27816 22596 27997 22624
rect 27985 22593 27997 22596
rect 28031 22593 28043 22627
rect 27985 22587 28043 22593
rect 28166 22584 28172 22636
rect 28224 22624 28230 22636
rect 28261 22627 28319 22633
rect 28261 22624 28273 22627
rect 28224 22596 28273 22624
rect 28224 22584 28230 22596
rect 28261 22593 28273 22596
rect 28307 22593 28319 22627
rect 28261 22587 28319 22593
rect 28905 22627 28963 22633
rect 28905 22593 28917 22627
rect 28951 22624 28963 22627
rect 29546 22624 29552 22636
rect 28951 22596 29552 22624
rect 28951 22593 28963 22596
rect 28905 22587 28963 22593
rect 29546 22584 29552 22596
rect 29604 22624 29610 22636
rect 30098 22624 30104 22636
rect 29604 22596 30104 22624
rect 29604 22584 29610 22596
rect 30098 22584 30104 22596
rect 30156 22584 30162 22636
rect 30558 22584 30564 22636
rect 30616 22633 30622 22636
rect 30616 22587 30628 22633
rect 30837 22627 30895 22633
rect 30837 22593 30849 22627
rect 30883 22624 30895 22627
rect 31386 22624 31392 22636
rect 30883 22596 31392 22624
rect 30883 22593 30895 22596
rect 30837 22587 30895 22593
rect 30616 22584 30622 22587
rect 31386 22584 31392 22596
rect 31444 22584 31450 22636
rect 34164 22633 34192 22664
rect 34333 22661 34345 22695
rect 34379 22692 34391 22695
rect 34379 22664 34560 22692
rect 34379 22661 34391 22664
rect 34333 22655 34391 22661
rect 34532 22636 34560 22664
rect 34149 22627 34207 22633
rect 34149 22593 34161 22627
rect 34195 22593 34207 22627
rect 34149 22587 34207 22593
rect 34238 22584 34244 22636
rect 34296 22624 34302 22636
rect 34425 22627 34483 22633
rect 34425 22624 34437 22627
rect 34296 22596 34437 22624
rect 34296 22584 34302 22596
rect 34425 22593 34437 22596
rect 34471 22593 34483 22627
rect 34425 22587 34483 22593
rect 34514 22584 34520 22636
rect 34572 22584 34578 22636
rect 29730 22556 29736 22568
rect 27724 22528 29736 22556
rect 29730 22516 29736 22528
rect 29788 22516 29794 22568
rect 34790 22516 34796 22568
rect 34848 22516 34854 22568
rect 20165 22491 20223 22497
rect 20165 22488 20177 22491
rect 8435 22460 9674 22488
rect 8435 22457 8447 22460
rect 8389 22451 8447 22457
rect 7929 22423 7987 22429
rect 7929 22389 7941 22423
rect 7975 22389 7987 22423
rect 7929 22383 7987 22389
rect 8757 22423 8815 22429
rect 8757 22389 8769 22423
rect 8803 22420 8815 22423
rect 8938 22420 8944 22432
rect 8803 22392 8944 22420
rect 8803 22389 8815 22392
rect 8757 22383 8815 22389
rect 8938 22380 8944 22392
rect 8996 22380 9002 22432
rect 9646 22420 9674 22460
rect 10796 22460 16988 22488
rect 17052 22460 20177 22488
rect 10796 22420 10824 22460
rect 9646 22392 10824 22420
rect 11238 22380 11244 22432
rect 11296 22380 11302 22432
rect 12250 22380 12256 22432
rect 12308 22420 12314 22432
rect 17052 22420 17080 22460
rect 20165 22457 20177 22460
rect 20211 22488 20223 22491
rect 23566 22488 23572 22500
rect 20211 22460 23572 22488
rect 20211 22457 20223 22460
rect 20165 22451 20223 22457
rect 23566 22448 23572 22460
rect 23624 22448 23630 22500
rect 29086 22448 29092 22500
rect 29144 22488 29150 22500
rect 29144 22460 29592 22488
rect 29144 22448 29150 22460
rect 12308 22392 17080 22420
rect 12308 22380 12314 22392
rect 17402 22380 17408 22432
rect 17460 22380 17466 22432
rect 19153 22423 19211 22429
rect 19153 22389 19165 22423
rect 19199 22420 19211 22423
rect 19242 22420 19248 22432
rect 19199 22392 19248 22420
rect 19199 22389 19211 22392
rect 19153 22383 19211 22389
rect 19242 22380 19248 22392
rect 19300 22380 19306 22432
rect 20441 22423 20499 22429
rect 20441 22389 20453 22423
rect 20487 22420 20499 22423
rect 20717 22423 20775 22429
rect 20717 22420 20729 22423
rect 20487 22392 20729 22420
rect 20487 22389 20499 22392
rect 20441 22383 20499 22389
rect 20717 22389 20729 22392
rect 20763 22420 20775 22423
rect 20806 22420 20812 22432
rect 20763 22392 20812 22420
rect 20763 22389 20775 22392
rect 20717 22383 20775 22389
rect 20806 22380 20812 22392
rect 20864 22380 20870 22432
rect 22005 22423 22063 22429
rect 22005 22389 22017 22423
rect 22051 22420 22063 22423
rect 22738 22420 22744 22432
rect 22051 22392 22744 22420
rect 22051 22389 22063 22392
rect 22005 22383 22063 22389
rect 22738 22380 22744 22392
rect 22796 22380 22802 22432
rect 29270 22380 29276 22432
rect 29328 22380 29334 22432
rect 29454 22380 29460 22432
rect 29512 22380 29518 22432
rect 29564 22420 29592 22460
rect 29730 22420 29736 22432
rect 29564 22392 29736 22420
rect 29730 22380 29736 22392
rect 29788 22380 29794 22432
rect 33042 22380 33048 22432
rect 33100 22420 33106 22432
rect 33965 22423 34023 22429
rect 33965 22420 33977 22423
rect 33100 22392 33977 22420
rect 33100 22380 33106 22392
rect 33965 22389 33977 22392
rect 34011 22389 34023 22423
rect 33965 22383 34023 22389
rect 1104 22330 35328 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 35328 22330
rect 1104 22256 35328 22278
rect 5350 22176 5356 22228
rect 5408 22216 5414 22228
rect 5626 22216 5632 22228
rect 5408 22188 5632 22216
rect 5408 22176 5414 22188
rect 5626 22176 5632 22188
rect 5684 22176 5690 22228
rect 6178 22176 6184 22228
rect 6236 22216 6242 22228
rect 12066 22216 12072 22228
rect 6236 22188 12072 22216
rect 6236 22176 6242 22188
rect 12066 22176 12072 22188
rect 12124 22176 12130 22228
rect 12894 22216 12900 22228
rect 12176 22188 12900 22216
rect 5166 22148 5172 22160
rect 4356 22120 5172 22148
rect 4356 22089 4384 22120
rect 5166 22108 5172 22120
rect 5224 22108 5230 22160
rect 8938 22108 8944 22160
rect 8996 22148 9002 22160
rect 12176 22148 12204 22188
rect 12894 22176 12900 22188
rect 12952 22176 12958 22228
rect 13262 22176 13268 22228
rect 13320 22216 13326 22228
rect 13633 22219 13691 22225
rect 13633 22216 13645 22219
rect 13320 22188 13645 22216
rect 13320 22176 13326 22188
rect 13633 22185 13645 22188
rect 13679 22185 13691 22219
rect 16850 22216 16856 22228
rect 13633 22179 13691 22185
rect 16132 22188 16856 22216
rect 15470 22148 15476 22160
rect 8996 22120 12204 22148
rect 15396 22120 15476 22148
rect 8996 22108 9002 22120
rect 4341 22083 4399 22089
rect 4341 22049 4353 22083
rect 4387 22049 4399 22083
rect 4341 22043 4399 22049
rect 4522 22040 4528 22092
rect 4580 22080 4586 22092
rect 4580 22052 4844 22080
rect 4580 22040 4586 22052
rect 4617 22015 4675 22021
rect 4617 22012 4629 22015
rect 4172 21984 4629 22012
rect 4172 21888 4200 21984
rect 4617 21981 4629 21984
rect 4663 21981 4675 22015
rect 4617 21975 4675 21981
rect 4706 21972 4712 22024
rect 4764 21972 4770 22024
rect 4816 22021 4844 22052
rect 9858 22040 9864 22092
rect 9916 22080 9922 22092
rect 15396 22089 15424 22120
rect 15470 22108 15476 22120
rect 15528 22148 15534 22160
rect 15657 22151 15715 22157
rect 15657 22148 15669 22151
rect 15528 22120 15669 22148
rect 15528 22108 15534 22120
rect 15657 22117 15669 22120
rect 15703 22148 15715 22151
rect 15746 22148 15752 22160
rect 15703 22120 15752 22148
rect 15703 22117 15715 22120
rect 15657 22111 15715 22117
rect 15746 22108 15752 22120
rect 15804 22108 15810 22160
rect 11057 22083 11115 22089
rect 11057 22080 11069 22083
rect 9916 22052 11069 22080
rect 9916 22040 9922 22052
rect 11057 22049 11069 22052
rect 11103 22080 11115 22083
rect 11333 22083 11391 22089
rect 11333 22080 11345 22083
rect 11103 22052 11345 22080
rect 11103 22049 11115 22052
rect 11057 22043 11115 22049
rect 11333 22049 11345 22052
rect 11379 22080 11391 22083
rect 15381 22083 15439 22089
rect 15381 22080 15393 22083
rect 11379 22052 12296 22080
rect 15359 22052 15393 22080
rect 11379 22049 11391 22052
rect 11333 22043 11391 22049
rect 4801 22015 4859 22021
rect 4801 21981 4813 22015
rect 4847 21981 4859 22015
rect 4801 21975 4859 21981
rect 4893 22015 4951 22021
rect 4893 21981 4905 22015
rect 4939 21981 4951 22015
rect 4893 21975 4951 21981
rect 4985 22015 5043 22021
rect 4985 21981 4997 22015
rect 5031 22012 5043 22015
rect 5261 22015 5319 22021
rect 5261 22012 5273 22015
rect 5031 21984 5273 22012
rect 5031 21981 5043 21984
rect 4985 21975 5043 21981
rect 5261 21981 5273 21984
rect 5307 22012 5319 22015
rect 8478 22012 8484 22024
rect 5307 21984 8484 22012
rect 5307 21981 5319 21984
rect 5261 21975 5319 21981
rect 4724 21944 4752 21972
rect 4540 21916 4752 21944
rect 4908 21944 4936 21975
rect 8478 21972 8484 21984
rect 8536 21972 8542 22024
rect 10781 22015 10839 22021
rect 10781 21981 10793 22015
rect 10827 22012 10839 22015
rect 11238 22012 11244 22024
rect 10827 21984 11244 22012
rect 10827 21981 10839 21984
rect 10781 21975 10839 21981
rect 11238 21972 11244 21984
rect 11296 21972 11302 22024
rect 12158 21972 12164 22024
rect 12216 21972 12222 22024
rect 12268 22012 12296 22052
rect 15381 22049 15393 22052
rect 15427 22049 15439 22083
rect 16132 22080 16160 22188
rect 16850 22176 16856 22188
rect 16908 22176 16914 22228
rect 17402 22176 17408 22228
rect 17460 22216 17466 22228
rect 17460 22188 25452 22216
rect 17460 22176 17466 22188
rect 17218 22108 17224 22160
rect 17276 22148 17282 22160
rect 17497 22151 17555 22157
rect 17497 22148 17509 22151
rect 17276 22120 17509 22148
rect 17276 22108 17282 22120
rect 17497 22117 17509 22120
rect 17543 22117 17555 22151
rect 17497 22111 17555 22117
rect 18966 22108 18972 22160
rect 19024 22148 19030 22160
rect 22189 22151 22247 22157
rect 19024 22120 20852 22148
rect 19024 22108 19030 22120
rect 19521 22083 19579 22089
rect 19521 22080 19533 22083
rect 15381 22043 15439 22049
rect 15488 22052 16160 22080
rect 18340 22052 19533 22080
rect 15488 22012 15516 22052
rect 12268 21984 15516 22012
rect 15930 21972 15936 22024
rect 15988 22012 15994 22024
rect 18340 22021 18368 22052
rect 19521 22049 19533 22052
rect 19567 22080 19579 22083
rect 20438 22080 20444 22092
rect 19567 22052 20444 22080
rect 19567 22049 19579 22052
rect 19521 22043 19579 22049
rect 20438 22040 20444 22052
rect 20496 22040 20502 22092
rect 20824 22089 20852 22120
rect 22189 22117 22201 22151
rect 22235 22117 22247 22151
rect 22189 22111 22247 22117
rect 20809 22083 20867 22089
rect 20809 22080 20821 22083
rect 20787 22052 20821 22080
rect 20809 22049 20821 22052
rect 20855 22049 20867 22083
rect 20809 22043 20867 22049
rect 16117 22015 16175 22021
rect 16117 22012 16129 22015
rect 15988 21984 16129 22012
rect 15988 21972 15994 21984
rect 16117 21981 16129 21984
rect 16163 21981 16175 22015
rect 16117 21975 16175 21981
rect 18325 22015 18383 22021
rect 18325 21981 18337 22015
rect 18371 21981 18383 22015
rect 18325 21975 18383 21981
rect 18601 22015 18659 22021
rect 18601 21981 18613 22015
rect 18647 21981 18659 22015
rect 18601 21975 18659 21981
rect 4908 21916 5028 21944
rect 4540 21888 4568 21916
rect 3142 21836 3148 21888
rect 3200 21876 3206 21888
rect 3789 21879 3847 21885
rect 3789 21876 3801 21879
rect 3200 21848 3801 21876
rect 3200 21836 3206 21848
rect 3789 21845 3801 21848
rect 3835 21845 3847 21879
rect 3789 21839 3847 21845
rect 4154 21836 4160 21888
rect 4212 21836 4218 21888
rect 4249 21879 4307 21885
rect 4249 21845 4261 21879
rect 4295 21876 4307 21879
rect 4522 21876 4528 21888
rect 4295 21848 4528 21876
rect 4295 21845 4307 21848
rect 4249 21839 4307 21845
rect 4522 21836 4528 21848
rect 4580 21836 4586 21888
rect 4706 21836 4712 21888
rect 4764 21876 4770 21888
rect 5000 21876 5028 21916
rect 5534 21904 5540 21956
rect 5592 21904 5598 21956
rect 9674 21904 9680 21956
rect 9732 21944 9738 21956
rect 9861 21947 9919 21953
rect 9861 21944 9873 21947
rect 9732 21916 9873 21944
rect 9732 21904 9738 21916
rect 9861 21913 9873 21916
rect 9907 21913 9919 21947
rect 9861 21907 9919 21913
rect 10873 21947 10931 21953
rect 10873 21913 10885 21947
rect 10919 21944 10931 21947
rect 12428 21947 12486 21953
rect 10919 21916 11652 21944
rect 10919 21913 10931 21916
rect 10873 21907 10931 21913
rect 4764 21848 5028 21876
rect 5169 21879 5227 21885
rect 4764 21836 4770 21848
rect 5169 21845 5181 21879
rect 5215 21876 5227 21879
rect 5552 21876 5580 21904
rect 5215 21848 5580 21876
rect 5215 21845 5227 21848
rect 5169 21839 5227 21845
rect 10410 21836 10416 21888
rect 10468 21836 10474 21888
rect 11624 21876 11652 21916
rect 12428 21913 12440 21947
rect 12474 21944 12486 21947
rect 12802 21944 12808 21956
rect 12474 21916 12808 21944
rect 12474 21913 12486 21916
rect 12428 21907 12486 21913
rect 12802 21904 12808 21916
rect 12860 21904 12866 21956
rect 13170 21904 13176 21956
rect 13228 21944 13234 21956
rect 15289 21947 15347 21953
rect 15289 21944 15301 21947
rect 13228 21916 15301 21944
rect 13228 21904 13234 21916
rect 15289 21913 15301 21916
rect 15335 21944 15347 21947
rect 16384 21947 16442 21953
rect 15335 21916 15976 21944
rect 15335 21913 15347 21916
rect 15289 21907 15347 21913
rect 13188 21876 13216 21904
rect 11624 21848 13216 21876
rect 13541 21879 13599 21885
rect 13541 21845 13553 21879
rect 13587 21876 13599 21879
rect 13814 21876 13820 21888
rect 13587 21848 13820 21876
rect 13587 21845 13599 21848
rect 13541 21839 13599 21845
rect 13814 21836 13820 21848
rect 13872 21836 13878 21888
rect 14826 21836 14832 21888
rect 14884 21836 14890 21888
rect 15194 21836 15200 21888
rect 15252 21836 15258 21888
rect 15838 21836 15844 21888
rect 15896 21836 15902 21888
rect 15948 21876 15976 21916
rect 16384 21913 16396 21947
rect 16430 21944 16442 21947
rect 16666 21944 16672 21956
rect 16430 21916 16672 21944
rect 16430 21913 16442 21916
rect 16384 21907 16442 21913
rect 16666 21904 16672 21916
rect 16724 21904 16730 21956
rect 18233 21947 18291 21953
rect 18233 21913 18245 21947
rect 18279 21944 18291 21947
rect 18616 21944 18644 21975
rect 19242 21972 19248 22024
rect 19300 21972 19306 22024
rect 20070 21972 20076 22024
rect 20128 22012 20134 22024
rect 20165 22015 20223 22021
rect 20165 22012 20177 22015
rect 20128 21984 20177 22012
rect 20128 21972 20134 21984
rect 20165 21981 20177 21984
rect 20211 21981 20223 22015
rect 20625 22015 20683 22021
rect 20625 22012 20637 22015
rect 20165 21975 20223 21981
rect 20364 21984 20637 22012
rect 20254 21944 20260 21956
rect 18279 21916 20260 21944
rect 18279 21913 18291 21916
rect 18233 21907 18291 21913
rect 20254 21904 20260 21916
rect 20312 21904 20318 21956
rect 17034 21876 17040 21888
rect 15948 21848 17040 21876
rect 17034 21836 17040 21848
rect 17092 21836 17098 21888
rect 18509 21879 18567 21885
rect 18509 21845 18521 21879
rect 18555 21876 18567 21879
rect 18690 21876 18696 21888
rect 18555 21848 18696 21876
rect 18555 21845 18567 21848
rect 18509 21839 18567 21845
rect 18690 21836 18696 21848
rect 18748 21836 18754 21888
rect 18782 21836 18788 21888
rect 18840 21876 18846 21888
rect 20364 21885 20392 21984
rect 20625 21981 20637 21984
rect 20671 22012 20683 22015
rect 20714 22012 20720 22024
rect 20671 21984 20720 22012
rect 20671 21981 20683 21984
rect 20625 21975 20683 21981
rect 20714 21972 20720 21984
rect 20772 21972 20778 22024
rect 22204 22012 22232 22111
rect 23658 22108 23664 22160
rect 23716 22148 23722 22160
rect 23753 22151 23811 22157
rect 23753 22148 23765 22151
rect 23716 22120 23765 22148
rect 23716 22108 23722 22120
rect 23753 22117 23765 22120
rect 23799 22117 23811 22151
rect 25424 22148 25452 22188
rect 25498 22176 25504 22228
rect 25556 22176 25562 22228
rect 26421 22219 26479 22225
rect 26421 22185 26433 22219
rect 26467 22216 26479 22219
rect 26510 22216 26516 22228
rect 26467 22188 26516 22216
rect 26467 22185 26479 22188
rect 26421 22179 26479 22185
rect 26510 22176 26516 22188
rect 26568 22176 26574 22228
rect 29086 22216 29092 22228
rect 26620 22188 29092 22216
rect 26620 22148 26648 22188
rect 29086 22176 29092 22188
rect 29144 22176 29150 22228
rect 29181 22219 29239 22225
rect 29181 22185 29193 22219
rect 29227 22216 29239 22219
rect 29227 22188 29316 22216
rect 29227 22185 29239 22188
rect 29181 22179 29239 22185
rect 28445 22151 28503 22157
rect 28445 22148 28457 22151
rect 25424 22120 26648 22148
rect 28368 22120 28457 22148
rect 23753 22111 23811 22117
rect 22830 22040 22836 22092
rect 22888 22040 22894 22092
rect 24026 22040 24032 22092
rect 24084 22080 24090 22092
rect 25774 22080 25780 22092
rect 24084 22052 25780 22080
rect 24084 22040 24090 22052
rect 25774 22040 25780 22052
rect 25832 22040 25838 22092
rect 25958 22040 25964 22092
rect 26016 22040 26022 22092
rect 26142 22040 26148 22092
rect 26200 22080 26206 22092
rect 26513 22083 26571 22089
rect 26513 22080 26525 22083
rect 26200 22052 26525 22080
rect 26200 22040 26206 22052
rect 26513 22049 26525 22052
rect 26559 22049 26571 22083
rect 26513 22043 26571 22049
rect 22462 22012 22468 22024
rect 22204 21984 22468 22012
rect 22462 21972 22468 21984
rect 22520 22012 22526 22024
rect 22649 22015 22707 22021
rect 22649 22012 22661 22015
rect 22520 21984 22661 22012
rect 22520 21972 22526 21984
rect 22649 21981 22661 21984
rect 22695 21981 22707 22015
rect 22649 21975 22707 21981
rect 24213 22015 24271 22021
rect 24213 21981 24225 22015
rect 24259 22012 24271 22015
rect 24302 22012 24308 22024
rect 24259 21984 24308 22012
rect 24259 21981 24271 21984
rect 24213 21975 24271 21981
rect 24302 21972 24308 21984
rect 24360 21972 24366 22024
rect 24489 22015 24547 22021
rect 24489 21981 24501 22015
rect 24535 22012 24547 22015
rect 26602 22012 26608 22024
rect 24535 21984 26608 22012
rect 24535 21981 24547 21984
rect 24489 21975 24547 21981
rect 26602 21972 26608 21984
rect 26660 21972 26666 22024
rect 27062 21972 27068 22024
rect 27120 21972 27126 22024
rect 28368 22012 28396 22120
rect 28445 22117 28457 22120
rect 28491 22117 28503 22151
rect 29288 22148 29316 22188
rect 30558 22176 30564 22228
rect 30616 22176 30622 22228
rect 33042 22225 33048 22228
rect 33032 22219 33048 22225
rect 33032 22185 33044 22219
rect 33032 22179 33048 22185
rect 33042 22176 33048 22179
rect 33100 22176 33106 22228
rect 34514 22176 34520 22228
rect 34572 22176 34578 22228
rect 29362 22148 29368 22160
rect 28445 22111 28503 22117
rect 28966 22120 29224 22148
rect 29288 22120 29368 22148
rect 28966 22080 28994 22120
rect 28828 22052 28994 22080
rect 29196 22080 29224 22120
rect 29362 22108 29368 22120
rect 29420 22108 29426 22160
rect 29454 22080 29460 22092
rect 29196 22052 29460 22080
rect 28534 22012 28540 22024
rect 28368 21984 28540 22012
rect 28534 21972 28540 21984
rect 28592 21972 28598 22024
rect 28626 21972 28632 22024
rect 28684 22012 28690 22024
rect 28828 22021 28856 22052
rect 29454 22040 29460 22052
rect 29512 22080 29518 22092
rect 29512 22052 30972 22080
rect 29512 22040 29518 22052
rect 28721 22015 28779 22021
rect 28721 22012 28733 22015
rect 28684 21984 28733 22012
rect 28684 21972 28690 21984
rect 28721 21981 28733 21984
rect 28767 21981 28779 22015
rect 28721 21975 28779 21981
rect 28813 22015 28871 22021
rect 28813 21981 28825 22015
rect 28859 21981 28871 22015
rect 28813 21975 28871 21981
rect 28951 22015 29009 22021
rect 28951 21981 28963 22015
rect 28997 21988 29009 22015
rect 29270 22012 29276 22024
rect 29196 21988 29276 22012
rect 28997 21984 29276 21988
rect 28997 21981 29224 21984
rect 28951 21975 29224 21981
rect 21076 21947 21134 21953
rect 21076 21913 21088 21947
rect 21122 21944 21134 21947
rect 21122 21916 22324 21944
rect 21122 21913 21134 21916
rect 21076 21907 21134 21913
rect 18969 21879 19027 21885
rect 18969 21876 18981 21879
rect 18840 21848 18981 21876
rect 18840 21836 18846 21848
rect 18969 21845 18981 21848
rect 19015 21845 19027 21879
rect 18969 21839 19027 21845
rect 20349 21879 20407 21885
rect 20349 21845 20361 21879
rect 20395 21876 20407 21879
rect 21174 21876 21180 21888
rect 20395 21848 21180 21876
rect 20395 21845 20407 21848
rect 20349 21839 20407 21845
rect 21174 21836 21180 21848
rect 21232 21836 21238 21888
rect 22296 21885 22324 21916
rect 22738 21904 22744 21956
rect 22796 21944 22802 21956
rect 24854 21944 24860 21956
rect 22796 21916 24164 21944
rect 22796 21904 22802 21916
rect 22281 21879 22339 21885
rect 22281 21845 22293 21879
rect 22327 21845 22339 21879
rect 22281 21839 22339 21845
rect 23014 21836 23020 21888
rect 23072 21876 23078 21888
rect 23109 21879 23167 21885
rect 23109 21876 23121 21879
rect 23072 21848 23121 21876
rect 23072 21836 23078 21848
rect 23109 21845 23121 21848
rect 23155 21876 23167 21879
rect 23382 21876 23388 21888
rect 23155 21848 23388 21876
rect 23155 21845 23167 21848
rect 23109 21839 23167 21845
rect 23382 21836 23388 21848
rect 23440 21836 23446 21888
rect 23658 21836 23664 21888
rect 23716 21876 23722 21888
rect 24026 21876 24032 21888
rect 23716 21848 24032 21876
rect 23716 21836 23722 21848
rect 24026 21836 24032 21848
rect 24084 21836 24090 21888
rect 24136 21876 24164 21916
rect 24412 21916 24860 21944
rect 24412 21876 24440 21916
rect 24854 21904 24860 21916
rect 24912 21904 24918 21956
rect 24946 21904 24952 21956
rect 25004 21944 25010 21956
rect 25222 21944 25228 21956
rect 25004 21916 25228 21944
rect 25004 21904 25010 21916
rect 25222 21904 25228 21916
rect 25280 21904 25286 21956
rect 25314 21904 25320 21956
rect 25372 21944 25378 21956
rect 25869 21947 25927 21953
rect 25869 21944 25881 21947
rect 25372 21916 25881 21944
rect 25372 21904 25378 21916
rect 25869 21913 25881 21916
rect 25915 21913 25927 21947
rect 25869 21907 25927 21913
rect 24136 21848 24440 21876
rect 26620 21876 26648 21972
rect 28966 21960 29224 21975
rect 29270 21972 29276 21984
rect 29328 21972 29334 22024
rect 29362 21972 29368 22024
rect 29420 21972 29426 22024
rect 29546 21972 29552 22024
rect 29604 22012 29610 22024
rect 30374 22012 30380 22024
rect 29604 21984 30380 22012
rect 29604 21972 29610 21984
rect 30374 21972 30380 21984
rect 30432 21972 30438 22024
rect 30944 22021 30972 22052
rect 31018 22040 31024 22092
rect 31076 22080 31082 22092
rect 31113 22083 31171 22089
rect 31113 22080 31125 22083
rect 31076 22052 31125 22080
rect 31076 22040 31082 22052
rect 31113 22049 31125 22052
rect 31159 22049 31171 22083
rect 32769 22083 32827 22089
rect 32769 22080 32781 22083
rect 31113 22043 31171 22049
rect 31726 22052 32781 22080
rect 30929 22015 30987 22021
rect 30929 21981 30941 22015
rect 30975 21981 30987 22015
rect 31386 22012 31392 22024
rect 30929 21975 30987 21981
rect 31312 21984 31392 22012
rect 27332 21947 27390 21953
rect 27332 21913 27344 21947
rect 27378 21944 27390 21947
rect 27614 21944 27620 21956
rect 27378 21916 27620 21944
rect 27378 21913 27390 21916
rect 27332 21907 27390 21913
rect 27614 21904 27620 21916
rect 27672 21904 27678 21956
rect 29638 21904 29644 21956
rect 29696 21944 29702 21956
rect 30285 21947 30343 21953
rect 30285 21944 30297 21947
rect 29696 21916 30297 21944
rect 29696 21904 29702 21916
rect 30285 21913 30297 21916
rect 30331 21944 30343 21947
rect 31312 21944 31340 21984
rect 31386 21972 31392 21984
rect 31444 22012 31450 22024
rect 31726 22012 31754 22052
rect 32769 22049 32781 22052
rect 32815 22080 32827 22083
rect 33134 22080 33140 22092
rect 32815 22052 33140 22080
rect 32815 22049 32827 22052
rect 32769 22043 32827 22049
rect 33134 22040 33140 22052
rect 33192 22040 33198 22092
rect 31444 21984 31754 22012
rect 31444 21972 31450 21984
rect 30331 21916 31340 21944
rect 30331 21913 30343 21916
rect 30285 21907 30343 21913
rect 33502 21904 33508 21956
rect 33560 21904 33566 21956
rect 28810 21876 28816 21888
rect 26620 21848 28816 21876
rect 28810 21836 28816 21848
rect 28868 21836 28874 21888
rect 28902 21836 28908 21888
rect 28960 21876 28966 21888
rect 28994 21876 29000 21888
rect 28960 21848 29000 21876
rect 28960 21836 28966 21848
rect 28994 21836 29000 21848
rect 29052 21836 29058 21888
rect 29089 21879 29147 21885
rect 29089 21845 29101 21879
rect 29135 21876 29147 21879
rect 29454 21876 29460 21888
rect 29135 21848 29460 21876
rect 29135 21845 29147 21848
rect 29089 21839 29147 21845
rect 29454 21836 29460 21848
rect 29512 21836 29518 21888
rect 31018 21836 31024 21888
rect 31076 21876 31082 21888
rect 31389 21879 31447 21885
rect 31389 21876 31401 21879
rect 31076 21848 31401 21876
rect 31076 21836 31082 21848
rect 31389 21845 31401 21848
rect 31435 21845 31447 21879
rect 31389 21839 31447 21845
rect 1104 21786 35328 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35328 21786
rect 1104 21712 35328 21734
rect 1857 21675 1915 21681
rect 1857 21641 1869 21675
rect 1903 21672 1915 21675
rect 4154 21672 4160 21684
rect 1903 21644 4160 21672
rect 1903 21641 1915 21644
rect 1857 21635 1915 21641
rect 4154 21632 4160 21644
rect 4212 21632 4218 21684
rect 4706 21632 4712 21684
rect 4764 21632 4770 21684
rect 7929 21675 7987 21681
rect 7929 21672 7941 21675
rect 7760 21644 7941 21672
rect 2992 21607 3050 21613
rect 2992 21573 3004 21607
rect 3038 21604 3050 21607
rect 3142 21604 3148 21616
rect 3038 21576 3148 21604
rect 3038 21573 3050 21576
rect 2992 21567 3050 21573
rect 3142 21564 3148 21576
rect 3200 21564 3206 21616
rect 4614 21604 4620 21616
rect 3344 21576 4620 21604
rect 3344 21545 3372 21576
rect 4614 21564 4620 21576
rect 4672 21564 4678 21616
rect 5350 21564 5356 21616
rect 5408 21604 5414 21616
rect 6454 21604 6460 21616
rect 5408 21576 6460 21604
rect 5408 21564 5414 21576
rect 6454 21564 6460 21576
rect 6512 21564 6518 21616
rect 7592 21607 7650 21613
rect 7592 21573 7604 21607
rect 7638 21604 7650 21607
rect 7760 21604 7788 21644
rect 7929 21641 7941 21644
rect 7975 21641 7987 21675
rect 7929 21635 7987 21641
rect 8294 21632 8300 21684
rect 8352 21672 8358 21684
rect 8389 21675 8447 21681
rect 8389 21672 8401 21675
rect 8352 21644 8401 21672
rect 8352 21632 8358 21644
rect 8389 21641 8401 21644
rect 8435 21641 8447 21675
rect 8389 21635 8447 21641
rect 9858 21632 9864 21684
rect 9916 21632 9922 21684
rect 10873 21675 10931 21681
rect 10873 21641 10885 21675
rect 10919 21672 10931 21675
rect 10962 21672 10968 21684
rect 10919 21644 10968 21672
rect 10919 21641 10931 21644
rect 10873 21635 10931 21641
rect 8110 21604 8116 21616
rect 7638 21576 7788 21604
rect 7852 21576 8116 21604
rect 7638 21573 7650 21576
rect 7592 21567 7650 21573
rect 3237 21539 3295 21545
rect 3237 21505 3249 21539
rect 3283 21536 3295 21539
rect 3329 21539 3387 21545
rect 3329 21536 3341 21539
rect 3283 21508 3341 21536
rect 3283 21505 3295 21508
rect 3237 21499 3295 21505
rect 3329 21505 3341 21508
rect 3375 21505 3387 21539
rect 3329 21499 3387 21505
rect 3596 21539 3654 21545
rect 3596 21505 3608 21539
rect 3642 21536 3654 21539
rect 4062 21536 4068 21548
rect 3642 21508 4068 21536
rect 3642 21505 3654 21508
rect 3596 21499 3654 21505
rect 4062 21496 4068 21508
rect 4120 21496 4126 21548
rect 5068 21539 5126 21545
rect 5068 21505 5080 21539
rect 5114 21536 5126 21539
rect 5810 21536 5816 21548
rect 5114 21508 5816 21536
rect 5114 21505 5126 21508
rect 5068 21499 5126 21505
rect 5810 21496 5816 21508
rect 5868 21496 5874 21548
rect 7852 21545 7880 21576
rect 8110 21564 8116 21576
rect 8168 21604 8174 21616
rect 9766 21604 9772 21616
rect 8168 21576 9772 21604
rect 8168 21564 8174 21576
rect 9766 21564 9772 21576
rect 9824 21564 9830 21616
rect 7837 21539 7895 21545
rect 7837 21505 7849 21539
rect 7883 21505 7895 21539
rect 8297 21539 8355 21545
rect 8297 21536 8309 21539
rect 7837 21499 7895 21505
rect 7944 21508 8309 21536
rect 4798 21428 4804 21480
rect 4856 21428 4862 21480
rect 4430 21292 4436 21344
rect 4488 21332 4494 21344
rect 4706 21332 4712 21344
rect 4488 21304 4712 21332
rect 4488 21292 4494 21304
rect 4706 21292 4712 21304
rect 4764 21292 4770 21344
rect 6178 21292 6184 21344
rect 6236 21292 6242 21344
rect 6457 21335 6515 21341
rect 6457 21301 6469 21335
rect 6503 21332 6515 21335
rect 7466 21332 7472 21344
rect 6503 21304 7472 21332
rect 6503 21301 6515 21304
rect 6457 21295 6515 21301
rect 7466 21292 7472 21304
rect 7524 21332 7530 21344
rect 7944 21332 7972 21508
rect 8297 21505 8309 21508
rect 8343 21505 8355 21539
rect 10229 21539 10287 21545
rect 8297 21499 8355 21505
rect 8404 21508 8984 21536
rect 8018 21428 8024 21480
rect 8076 21468 8082 21480
rect 8404 21468 8432 21508
rect 8076 21440 8432 21468
rect 8573 21471 8631 21477
rect 8076 21428 8082 21440
rect 8573 21437 8585 21471
rect 8619 21468 8631 21471
rect 8846 21468 8852 21480
rect 8619 21440 8852 21468
rect 8619 21437 8631 21440
rect 8573 21431 8631 21437
rect 8846 21428 8852 21440
rect 8904 21428 8910 21480
rect 8956 21468 8984 21508
rect 10229 21505 10241 21539
rect 10275 21536 10287 21539
rect 10888 21536 10916 21635
rect 10962 21632 10968 21644
rect 11020 21632 11026 21684
rect 12802 21632 12808 21684
rect 12860 21632 12866 21684
rect 13170 21632 13176 21684
rect 13228 21632 13234 21684
rect 15194 21632 15200 21684
rect 15252 21672 15258 21684
rect 15657 21675 15715 21681
rect 15657 21672 15669 21675
rect 15252 21644 15669 21672
rect 15252 21632 15258 21644
rect 15657 21641 15669 21644
rect 15703 21672 15715 21675
rect 16114 21672 16120 21684
rect 15703 21644 16120 21672
rect 15703 21641 15715 21644
rect 15657 21635 15715 21641
rect 16114 21632 16120 21644
rect 16172 21632 16178 21684
rect 16666 21632 16672 21684
rect 16724 21632 16730 21684
rect 17034 21632 17040 21684
rect 17092 21632 17098 21684
rect 17129 21675 17187 21681
rect 17129 21641 17141 21675
rect 17175 21672 17187 21675
rect 17218 21672 17224 21684
rect 17175 21644 17224 21672
rect 17175 21641 17187 21644
rect 17129 21635 17187 21641
rect 17218 21632 17224 21644
rect 17276 21632 17282 21684
rect 18598 21632 18604 21684
rect 18656 21672 18662 21684
rect 18969 21675 19027 21681
rect 18969 21672 18981 21675
rect 18656 21644 18981 21672
rect 18656 21632 18662 21644
rect 18969 21641 18981 21644
rect 19015 21672 19027 21675
rect 19015 21644 20576 21672
rect 19015 21641 19027 21644
rect 18969 21635 19027 21641
rect 13265 21607 13323 21613
rect 13265 21573 13277 21607
rect 13311 21604 13323 21607
rect 13814 21604 13820 21616
rect 13311 21576 13820 21604
rect 13311 21573 13323 21576
rect 13265 21567 13323 21573
rect 13814 21564 13820 21576
rect 13872 21564 13878 21616
rect 14544 21607 14602 21613
rect 14544 21573 14556 21607
rect 14590 21604 14602 21607
rect 14826 21604 14832 21616
rect 14590 21576 14832 21604
rect 14590 21573 14602 21576
rect 14544 21567 14602 21573
rect 14826 21564 14832 21576
rect 14884 21564 14890 21616
rect 15746 21564 15752 21616
rect 15804 21564 15810 21616
rect 17494 21604 17500 21616
rect 16040 21576 17500 21604
rect 16040 21536 16068 21576
rect 17494 21564 17500 21576
rect 17552 21564 17558 21616
rect 17604 21576 19012 21604
rect 17604 21545 17632 21576
rect 18984 21548 19012 21576
rect 10275 21508 10916 21536
rect 12406 21508 16068 21536
rect 16117 21539 16175 21545
rect 10275 21505 10287 21508
rect 10229 21499 10287 21505
rect 12406 21468 12434 21508
rect 16117 21505 16129 21539
rect 16163 21536 16175 21539
rect 17589 21539 17647 21545
rect 16163 21508 16528 21536
rect 16163 21505 16175 21508
rect 16117 21499 16175 21505
rect 8956 21440 12434 21468
rect 13354 21428 13360 21480
rect 13412 21468 13418 21480
rect 13633 21471 13691 21477
rect 13633 21468 13645 21471
rect 13412 21440 13645 21468
rect 13412 21428 13418 21440
rect 13633 21437 13645 21440
rect 13679 21437 13691 21471
rect 13633 21431 13691 21437
rect 14277 21471 14335 21477
rect 14277 21437 14289 21471
rect 14323 21437 14335 21471
rect 14277 21431 14335 21437
rect 8864 21341 8892 21428
rect 7524 21304 7972 21332
rect 8849 21335 8907 21341
rect 7524 21292 7530 21304
rect 8849 21301 8861 21335
rect 8895 21332 8907 21335
rect 9582 21332 9588 21344
rect 8895 21304 9588 21332
rect 8895 21301 8907 21304
rect 8849 21295 8907 21301
rect 9582 21292 9588 21304
rect 9640 21292 9646 21344
rect 10410 21292 10416 21344
rect 10468 21332 10474 21344
rect 10597 21335 10655 21341
rect 10597 21332 10609 21335
rect 10468 21304 10609 21332
rect 10468 21292 10474 21304
rect 10597 21301 10609 21304
rect 10643 21301 10655 21335
rect 14292 21332 14320 21431
rect 14550 21332 14556 21344
rect 14292 21304 14556 21332
rect 10597 21295 10655 21301
rect 14550 21292 14556 21304
rect 14608 21292 14614 21344
rect 16500 21341 16528 21508
rect 17589 21505 17601 21539
rect 17635 21505 17647 21539
rect 17589 21499 17647 21505
rect 17856 21539 17914 21545
rect 17856 21505 17868 21539
rect 17902 21536 17914 21539
rect 18138 21536 18144 21548
rect 17902 21508 18144 21536
rect 17902 21505 17914 21508
rect 17856 21499 17914 21505
rect 18138 21496 18144 21508
rect 18196 21496 18202 21548
rect 18966 21496 18972 21548
rect 19024 21536 19030 21548
rect 19061 21539 19119 21545
rect 19061 21536 19073 21539
rect 19024 21508 19073 21536
rect 19024 21496 19030 21508
rect 19061 21505 19073 21508
rect 19107 21505 19119 21539
rect 19061 21499 19119 21505
rect 19328 21539 19386 21545
rect 19328 21505 19340 21539
rect 19374 21536 19386 21539
rect 19610 21536 19616 21548
rect 19374 21508 19616 21536
rect 19374 21505 19386 21508
rect 19328 21499 19386 21505
rect 19610 21496 19616 21508
rect 19668 21496 19674 21548
rect 20548 21545 20576 21644
rect 21174 21632 21180 21684
rect 21232 21632 21238 21684
rect 22094 21632 22100 21684
rect 22152 21672 22158 21684
rect 22922 21672 22928 21684
rect 22152 21644 22928 21672
rect 22152 21632 22158 21644
rect 22922 21632 22928 21644
rect 22980 21632 22986 21684
rect 23017 21675 23075 21681
rect 23017 21641 23029 21675
rect 23063 21672 23075 21675
rect 24210 21672 24216 21684
rect 23063 21644 24216 21672
rect 23063 21641 23075 21644
rect 23017 21635 23075 21641
rect 24210 21632 24216 21644
rect 24268 21632 24274 21684
rect 24765 21675 24823 21681
rect 24765 21672 24777 21675
rect 24320 21644 24777 21672
rect 20717 21607 20775 21613
rect 20717 21573 20729 21607
rect 20763 21573 20775 21607
rect 20717 21567 20775 21573
rect 20533 21539 20591 21545
rect 20533 21505 20545 21539
rect 20579 21505 20591 21539
rect 20533 21499 20591 21505
rect 20732 21480 20760 21567
rect 22002 21564 22008 21616
rect 22060 21604 22066 21616
rect 22649 21607 22707 21613
rect 22649 21604 22661 21607
rect 22060 21576 22661 21604
rect 22060 21564 22066 21576
rect 22649 21573 22661 21576
rect 22695 21573 22707 21607
rect 22940 21604 22968 21632
rect 23109 21607 23167 21613
rect 23109 21604 23121 21607
rect 22940 21576 23121 21604
rect 22649 21567 22707 21573
rect 23109 21573 23121 21576
rect 23155 21573 23167 21607
rect 23109 21567 23167 21573
rect 23560 21607 23618 21613
rect 23560 21573 23572 21607
rect 23606 21604 23618 21607
rect 24320 21604 24348 21644
rect 24765 21641 24777 21644
rect 24811 21641 24823 21675
rect 24765 21635 24823 21641
rect 24854 21632 24860 21684
rect 24912 21672 24918 21684
rect 25225 21675 25283 21681
rect 25225 21672 25237 21675
rect 24912 21644 25237 21672
rect 24912 21632 24918 21644
rect 25225 21641 25237 21644
rect 25271 21641 25283 21675
rect 25225 21635 25283 21641
rect 26050 21632 26056 21684
rect 26108 21632 26114 21684
rect 27522 21632 27528 21684
rect 27580 21632 27586 21684
rect 27614 21632 27620 21684
rect 27672 21632 27678 21684
rect 27985 21675 28043 21681
rect 27985 21641 27997 21675
rect 28031 21672 28043 21675
rect 28534 21672 28540 21684
rect 28031 21644 28540 21672
rect 28031 21641 28043 21644
rect 27985 21635 28043 21641
rect 28534 21632 28540 21644
rect 28592 21632 28598 21684
rect 28810 21632 28816 21684
rect 28868 21672 28874 21684
rect 29457 21675 29515 21681
rect 29457 21672 29469 21675
rect 28868 21644 28994 21672
rect 28868 21632 28874 21644
rect 26145 21607 26203 21613
rect 26145 21604 26157 21607
rect 23606 21576 24348 21604
rect 25056 21576 26157 21604
rect 23606 21573 23618 21576
rect 23560 21567 23618 21573
rect 20809 21539 20867 21545
rect 20809 21505 20821 21539
rect 20855 21505 20867 21539
rect 20809 21499 20867 21505
rect 17310 21428 17316 21480
rect 17368 21428 17374 21480
rect 20714 21428 20720 21480
rect 20772 21428 20778 21480
rect 20824 21400 20852 21499
rect 20898 21496 20904 21548
rect 20956 21496 20962 21548
rect 22278 21496 22284 21548
rect 22336 21496 22342 21548
rect 22373 21539 22431 21545
rect 22373 21505 22385 21539
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 20456 21372 20852 21400
rect 21085 21403 21143 21409
rect 20456 21344 20484 21372
rect 21085 21369 21097 21403
rect 21131 21400 21143 21403
rect 22388 21400 22416 21499
rect 22462 21496 22468 21548
rect 22520 21536 22526 21548
rect 22520 21508 22565 21536
rect 22520 21496 22526 21508
rect 22738 21496 22744 21548
rect 22796 21496 22802 21548
rect 22879 21539 22937 21545
rect 22879 21505 22891 21539
rect 22925 21536 22937 21539
rect 23014 21536 23020 21548
rect 22925 21508 23020 21536
rect 22925 21505 22937 21508
rect 22879 21499 22937 21505
rect 23014 21496 23020 21508
rect 23072 21496 23078 21548
rect 24026 21496 24032 21548
rect 24084 21536 24090 21548
rect 25056 21536 25084 21576
rect 25608 21545 25636 21576
rect 26145 21573 26157 21576
rect 26191 21573 26203 21607
rect 26145 21567 26203 21573
rect 27430 21564 27436 21616
rect 27488 21604 27494 21616
rect 28721 21607 28779 21613
rect 28721 21604 28733 21607
rect 27488 21576 28733 21604
rect 27488 21564 27494 21576
rect 28721 21573 28733 21576
rect 28767 21573 28779 21607
rect 28966 21604 28994 21644
rect 29196 21644 29469 21672
rect 29196 21604 29224 21644
rect 29457 21641 29469 21644
rect 29503 21672 29515 21675
rect 29546 21672 29552 21684
rect 29503 21644 29552 21672
rect 29503 21641 29515 21644
rect 29457 21635 29515 21641
rect 29546 21632 29552 21644
rect 29604 21632 29610 21684
rect 29730 21632 29736 21684
rect 29788 21632 29794 21684
rect 29914 21632 29920 21684
rect 29972 21632 29978 21684
rect 28966 21576 29224 21604
rect 29273 21607 29331 21613
rect 28721 21567 28779 21573
rect 29273 21573 29285 21607
rect 29319 21604 29331 21607
rect 29362 21604 29368 21616
rect 29319 21576 29368 21604
rect 29319 21573 29331 21576
rect 29273 21567 29331 21573
rect 29362 21564 29368 21576
rect 29420 21564 29426 21616
rect 24084 21508 25084 21536
rect 25133 21539 25191 21545
rect 24084 21496 24090 21508
rect 25133 21505 25145 21539
rect 25179 21505 25191 21539
rect 25133 21499 25191 21505
rect 25593 21539 25651 21545
rect 25593 21505 25605 21539
rect 25639 21505 25651 21539
rect 28624 21539 28682 21545
rect 28624 21536 28636 21539
rect 25593 21499 25651 21505
rect 28552 21508 28636 21536
rect 23293 21471 23351 21477
rect 23293 21437 23305 21471
rect 23339 21437 23351 21471
rect 23293 21431 23351 21437
rect 21131 21372 22416 21400
rect 21131 21369 21143 21372
rect 21085 21363 21143 21369
rect 16485 21335 16543 21341
rect 16485 21301 16497 21335
rect 16531 21332 16543 21335
rect 18506 21332 18512 21344
rect 16531 21304 18512 21332
rect 16531 21301 16543 21304
rect 16485 21295 16543 21301
rect 18506 21292 18512 21304
rect 18564 21292 18570 21344
rect 20438 21292 20444 21344
rect 20496 21292 20502 21344
rect 20898 21292 20904 21344
rect 20956 21332 20962 21344
rect 21821 21335 21879 21341
rect 21821 21332 21833 21335
rect 20956 21304 21833 21332
rect 20956 21292 20962 21304
rect 21821 21301 21833 21304
rect 21867 21332 21879 21335
rect 22002 21332 22008 21344
rect 21867 21304 22008 21332
rect 21867 21301 21879 21304
rect 21821 21295 21879 21301
rect 22002 21292 22008 21304
rect 22060 21332 22066 21344
rect 22094 21332 22100 21344
rect 22060 21304 22100 21332
rect 22060 21292 22066 21304
rect 22094 21292 22100 21304
rect 22152 21292 22158 21344
rect 23308 21332 23336 21431
rect 24302 21360 24308 21412
rect 24360 21400 24366 21412
rect 24673 21403 24731 21409
rect 24673 21400 24685 21403
rect 24360 21372 24685 21400
rect 24360 21360 24366 21372
rect 24673 21369 24685 21372
rect 24719 21400 24731 21403
rect 25148 21400 25176 21499
rect 25409 21471 25467 21477
rect 25409 21437 25421 21471
rect 25455 21468 25467 21471
rect 25498 21468 25504 21480
rect 25455 21440 25504 21468
rect 25455 21437 25467 21440
rect 25409 21431 25467 21437
rect 25498 21428 25504 21440
rect 25556 21468 25562 21480
rect 26050 21468 26056 21480
rect 25556 21440 26056 21468
rect 25556 21428 25562 21440
rect 26050 21428 26056 21440
rect 26108 21428 26114 21480
rect 27890 21428 27896 21480
rect 27948 21468 27954 21480
rect 28077 21471 28135 21477
rect 28077 21468 28089 21471
rect 27948 21440 28089 21468
rect 27948 21428 27954 21440
rect 28077 21437 28089 21440
rect 28123 21437 28135 21471
rect 28077 21431 28135 21437
rect 28166 21428 28172 21480
rect 28224 21428 28230 21480
rect 28552 21468 28580 21508
rect 28624 21505 28636 21508
rect 28670 21505 28682 21539
rect 28624 21499 28682 21505
rect 28810 21496 28816 21548
rect 28868 21496 28874 21548
rect 28902 21496 28908 21548
rect 28960 21545 28966 21548
rect 28960 21539 28999 21545
rect 28987 21505 28999 21539
rect 28960 21499 28999 21505
rect 29089 21539 29147 21545
rect 29089 21505 29101 21539
rect 29135 21536 29147 21539
rect 29454 21536 29460 21548
rect 29135 21508 29460 21536
rect 29135 21505 29147 21508
rect 29089 21499 29147 21505
rect 28960 21496 28966 21499
rect 29454 21496 29460 21508
rect 29512 21496 29518 21548
rect 30285 21539 30343 21545
rect 30285 21505 30297 21539
rect 30331 21505 30343 21539
rect 30285 21499 30343 21505
rect 28267 21440 28580 21468
rect 24719 21372 25176 21400
rect 24719 21369 24731 21372
rect 24673 21363 24731 21369
rect 26878 21360 26884 21412
rect 26936 21400 26942 21412
rect 27522 21400 27528 21412
rect 26936 21372 27528 21400
rect 26936 21360 26942 21372
rect 27522 21360 27528 21372
rect 27580 21400 27586 21412
rect 28267 21400 28295 21440
rect 28718 21428 28724 21480
rect 28776 21468 28782 21480
rect 30300 21468 30328 21499
rect 28776 21440 30328 21468
rect 30377 21471 30435 21477
rect 28776 21428 28782 21440
rect 30377 21437 30389 21471
rect 30423 21437 30435 21471
rect 30377 21431 30435 21437
rect 30469 21471 30527 21477
rect 30469 21437 30481 21471
rect 30515 21437 30527 21471
rect 30469 21431 30527 21437
rect 27580 21372 28295 21400
rect 28445 21403 28503 21409
rect 27580 21360 27586 21372
rect 28445 21369 28457 21403
rect 28491 21400 28503 21403
rect 29822 21400 29828 21412
rect 28491 21372 29828 21400
rect 28491 21369 28503 21372
rect 28445 21363 28503 21369
rect 29822 21360 29828 21372
rect 29880 21360 29886 21412
rect 30282 21360 30288 21412
rect 30340 21400 30346 21412
rect 30392 21400 30420 21431
rect 30340 21372 30420 21400
rect 30484 21400 30512 21431
rect 30926 21400 30932 21412
rect 30484 21372 30932 21400
rect 30340 21360 30346 21372
rect 23474 21332 23480 21344
rect 23308 21304 23480 21332
rect 23474 21292 23480 21304
rect 23532 21292 23538 21344
rect 25774 21292 25780 21344
rect 25832 21332 25838 21344
rect 26329 21335 26387 21341
rect 26329 21332 26341 21335
rect 25832 21304 26341 21332
rect 25832 21292 25838 21304
rect 26329 21301 26341 21304
rect 26375 21301 26387 21335
rect 26329 21295 26387 21301
rect 28350 21292 28356 21344
rect 28408 21332 28414 21344
rect 30484 21332 30512 21372
rect 30926 21360 30932 21372
rect 30984 21400 30990 21412
rect 31202 21400 31208 21412
rect 30984 21372 31208 21400
rect 30984 21360 30990 21372
rect 31202 21360 31208 21372
rect 31260 21360 31266 21412
rect 28408 21304 30512 21332
rect 28408 21292 28414 21304
rect 30742 21292 30748 21344
rect 30800 21292 30806 21344
rect 1104 21242 35328 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 35328 21242
rect 1104 21168 35328 21190
rect 4062 21088 4068 21140
rect 4120 21128 4126 21140
rect 4157 21131 4215 21137
rect 4157 21128 4169 21131
rect 4120 21100 4169 21128
rect 4120 21088 4126 21100
rect 4157 21097 4169 21100
rect 4203 21097 4215 21131
rect 4157 21091 4215 21097
rect 5810 21088 5816 21140
rect 5868 21088 5874 21140
rect 7190 21128 7196 21140
rect 6196 21100 7196 21128
rect 6196 21060 6224 21100
rect 7190 21088 7196 21100
rect 7248 21088 7254 21140
rect 7745 21131 7803 21137
rect 7745 21097 7757 21131
rect 7791 21128 7803 21131
rect 7834 21128 7840 21140
rect 7791 21100 7840 21128
rect 7791 21097 7803 21100
rect 7745 21091 7803 21097
rect 7834 21088 7840 21100
rect 7892 21088 7898 21140
rect 7929 21131 7987 21137
rect 7929 21097 7941 21131
rect 7975 21128 7987 21131
rect 8018 21128 8024 21140
rect 7975 21100 8024 21128
rect 7975 21097 7987 21100
rect 7929 21091 7987 21097
rect 8018 21088 8024 21100
rect 8076 21088 8082 21140
rect 8113 21131 8171 21137
rect 8113 21097 8125 21131
rect 8159 21128 8171 21131
rect 8386 21128 8392 21140
rect 8159 21100 8392 21128
rect 8159 21097 8171 21100
rect 8113 21091 8171 21097
rect 8386 21088 8392 21100
rect 8444 21088 8450 21140
rect 8496 21100 14044 21128
rect 5000 21032 6224 21060
rect 5000 21001 5028 21032
rect 6454 21020 6460 21072
rect 6512 21060 6518 21072
rect 8496 21060 8524 21100
rect 6512 21032 8524 21060
rect 14016 21060 14044 21100
rect 14090 21088 14096 21140
rect 14148 21128 14154 21140
rect 14277 21131 14335 21137
rect 14277 21128 14289 21131
rect 14148 21100 14289 21128
rect 14148 21088 14154 21100
rect 14277 21097 14289 21100
rect 14323 21097 14335 21131
rect 14277 21091 14335 21097
rect 15746 21088 15752 21140
rect 15804 21128 15810 21140
rect 16485 21131 16543 21137
rect 16485 21128 16497 21131
rect 15804 21100 16497 21128
rect 15804 21088 15810 21100
rect 16485 21097 16497 21100
rect 16531 21097 16543 21131
rect 16485 21091 16543 21097
rect 18138 21088 18144 21140
rect 18196 21088 18202 21140
rect 19610 21088 19616 21140
rect 19668 21088 19674 21140
rect 20441 21131 20499 21137
rect 20441 21128 20453 21131
rect 19720 21100 20453 21128
rect 18782 21060 18788 21072
rect 14016 21032 18788 21060
rect 6512 21020 6518 21032
rect 4801 20995 4859 21001
rect 4801 20961 4813 20995
rect 4847 20992 4859 20995
rect 4985 20995 5043 21001
rect 4985 20992 4997 20995
rect 4847 20964 4997 20992
rect 4847 20961 4859 20964
rect 4801 20955 4859 20961
rect 4985 20961 4997 20964
rect 5031 20961 5043 20995
rect 4985 20955 5043 20961
rect 6362 20952 6368 21004
rect 6420 20952 6426 21004
rect 9585 20995 9643 21001
rect 9585 20961 9597 20995
rect 9631 20961 9643 20995
rect 9585 20955 9643 20961
rect 4525 20927 4583 20933
rect 4525 20893 4537 20927
rect 4571 20924 4583 20927
rect 4890 20924 4896 20936
rect 4571 20896 4896 20924
rect 4571 20893 4583 20896
rect 4525 20887 4583 20893
rect 4890 20884 4896 20896
rect 4948 20884 4954 20936
rect 6178 20884 6184 20936
rect 6236 20924 6242 20936
rect 7193 20927 7251 20933
rect 7193 20924 7205 20927
rect 6236 20896 7205 20924
rect 6236 20884 6242 20896
rect 7193 20893 7205 20896
rect 7239 20893 7251 20927
rect 7193 20887 7251 20893
rect 7466 20884 7472 20936
rect 7524 20884 7530 20936
rect 7561 20927 7619 20933
rect 7561 20893 7573 20927
rect 7607 20924 7619 20927
rect 8386 20924 8392 20936
rect 7607 20896 8392 20924
rect 7607 20893 7619 20896
rect 7561 20887 7619 20893
rect 8386 20884 8392 20896
rect 8444 20884 8450 20936
rect 9600 20924 9628 20955
rect 9766 20952 9772 21004
rect 9824 20952 9830 21004
rect 18598 20952 18604 21004
rect 18656 20952 18662 21004
rect 18708 21001 18736 21032
rect 18782 21020 18788 21032
rect 18840 21060 18846 21072
rect 18969 21063 19027 21069
rect 18969 21060 18981 21063
rect 18840 21032 18981 21060
rect 18840 21020 18846 21032
rect 18969 21029 18981 21032
rect 19015 21029 19027 21063
rect 19720 21060 19748 21100
rect 20441 21097 20453 21100
rect 20487 21128 20499 21131
rect 20806 21128 20812 21140
rect 20487 21100 20812 21128
rect 20487 21097 20499 21100
rect 20441 21091 20499 21097
rect 20806 21088 20812 21100
rect 20864 21088 20870 21140
rect 25866 21088 25872 21140
rect 25924 21128 25930 21140
rect 25924 21100 27384 21128
rect 25924 21088 25930 21100
rect 18969 21023 19027 21029
rect 19076 21032 19748 21060
rect 18693 20995 18751 21001
rect 18693 20961 18705 20995
rect 18739 20961 18751 20995
rect 19076 20992 19104 21032
rect 20070 21020 20076 21072
rect 20128 21060 20134 21072
rect 22002 21060 22008 21072
rect 20128 21032 22008 21060
rect 20128 21020 20134 21032
rect 22002 21020 22008 21032
rect 22060 21020 22066 21072
rect 23842 21020 23848 21072
rect 23900 21060 23906 21072
rect 24118 21060 24124 21072
rect 23900 21032 24124 21060
rect 23900 21020 23906 21032
rect 24118 21020 24124 21032
rect 24176 21060 24182 21072
rect 24397 21063 24455 21069
rect 24397 21060 24409 21063
rect 24176 21032 24409 21060
rect 24176 21020 24182 21032
rect 24397 21029 24409 21032
rect 24443 21029 24455 21063
rect 27356 21060 27384 21100
rect 27430 21088 27436 21140
rect 27488 21088 27494 21140
rect 29273 21131 29331 21137
rect 27540 21100 28994 21128
rect 27540 21060 27568 21100
rect 27356 21032 27568 21060
rect 28966 21060 28994 21100
rect 29273 21097 29285 21131
rect 29319 21128 29331 21131
rect 29362 21128 29368 21140
rect 29319 21100 29368 21128
rect 29319 21097 29331 21100
rect 29273 21091 29331 21097
rect 29362 21088 29368 21100
rect 29420 21128 29426 21140
rect 30006 21128 30012 21140
rect 29420 21100 30012 21128
rect 29420 21088 29426 21100
rect 30006 21088 30012 21100
rect 30064 21088 30070 21140
rect 30282 21088 30288 21140
rect 30340 21128 30346 21140
rect 31021 21131 31079 21137
rect 31021 21128 31033 21131
rect 30340 21100 31033 21128
rect 30340 21088 30346 21100
rect 31021 21097 31033 21100
rect 31067 21097 31079 21131
rect 31021 21091 31079 21097
rect 31202 21088 31208 21140
rect 31260 21128 31266 21140
rect 31665 21131 31723 21137
rect 31665 21128 31677 21131
rect 31260 21100 31677 21128
rect 31260 21088 31266 21100
rect 31665 21097 31677 21100
rect 31711 21097 31723 21131
rect 31665 21091 31723 21097
rect 29454 21060 29460 21072
rect 28966 21032 29460 21060
rect 24397 21023 24455 21029
rect 29454 21020 29460 21032
rect 29512 21020 29518 21072
rect 18693 20955 18751 20961
rect 18800 20964 19104 20992
rect 9858 20924 9864 20936
rect 9600 20896 9864 20924
rect 9858 20884 9864 20896
rect 9916 20884 9922 20936
rect 11609 20927 11667 20933
rect 11609 20893 11621 20927
rect 11655 20924 11667 20927
rect 12158 20924 12164 20936
rect 11655 20896 12164 20924
rect 11655 20893 11667 20896
rect 11609 20887 11667 20893
rect 12158 20884 12164 20896
rect 12216 20924 12222 20936
rect 12342 20924 12348 20936
rect 12216 20896 12348 20924
rect 12216 20884 12222 20896
rect 12342 20884 12348 20896
rect 12400 20884 12406 20936
rect 14090 20884 14096 20936
rect 14148 20924 14154 20936
rect 15381 20927 15439 20933
rect 15381 20924 15393 20927
rect 14148 20896 15393 20924
rect 14148 20884 14154 20896
rect 15381 20893 15393 20896
rect 15427 20893 15439 20927
rect 15381 20887 15439 20893
rect 17678 20884 17684 20936
rect 17736 20924 17742 20936
rect 18800 20924 18828 20964
rect 19334 20952 19340 21004
rect 19392 20992 19398 21004
rect 20165 20995 20223 21001
rect 20165 20992 20177 20995
rect 19392 20964 20177 20992
rect 19392 20952 19398 20964
rect 20165 20961 20177 20964
rect 20211 20961 20223 20995
rect 20165 20955 20223 20961
rect 23201 20995 23259 21001
rect 23201 20961 23213 20995
rect 23247 20992 23259 20995
rect 23474 20992 23480 21004
rect 23247 20964 23480 20992
rect 23247 20961 23259 20964
rect 23201 20955 23259 20961
rect 23474 20952 23480 20964
rect 23532 20992 23538 21004
rect 23532 20964 24624 20992
rect 23532 20952 23538 20964
rect 17736 20896 18828 20924
rect 19981 20927 20039 20933
rect 17736 20884 17742 20896
rect 19981 20893 19993 20927
rect 20027 20924 20039 20927
rect 20438 20924 20444 20936
rect 20027 20896 20444 20924
rect 20027 20893 20039 20896
rect 19981 20887 20039 20893
rect 20438 20884 20444 20896
rect 20496 20884 20502 20936
rect 23842 20884 23848 20936
rect 23900 20884 23906 20936
rect 23937 20927 23995 20933
rect 23937 20893 23949 20927
rect 23983 20924 23995 20927
rect 24213 20927 24271 20933
rect 23983 20896 24164 20924
rect 23983 20893 23995 20896
rect 23937 20887 23995 20893
rect 4614 20816 4620 20868
rect 4672 20856 4678 20868
rect 6273 20859 6331 20865
rect 6273 20856 6285 20859
rect 4672 20828 6285 20856
rect 4672 20816 4678 20828
rect 6273 20825 6285 20828
rect 6319 20825 6331 20859
rect 6273 20819 6331 20825
rect 7377 20859 7435 20865
rect 7377 20825 7389 20859
rect 7423 20856 7435 20859
rect 7650 20856 7656 20868
rect 7423 20828 7656 20856
rect 7423 20825 7435 20828
rect 7377 20819 7435 20825
rect 7650 20816 7656 20828
rect 7708 20856 7714 20868
rect 8018 20856 8024 20868
rect 7708 20828 8024 20856
rect 7708 20816 7714 20828
rect 8018 20816 8024 20828
rect 8076 20816 8082 20868
rect 10036 20859 10094 20865
rect 10036 20825 10048 20859
rect 10082 20856 10094 20859
rect 10318 20856 10324 20868
rect 10082 20828 10324 20856
rect 10082 20825 10094 20828
rect 10036 20819 10094 20825
rect 10318 20816 10324 20828
rect 10376 20816 10382 20868
rect 11876 20859 11934 20865
rect 11876 20825 11888 20859
rect 11922 20856 11934 20859
rect 12434 20856 12440 20868
rect 11922 20828 12440 20856
rect 11922 20825 11934 20828
rect 11876 20819 11934 20825
rect 12434 20816 12440 20828
rect 12492 20816 12498 20868
rect 14550 20816 14556 20868
rect 14608 20856 14614 20868
rect 15473 20859 15531 20865
rect 15473 20856 15485 20859
rect 14608 20828 15485 20856
rect 14608 20816 14614 20828
rect 15473 20825 15485 20828
rect 15519 20825 15531 20859
rect 15473 20819 15531 20825
rect 17310 20816 17316 20868
rect 17368 20856 17374 20868
rect 17589 20859 17647 20865
rect 17589 20856 17601 20859
rect 17368 20828 17601 20856
rect 17368 20816 17374 20828
rect 17589 20825 17601 20828
rect 17635 20856 17647 20859
rect 20530 20856 20536 20868
rect 17635 20828 20536 20856
rect 17635 20825 17647 20828
rect 17589 20819 17647 20825
rect 20530 20816 20536 20828
rect 20588 20816 20594 20868
rect 20622 20816 20628 20868
rect 20680 20856 20686 20868
rect 20680 20828 22876 20856
rect 20680 20816 20686 20828
rect 6362 20748 6368 20800
rect 6420 20788 6426 20800
rect 6641 20791 6699 20797
rect 6641 20788 6653 20791
rect 6420 20760 6653 20788
rect 6420 20748 6426 20760
rect 6641 20757 6653 20760
rect 6687 20757 6699 20791
rect 6641 20751 6699 20757
rect 8938 20748 8944 20800
rect 8996 20748 9002 20800
rect 9306 20748 9312 20800
rect 9364 20748 9370 20800
rect 9398 20748 9404 20800
rect 9456 20748 9462 20800
rect 11146 20748 11152 20800
rect 11204 20748 11210 20800
rect 12989 20791 13047 20797
rect 12989 20757 13001 20791
rect 13035 20788 13047 20791
rect 13446 20788 13452 20800
rect 13035 20760 13452 20788
rect 13035 20757 13047 20760
rect 12989 20751 13047 20757
rect 13446 20748 13452 20760
rect 13504 20748 13510 20800
rect 18509 20791 18567 20797
rect 18509 20757 18521 20791
rect 18555 20788 18567 20791
rect 18690 20788 18696 20800
rect 18555 20760 18696 20788
rect 18555 20757 18567 20760
rect 18509 20751 18567 20757
rect 18690 20748 18696 20760
rect 18748 20748 18754 20800
rect 19334 20748 19340 20800
rect 19392 20788 19398 20800
rect 19429 20791 19487 20797
rect 19429 20788 19441 20791
rect 19392 20760 19441 20788
rect 19392 20748 19398 20760
rect 19429 20757 19441 20760
rect 19475 20757 19487 20791
rect 19429 20751 19487 20757
rect 20070 20748 20076 20800
rect 20128 20748 20134 20800
rect 21821 20791 21879 20797
rect 21821 20757 21833 20791
rect 21867 20788 21879 20791
rect 22738 20788 22744 20800
rect 21867 20760 22744 20788
rect 21867 20757 21879 20760
rect 21821 20751 21879 20757
rect 22738 20748 22744 20760
rect 22796 20748 22802 20800
rect 22848 20788 22876 20828
rect 22922 20816 22928 20868
rect 22980 20865 22986 20868
rect 22980 20819 22992 20865
rect 23860 20856 23888 20884
rect 23584 20828 23888 20856
rect 24029 20859 24087 20865
rect 22980 20816 22986 20819
rect 23584 20788 23612 20828
rect 24029 20825 24041 20859
rect 24075 20825 24087 20859
rect 24136 20856 24164 20896
rect 24213 20893 24225 20927
rect 24259 20924 24271 20927
rect 24302 20924 24308 20936
rect 24259 20896 24308 20924
rect 24259 20893 24271 20896
rect 24213 20887 24271 20893
rect 24302 20884 24308 20896
rect 24360 20884 24366 20936
rect 24596 20933 24624 20964
rect 27062 20952 27068 21004
rect 27120 20992 27126 21004
rect 27525 20995 27583 21001
rect 27525 20992 27537 20995
rect 27120 20964 27537 20992
rect 27120 20952 27126 20964
rect 27525 20961 27537 20964
rect 27571 20961 27583 20995
rect 29638 20992 29644 21004
rect 27525 20955 27583 20961
rect 29012 20964 29644 20992
rect 24581 20927 24639 20933
rect 24581 20893 24593 20927
rect 24627 20924 24639 20927
rect 25222 20924 25228 20936
rect 24627 20896 25228 20924
rect 24627 20893 24639 20896
rect 24581 20887 24639 20893
rect 25222 20884 25228 20896
rect 25280 20924 25286 20936
rect 26053 20927 26111 20933
rect 26053 20924 26065 20927
rect 25280 20896 26065 20924
rect 25280 20884 25286 20896
rect 26053 20893 26065 20896
rect 26099 20893 26111 20927
rect 27540 20924 27568 20955
rect 29012 20924 29040 20964
rect 29638 20952 29644 20964
rect 29696 20952 29702 21004
rect 27540 20896 29040 20924
rect 29089 20927 29147 20933
rect 26053 20887 26111 20893
rect 29089 20893 29101 20927
rect 29135 20924 29147 20927
rect 29454 20924 29460 20936
rect 29135 20896 29460 20924
rect 29135 20893 29147 20896
rect 29089 20887 29147 20893
rect 29454 20884 29460 20896
rect 29512 20924 29518 20936
rect 29730 20924 29736 20936
rect 29512 20896 29736 20924
rect 29512 20884 29518 20896
rect 29730 20884 29736 20896
rect 29788 20884 29794 20936
rect 29914 20933 29920 20936
rect 29908 20924 29920 20933
rect 29875 20896 29920 20924
rect 29908 20887 29920 20896
rect 29914 20884 29920 20887
rect 29972 20884 29978 20936
rect 31389 20927 31447 20933
rect 31389 20893 31401 20927
rect 31435 20924 31447 20927
rect 34517 20927 34575 20933
rect 31435 20896 31469 20924
rect 31435 20893 31447 20896
rect 31389 20887 31447 20893
rect 34517 20893 34529 20927
rect 34563 20924 34575 20927
rect 34698 20924 34704 20936
rect 34563 20896 34704 20924
rect 34563 20893 34575 20896
rect 34517 20887 34575 20893
rect 24848 20859 24906 20865
rect 24136 20828 24808 20856
rect 24029 20819 24087 20825
rect 22848 20760 23612 20788
rect 23658 20748 23664 20800
rect 23716 20748 23722 20800
rect 24044 20788 24072 20819
rect 24302 20788 24308 20800
rect 24044 20760 24308 20788
rect 24302 20748 24308 20760
rect 24360 20748 24366 20800
rect 24780 20788 24808 20828
rect 24848 20825 24860 20859
rect 24894 20856 24906 20859
rect 24946 20856 24952 20868
rect 24894 20828 24952 20856
rect 24894 20825 24906 20828
rect 24848 20819 24906 20825
rect 24946 20816 24952 20828
rect 25004 20816 25010 20868
rect 25038 20816 25044 20868
rect 25096 20856 25102 20868
rect 25682 20856 25688 20868
rect 25096 20828 25688 20856
rect 25096 20816 25102 20828
rect 25682 20816 25688 20828
rect 25740 20816 25746 20868
rect 26320 20859 26378 20865
rect 26320 20825 26332 20859
rect 26366 20856 26378 20859
rect 26970 20856 26976 20868
rect 26366 20828 26976 20856
rect 26366 20825 26378 20828
rect 26320 20819 26378 20825
rect 26970 20816 26976 20828
rect 27028 20816 27034 20868
rect 27798 20865 27804 20868
rect 27792 20819 27804 20865
rect 27798 20816 27804 20819
rect 27856 20816 27862 20868
rect 31110 20816 31116 20868
rect 31168 20856 31174 20868
rect 31404 20856 31432 20887
rect 34698 20884 34704 20896
rect 34756 20884 34762 20936
rect 31481 20859 31539 20865
rect 31481 20856 31493 20859
rect 31168 20828 31493 20856
rect 31168 20816 31174 20828
rect 31481 20825 31493 20828
rect 31527 20856 31539 20859
rect 31570 20856 31576 20868
rect 31527 20828 31576 20856
rect 31527 20825 31539 20828
rect 31481 20819 31539 20825
rect 31570 20816 31576 20828
rect 31628 20816 31634 20868
rect 34241 20859 34299 20865
rect 34241 20825 34253 20859
rect 34287 20856 34299 20859
rect 35342 20856 35348 20868
rect 34287 20828 35348 20856
rect 34287 20825 34299 20828
rect 34241 20819 34299 20825
rect 35342 20816 35348 20828
rect 35400 20816 35406 20868
rect 25314 20788 25320 20800
rect 24780 20760 25320 20788
rect 25314 20748 25320 20760
rect 25372 20788 25378 20800
rect 25961 20791 26019 20797
rect 25961 20788 25973 20791
rect 25372 20760 25973 20788
rect 25372 20748 25378 20760
rect 25961 20757 25973 20760
rect 26007 20757 26019 20791
rect 25961 20751 26019 20757
rect 26050 20748 26056 20800
rect 26108 20788 26114 20800
rect 27522 20788 27528 20800
rect 26108 20760 27528 20788
rect 26108 20748 26114 20760
rect 27522 20748 27528 20760
rect 27580 20788 27586 20800
rect 28258 20788 28264 20800
rect 27580 20760 28264 20788
rect 27580 20748 27586 20760
rect 28258 20748 28264 20760
rect 28316 20748 28322 20800
rect 28902 20748 28908 20800
rect 28960 20748 28966 20800
rect 1104 20698 35328 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35328 20698
rect 1104 20624 35328 20646
rect 9306 20544 9312 20596
rect 9364 20584 9370 20596
rect 9493 20587 9551 20593
rect 9493 20584 9505 20587
rect 9364 20556 9505 20584
rect 9364 20544 9370 20556
rect 9493 20553 9505 20556
rect 9539 20553 9551 20587
rect 9493 20547 9551 20553
rect 8380 20519 8438 20525
rect 8380 20485 8392 20519
rect 8426 20516 8438 20519
rect 8938 20516 8944 20528
rect 8426 20488 8944 20516
rect 8426 20485 8438 20488
rect 8380 20479 8438 20485
rect 8938 20476 8944 20488
rect 8996 20476 9002 20528
rect 1302 20408 1308 20460
rect 1360 20448 1366 20460
rect 1397 20451 1455 20457
rect 1397 20448 1409 20451
rect 1360 20420 1409 20448
rect 1360 20408 1366 20420
rect 1397 20417 1409 20420
rect 1443 20448 1455 20451
rect 1673 20451 1731 20457
rect 1673 20448 1685 20451
rect 1443 20420 1685 20448
rect 1443 20417 1455 20420
rect 1397 20411 1455 20417
rect 1673 20417 1685 20420
rect 1719 20417 1731 20451
rect 1673 20411 1731 20417
rect 8110 20408 8116 20460
rect 8168 20408 8174 20460
rect 9508 20448 9536 20547
rect 10318 20544 10324 20596
rect 10376 20544 10382 20596
rect 10689 20587 10747 20593
rect 10689 20553 10701 20587
rect 10735 20584 10747 20587
rect 11146 20584 11152 20596
rect 10735 20556 11152 20584
rect 10735 20553 10747 20556
rect 10689 20547 10747 20553
rect 9953 20519 10011 20525
rect 9953 20485 9965 20519
rect 9999 20516 10011 20519
rect 10704 20516 10732 20547
rect 11146 20544 11152 20556
rect 11204 20544 11210 20596
rect 11606 20544 11612 20596
rect 11664 20584 11670 20596
rect 15562 20584 15568 20596
rect 11664 20556 15568 20584
rect 11664 20544 11670 20556
rect 15562 20544 15568 20556
rect 15620 20544 15626 20596
rect 19978 20544 19984 20596
rect 20036 20584 20042 20596
rect 20257 20587 20315 20593
rect 20257 20584 20269 20587
rect 20036 20556 20269 20584
rect 20036 20544 20042 20556
rect 20257 20553 20269 20556
rect 20303 20584 20315 20587
rect 20809 20587 20867 20593
rect 20809 20584 20821 20587
rect 20303 20556 20821 20584
rect 20303 20553 20315 20556
rect 20257 20547 20315 20553
rect 20809 20553 20821 20556
rect 20855 20553 20867 20587
rect 20809 20547 20867 20553
rect 22649 20587 22707 20593
rect 22649 20553 22661 20587
rect 22695 20584 22707 20587
rect 22738 20584 22744 20596
rect 22695 20556 22744 20584
rect 22695 20553 22707 20556
rect 22649 20547 22707 20553
rect 22738 20544 22744 20556
rect 22796 20544 22802 20596
rect 22922 20544 22928 20596
rect 22980 20584 22986 20596
rect 23017 20587 23075 20593
rect 23017 20584 23029 20587
rect 22980 20556 23029 20584
rect 22980 20544 22986 20556
rect 23017 20553 23029 20556
rect 23063 20553 23075 20587
rect 23017 20547 23075 20553
rect 24394 20544 24400 20596
rect 24452 20584 24458 20596
rect 24489 20587 24547 20593
rect 24489 20584 24501 20587
rect 24452 20556 24501 20584
rect 24452 20544 24458 20556
rect 24489 20553 24501 20556
rect 24535 20553 24547 20587
rect 24489 20547 24547 20553
rect 25314 20544 25320 20596
rect 25372 20544 25378 20596
rect 25869 20587 25927 20593
rect 25869 20553 25881 20587
rect 25915 20584 25927 20587
rect 26050 20584 26056 20596
rect 25915 20556 26056 20584
rect 25915 20553 25927 20556
rect 25869 20547 25927 20553
rect 26050 20544 26056 20556
rect 26108 20544 26114 20596
rect 26418 20544 26424 20596
rect 26476 20544 26482 20596
rect 26970 20544 26976 20596
rect 27028 20544 27034 20596
rect 27341 20587 27399 20593
rect 27341 20553 27353 20587
rect 27387 20584 27399 20587
rect 27430 20584 27436 20596
rect 27387 20556 27436 20584
rect 27387 20553 27399 20556
rect 27341 20547 27399 20553
rect 27430 20544 27436 20556
rect 27488 20544 27494 20596
rect 27798 20544 27804 20596
rect 27856 20544 27862 20596
rect 28169 20587 28227 20593
rect 28169 20553 28181 20587
rect 28215 20584 28227 20587
rect 28902 20584 28908 20596
rect 28215 20556 28908 20584
rect 28215 20553 28227 20556
rect 28169 20547 28227 20553
rect 28902 20544 28908 20556
rect 28960 20544 28966 20596
rect 29362 20544 29368 20596
rect 29420 20584 29426 20596
rect 29457 20587 29515 20593
rect 29457 20584 29469 20587
rect 29420 20556 29469 20584
rect 29420 20544 29426 20556
rect 29457 20553 29469 20556
rect 29503 20553 29515 20587
rect 29457 20547 29515 20553
rect 9999 20488 10732 20516
rect 9999 20485 10011 20488
rect 9953 20479 10011 20485
rect 12342 20476 12348 20528
rect 12400 20516 12406 20528
rect 14550 20516 14556 20528
rect 12400 20488 14556 20516
rect 12400 20476 12406 20488
rect 9677 20451 9735 20457
rect 9677 20448 9689 20451
rect 9508 20420 9689 20448
rect 9677 20417 9689 20420
rect 9723 20417 9735 20451
rect 9677 20411 9735 20417
rect 9861 20451 9919 20457
rect 9861 20417 9873 20451
rect 9907 20417 9919 20451
rect 9861 20411 9919 20417
rect 10045 20451 10103 20457
rect 10045 20417 10057 20451
rect 10091 20448 10103 20451
rect 10318 20448 10324 20460
rect 10091 20420 10324 20448
rect 10091 20417 10103 20420
rect 10045 20411 10103 20417
rect 9876 20380 9904 20411
rect 10318 20408 10324 20420
rect 10376 20408 10382 20460
rect 10781 20451 10839 20457
rect 10781 20417 10793 20451
rect 10827 20448 10839 20451
rect 12069 20451 12127 20457
rect 12069 20448 12081 20451
rect 10827 20420 12081 20448
rect 10827 20417 10839 20420
rect 10781 20411 10839 20417
rect 12069 20417 12081 20420
rect 12115 20448 12127 20451
rect 12805 20451 12863 20457
rect 12115 20420 12756 20448
rect 12115 20417 12127 20420
rect 12069 20411 12127 20417
rect 10410 20380 10416 20392
rect 9876 20352 10416 20380
rect 1581 20247 1639 20253
rect 1581 20213 1593 20247
rect 1627 20244 1639 20247
rect 3786 20244 3792 20256
rect 1627 20216 3792 20244
rect 1627 20213 1639 20216
rect 1581 20207 1639 20213
rect 3786 20204 3792 20216
rect 3844 20204 3850 20256
rect 5534 20204 5540 20256
rect 5592 20244 5598 20256
rect 9876 20244 9904 20352
rect 10410 20340 10416 20352
rect 10468 20340 10474 20392
rect 10965 20383 11023 20389
rect 10965 20349 10977 20383
rect 11011 20380 11023 20383
rect 11011 20352 11284 20380
rect 11011 20349 11023 20352
rect 10965 20343 11023 20349
rect 5592 20216 9904 20244
rect 5592 20204 5598 20216
rect 10226 20204 10232 20256
rect 10284 20204 10290 20256
rect 11256 20253 11284 20352
rect 12342 20340 12348 20392
rect 12400 20340 12406 20392
rect 12728 20380 12756 20420
rect 12805 20417 12817 20451
rect 12851 20448 12863 20451
rect 13446 20448 13452 20460
rect 12851 20420 13452 20448
rect 12851 20417 12863 20420
rect 12805 20411 12863 20417
rect 13446 20408 13452 20420
rect 13504 20408 13510 20460
rect 13556 20457 13584 20488
rect 14550 20476 14556 20488
rect 14608 20476 14614 20528
rect 20717 20519 20775 20525
rect 20717 20516 20729 20519
rect 20180 20488 20729 20516
rect 13541 20451 13599 20457
rect 13541 20417 13553 20451
rect 13587 20417 13599 20451
rect 13541 20411 13599 20417
rect 13808 20451 13866 20457
rect 13808 20417 13820 20451
rect 13854 20448 13866 20451
rect 14090 20448 14096 20460
rect 13854 20420 14096 20448
rect 13854 20417 13866 20420
rect 13808 20411 13866 20417
rect 14090 20408 14096 20420
rect 14148 20408 14154 20460
rect 17034 20408 17040 20460
rect 17092 20408 17098 20460
rect 20180 20457 20208 20488
rect 20717 20485 20729 20488
rect 20763 20516 20775 20519
rect 22094 20516 22100 20528
rect 20763 20488 22100 20516
rect 20763 20485 20775 20488
rect 20717 20479 20775 20485
rect 22094 20476 22100 20488
rect 22152 20476 22158 20528
rect 23750 20476 23756 20528
rect 23808 20516 23814 20528
rect 25409 20519 25467 20525
rect 25409 20516 25421 20519
rect 23808 20488 25421 20516
rect 23808 20476 23814 20488
rect 25409 20485 25421 20488
rect 25455 20516 25467 20519
rect 27890 20516 27896 20528
rect 25455 20488 27896 20516
rect 25455 20485 25467 20488
rect 25409 20479 25467 20485
rect 27890 20476 27896 20488
rect 27948 20516 27954 20528
rect 28261 20519 28319 20525
rect 28261 20516 28273 20519
rect 27948 20488 28273 20516
rect 27948 20476 27954 20488
rect 28261 20485 28273 20488
rect 28307 20516 28319 20519
rect 28718 20516 28724 20528
rect 28307 20488 28724 20516
rect 28307 20485 28319 20488
rect 28261 20479 28319 20485
rect 28718 20476 28724 20488
rect 28776 20476 28782 20528
rect 20165 20451 20223 20457
rect 20165 20417 20177 20451
rect 20211 20417 20223 20451
rect 20165 20411 20223 20417
rect 22557 20451 22615 20457
rect 22557 20417 22569 20451
rect 22603 20448 22615 20451
rect 22646 20448 22652 20460
rect 22603 20420 22652 20448
rect 22603 20417 22615 20420
rect 22557 20411 22615 20417
rect 22646 20408 22652 20420
rect 22704 20408 22710 20460
rect 24026 20408 24032 20460
rect 24084 20408 24090 20460
rect 24210 20408 24216 20460
rect 24268 20448 24274 20460
rect 24305 20451 24363 20457
rect 24305 20448 24317 20451
rect 24268 20420 24317 20448
rect 24268 20408 24274 20420
rect 24305 20417 24317 20420
rect 24351 20417 24363 20451
rect 24305 20411 24363 20417
rect 26602 20408 26608 20460
rect 26660 20448 26666 20460
rect 29472 20448 29500 20547
rect 32214 20476 32220 20528
rect 32272 20516 32278 20528
rect 33502 20516 33508 20528
rect 32272 20488 33508 20516
rect 32272 20476 32278 20488
rect 33502 20476 33508 20488
rect 33560 20516 33566 20528
rect 33560 20488 33994 20516
rect 33560 20476 33566 20488
rect 29641 20451 29699 20457
rect 29641 20448 29653 20451
rect 26660 20420 27568 20448
rect 29472 20420 29653 20448
rect 26660 20408 26666 20420
rect 12894 20380 12900 20392
rect 12728 20352 12900 20380
rect 12894 20340 12900 20352
rect 12952 20340 12958 20392
rect 12986 20340 12992 20392
rect 13044 20380 13050 20392
rect 13081 20383 13139 20389
rect 13081 20380 13093 20383
rect 13044 20352 13093 20380
rect 13044 20340 13050 20352
rect 13081 20349 13093 20352
rect 13127 20380 13139 20383
rect 13265 20383 13323 20389
rect 13265 20380 13277 20383
rect 13127 20352 13277 20380
rect 13127 20349 13139 20352
rect 13081 20343 13139 20349
rect 13265 20349 13277 20352
rect 13311 20349 13323 20383
rect 13265 20343 13323 20349
rect 15930 20340 15936 20392
rect 15988 20380 15994 20392
rect 17129 20383 17187 20389
rect 17129 20380 17141 20383
rect 15988 20352 17141 20380
rect 15988 20340 15994 20352
rect 17129 20349 17141 20352
rect 17175 20349 17187 20383
rect 17129 20343 17187 20349
rect 17218 20340 17224 20392
rect 17276 20380 17282 20392
rect 17497 20383 17555 20389
rect 17497 20380 17509 20383
rect 17276 20352 17509 20380
rect 17276 20340 17282 20352
rect 17497 20349 17509 20352
rect 17543 20349 17555 20383
rect 17497 20343 17555 20349
rect 22189 20383 22247 20389
rect 22189 20349 22201 20383
rect 22235 20380 22247 20383
rect 22462 20380 22468 20392
rect 22235 20352 22468 20380
rect 22235 20349 22247 20352
rect 22189 20343 22247 20349
rect 22462 20340 22468 20352
rect 22520 20340 22526 20392
rect 24118 20340 24124 20392
rect 24176 20340 24182 20392
rect 24946 20340 24952 20392
rect 25004 20340 25010 20392
rect 25593 20383 25651 20389
rect 25593 20349 25605 20383
rect 25639 20380 25651 20383
rect 26050 20380 26056 20392
rect 25639 20352 26056 20380
rect 25639 20349 25651 20352
rect 25593 20343 25651 20349
rect 26050 20340 26056 20352
rect 26108 20340 26114 20392
rect 26418 20340 26424 20392
rect 26476 20380 26482 20392
rect 27540 20389 27568 20420
rect 29641 20417 29653 20420
rect 29687 20417 29699 20451
rect 29641 20411 29699 20417
rect 29822 20408 29828 20460
rect 29880 20408 29886 20460
rect 30193 20451 30251 20457
rect 30193 20417 30205 20451
rect 30239 20448 30251 20451
rect 30282 20448 30288 20460
rect 30239 20420 30288 20448
rect 30239 20417 30251 20420
rect 30193 20411 30251 20417
rect 30282 20408 30288 20420
rect 30340 20408 30346 20460
rect 30745 20451 30803 20457
rect 30745 20417 30757 20451
rect 30791 20448 30803 20451
rect 30791 20420 31340 20448
rect 30791 20417 30803 20420
rect 30745 20411 30803 20417
rect 27433 20383 27491 20389
rect 27433 20380 27445 20383
rect 26476 20352 27445 20380
rect 26476 20340 26482 20352
rect 27433 20349 27445 20352
rect 27479 20349 27491 20383
rect 27433 20343 27491 20349
rect 27525 20383 27583 20389
rect 27525 20349 27537 20383
rect 27571 20349 27583 20383
rect 27525 20343 27583 20349
rect 28350 20340 28356 20392
rect 28408 20340 28414 20392
rect 29917 20383 29975 20389
rect 29917 20349 29929 20383
rect 29963 20349 29975 20383
rect 29917 20343 29975 20349
rect 30009 20383 30067 20389
rect 30009 20349 30021 20383
rect 30055 20349 30067 20383
rect 30009 20343 30067 20349
rect 12434 20272 12440 20324
rect 12492 20272 12498 20324
rect 15838 20312 15844 20324
rect 13188 20284 13584 20312
rect 11241 20247 11299 20253
rect 11241 20213 11253 20247
rect 11287 20244 11299 20247
rect 13188 20244 13216 20284
rect 11287 20216 13216 20244
rect 13556 20244 13584 20284
rect 14568 20284 15844 20312
rect 14568 20244 14596 20284
rect 15838 20272 15844 20284
rect 15896 20272 15902 20324
rect 19426 20272 19432 20324
rect 19484 20312 19490 20324
rect 20533 20315 20591 20321
rect 20533 20312 20545 20315
rect 19484 20284 20545 20312
rect 19484 20272 19490 20284
rect 20533 20281 20545 20284
rect 20579 20312 20591 20315
rect 20579 20284 20944 20312
rect 20579 20281 20591 20284
rect 20533 20275 20591 20281
rect 13556 20216 14596 20244
rect 11287 20213 11299 20216
rect 11241 20207 11299 20213
rect 14642 20204 14648 20256
rect 14700 20244 14706 20256
rect 14921 20247 14979 20253
rect 14921 20244 14933 20247
rect 14700 20216 14933 20244
rect 14700 20204 14706 20216
rect 14921 20213 14933 20216
rect 14967 20213 14979 20247
rect 14921 20207 14979 20213
rect 16666 20204 16672 20256
rect 16724 20204 16730 20256
rect 20916 20244 20944 20284
rect 23566 20244 23572 20256
rect 20916 20216 23572 20244
rect 23566 20204 23572 20216
rect 23624 20204 23630 20256
rect 23658 20204 23664 20256
rect 23716 20244 23722 20256
rect 24029 20247 24087 20253
rect 24029 20244 24041 20247
rect 23716 20216 24041 20244
rect 23716 20204 23722 20216
rect 24029 20213 24041 20216
rect 24075 20213 24087 20247
rect 24029 20207 24087 20213
rect 24302 20204 24308 20256
rect 24360 20244 24366 20256
rect 24673 20247 24731 20253
rect 24673 20244 24685 20247
rect 24360 20216 24685 20244
rect 24360 20204 24366 20216
rect 24673 20213 24685 20216
rect 24719 20244 24731 20247
rect 24854 20244 24860 20256
rect 24719 20216 24860 20244
rect 24719 20213 24731 20216
rect 24673 20207 24731 20213
rect 24854 20204 24860 20216
rect 24912 20204 24918 20256
rect 24964 20253 24992 20340
rect 26602 20272 26608 20324
rect 26660 20272 26666 20324
rect 26786 20272 26792 20324
rect 26844 20312 26850 20324
rect 29932 20312 29960 20343
rect 26844 20284 29960 20312
rect 30024 20312 30052 20343
rect 30561 20315 30619 20321
rect 30561 20312 30573 20315
rect 30024 20284 30573 20312
rect 26844 20272 26850 20284
rect 24949 20247 25007 20253
rect 24949 20213 24961 20247
rect 24995 20213 25007 20247
rect 24949 20207 25007 20213
rect 27798 20204 27804 20256
rect 27856 20244 27862 20256
rect 30024 20244 30052 20284
rect 30561 20281 30573 20284
rect 30607 20312 30619 20315
rect 30837 20315 30895 20321
rect 30837 20312 30849 20315
rect 30607 20284 30849 20312
rect 30607 20281 30619 20284
rect 30561 20275 30619 20281
rect 30837 20281 30849 20284
rect 30883 20312 30895 20315
rect 31021 20315 31079 20321
rect 31021 20312 31033 20315
rect 30883 20284 31033 20312
rect 30883 20281 30895 20284
rect 30837 20275 30895 20281
rect 31021 20281 31033 20284
rect 31067 20281 31079 20315
rect 31021 20275 31079 20281
rect 27856 20216 30052 20244
rect 27856 20204 27862 20216
rect 30374 20204 30380 20256
rect 30432 20204 30438 20256
rect 31312 20253 31340 20420
rect 33134 20408 33140 20460
rect 33192 20448 33198 20460
rect 33229 20451 33287 20457
rect 33229 20448 33241 20451
rect 33192 20420 33241 20448
rect 33192 20408 33198 20420
rect 33229 20417 33241 20420
rect 33275 20417 33287 20451
rect 33229 20411 33287 20417
rect 33505 20383 33563 20389
rect 33505 20349 33517 20383
rect 33551 20380 33563 20383
rect 33962 20380 33968 20392
rect 33551 20352 33968 20380
rect 33551 20349 33563 20352
rect 33505 20343 33563 20349
rect 33962 20340 33968 20352
rect 34020 20340 34026 20392
rect 31297 20247 31355 20253
rect 31297 20213 31309 20247
rect 31343 20244 31355 20247
rect 31386 20244 31392 20256
rect 31343 20216 31392 20244
rect 31343 20213 31355 20216
rect 31297 20207 31355 20213
rect 31386 20204 31392 20216
rect 31444 20204 31450 20256
rect 34698 20204 34704 20256
rect 34756 20244 34762 20256
rect 34977 20247 35035 20253
rect 34977 20244 34989 20247
rect 34756 20216 34989 20244
rect 34756 20204 34762 20216
rect 34977 20213 34989 20216
rect 35023 20213 35035 20247
rect 34977 20207 35035 20213
rect 1104 20154 35328 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 35328 20154
rect 1104 20080 35328 20102
rect 3973 20043 4031 20049
rect 3973 20040 3985 20043
rect 3436 20012 3985 20040
rect 3436 19845 3464 20012
rect 3973 20009 3985 20012
rect 4019 20040 4031 20043
rect 9674 20040 9680 20052
rect 4019 20012 9680 20040
rect 4019 20009 4031 20012
rect 3973 20003 4031 20009
rect 9674 20000 9680 20012
rect 9732 20000 9738 20052
rect 16758 20040 16764 20052
rect 14835 20012 16764 20040
rect 3605 19975 3663 19981
rect 3605 19941 3617 19975
rect 3651 19972 3663 19975
rect 4154 19972 4160 19984
rect 3651 19944 4160 19972
rect 3651 19941 3663 19944
rect 3605 19935 3663 19941
rect 4154 19932 4160 19944
rect 4212 19932 4218 19984
rect 8478 19932 8484 19984
rect 8536 19972 8542 19984
rect 8536 19944 12434 19972
rect 8536 19932 8542 19944
rect 4798 19864 4804 19916
rect 4856 19864 4862 19916
rect 10410 19864 10416 19916
rect 10468 19904 10474 19916
rect 10505 19907 10563 19913
rect 10505 19904 10517 19907
rect 10468 19876 10517 19904
rect 10468 19864 10474 19876
rect 10505 19873 10517 19876
rect 10551 19873 10563 19907
rect 12406 19904 12434 19944
rect 12526 19932 12532 19984
rect 12584 19972 12590 19984
rect 12894 19972 12900 19984
rect 12584 19944 12900 19972
rect 12584 19932 12590 19944
rect 12894 19932 12900 19944
rect 12952 19972 12958 19984
rect 14835 19972 14863 20012
rect 16758 20000 16764 20012
rect 16816 20000 16822 20052
rect 17034 20000 17040 20052
rect 17092 20040 17098 20052
rect 17129 20043 17187 20049
rect 17129 20040 17141 20043
rect 17092 20012 17141 20040
rect 17092 20000 17098 20012
rect 17129 20009 17141 20012
rect 17175 20009 17187 20043
rect 17129 20003 17187 20009
rect 21913 20043 21971 20049
rect 21913 20009 21925 20043
rect 21959 20040 21971 20043
rect 24026 20040 24032 20052
rect 21959 20012 24032 20040
rect 21959 20009 21971 20012
rect 21913 20003 21971 20009
rect 24026 20000 24032 20012
rect 24084 20000 24090 20052
rect 24489 20043 24547 20049
rect 24489 20009 24501 20043
rect 24535 20040 24547 20043
rect 24854 20040 24860 20052
rect 24535 20012 24860 20040
rect 24535 20009 24547 20012
rect 24489 20003 24547 20009
rect 24854 20000 24860 20012
rect 24912 20000 24918 20052
rect 31849 20043 31907 20049
rect 31849 20009 31861 20043
rect 31895 20040 31907 20043
rect 32030 20040 32036 20052
rect 31895 20012 32036 20040
rect 31895 20009 31907 20012
rect 31849 20003 31907 20009
rect 32030 20000 32036 20012
rect 32088 20040 32094 20052
rect 33410 20040 33416 20052
rect 32088 20012 33416 20040
rect 32088 20000 32094 20012
rect 33410 20000 33416 20012
rect 33468 20000 33474 20052
rect 33962 20000 33968 20052
rect 34020 20000 34026 20052
rect 12952 19944 14863 19972
rect 12952 19932 12958 19944
rect 13906 19904 13912 19916
rect 12406 19876 13912 19904
rect 10505 19867 10563 19873
rect 13906 19864 13912 19876
rect 13964 19864 13970 19916
rect 14559 19904 14587 19944
rect 22094 19932 22100 19984
rect 22152 19972 22158 19984
rect 22152 19944 23336 19972
rect 22152 19932 22158 19944
rect 23308 19916 23336 19944
rect 23566 19932 23572 19984
rect 23624 19972 23630 19984
rect 25590 19972 25596 19984
rect 23624 19944 25596 19972
rect 23624 19932 23630 19944
rect 25590 19932 25596 19944
rect 25648 19932 25654 19984
rect 14476 19876 14587 19904
rect 14737 19907 14795 19913
rect 3421 19839 3479 19845
rect 3421 19805 3433 19839
rect 3467 19805 3479 19839
rect 3421 19799 3479 19805
rect 3786 19796 3792 19848
rect 3844 19796 3850 19848
rect 4430 19796 4436 19848
rect 4488 19836 4494 19848
rect 4709 19839 4767 19845
rect 4709 19836 4721 19839
rect 4488 19808 4721 19836
rect 4488 19796 4494 19808
rect 4709 19805 4721 19808
rect 4755 19836 4767 19839
rect 5442 19836 5448 19848
rect 4755 19808 5448 19836
rect 4755 19805 4767 19808
rect 4709 19799 4767 19805
rect 5442 19796 5448 19808
rect 5500 19796 5506 19848
rect 14476 19845 14504 19876
rect 14737 19873 14749 19907
rect 14783 19904 14795 19907
rect 15010 19904 15016 19916
rect 14783 19876 15016 19904
rect 14783 19873 14795 19876
rect 14737 19867 14795 19873
rect 15010 19864 15016 19876
rect 15068 19864 15074 19916
rect 22281 19907 22339 19913
rect 22281 19904 22293 19907
rect 21468 19876 22293 19904
rect 21468 19848 21496 19876
rect 22281 19873 22293 19876
rect 22327 19904 22339 19907
rect 22327 19876 22600 19904
rect 22327 19873 22339 19876
rect 22281 19867 22339 19873
rect 14461 19839 14519 19845
rect 14461 19805 14473 19839
rect 14507 19805 14519 19839
rect 14461 19799 14519 19805
rect 14550 19796 14556 19848
rect 14608 19836 14614 19848
rect 14918 19836 14924 19848
rect 14608 19808 14924 19836
rect 14608 19796 14614 19808
rect 14918 19796 14924 19808
rect 14976 19836 14982 19848
rect 15749 19839 15807 19845
rect 15749 19836 15761 19839
rect 14976 19808 15761 19836
rect 14976 19796 14982 19808
rect 15749 19805 15761 19808
rect 15795 19836 15807 19839
rect 16574 19836 16580 19848
rect 15795 19808 16580 19836
rect 15795 19805 15807 19808
rect 15749 19799 15807 19805
rect 16574 19796 16580 19808
rect 16632 19836 16638 19848
rect 17681 19839 17739 19845
rect 17681 19836 17693 19839
rect 16632 19808 17693 19836
rect 16632 19796 16638 19808
rect 17681 19805 17693 19808
rect 17727 19805 17739 19839
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 17681 19799 17739 19805
rect 19076 19808 19257 19836
rect 5068 19771 5126 19777
rect 5068 19737 5080 19771
rect 5114 19768 5126 19771
rect 5350 19768 5356 19780
rect 5114 19740 5356 19768
rect 5114 19737 5126 19740
rect 5068 19731 5126 19737
rect 5350 19728 5356 19740
rect 5408 19728 5414 19780
rect 5994 19728 6000 19780
rect 6052 19768 6058 19780
rect 6273 19771 6331 19777
rect 6273 19768 6285 19771
rect 6052 19740 6285 19768
rect 6052 19728 6058 19740
rect 6273 19737 6285 19740
rect 6319 19737 6331 19771
rect 6273 19731 6331 19737
rect 10410 19728 10416 19780
rect 10468 19728 10474 19780
rect 12802 19728 12808 19780
rect 12860 19768 12866 19780
rect 16016 19771 16074 19777
rect 12860 19740 15332 19768
rect 12860 19728 12866 19740
rect 6178 19660 6184 19712
rect 6236 19660 6242 19712
rect 6638 19660 6644 19712
rect 6696 19700 6702 19712
rect 7193 19703 7251 19709
rect 7193 19700 7205 19703
rect 6696 19672 7205 19700
rect 6696 19660 6702 19672
rect 7193 19669 7205 19672
rect 7239 19700 7251 19703
rect 11606 19700 11612 19712
rect 7239 19672 11612 19700
rect 7239 19669 7251 19672
rect 7193 19663 7251 19669
rect 11606 19660 11612 19672
rect 11664 19660 11670 19712
rect 12710 19660 12716 19712
rect 12768 19700 12774 19712
rect 12897 19703 12955 19709
rect 12897 19700 12909 19703
rect 12768 19672 12909 19700
rect 12768 19660 12774 19672
rect 12897 19669 12909 19672
rect 12943 19669 12955 19703
rect 12897 19663 12955 19669
rect 14090 19660 14096 19712
rect 14148 19660 14154 19712
rect 14553 19703 14611 19709
rect 14553 19669 14565 19703
rect 14599 19700 14611 19703
rect 14642 19700 14648 19712
rect 14599 19672 14648 19700
rect 14599 19669 14611 19672
rect 14553 19663 14611 19669
rect 14642 19660 14648 19672
rect 14700 19700 14706 19712
rect 14826 19700 14832 19712
rect 14700 19672 14832 19700
rect 14700 19660 14706 19672
rect 14826 19660 14832 19672
rect 14884 19660 14890 19712
rect 15102 19660 15108 19712
rect 15160 19700 15166 19712
rect 15197 19703 15255 19709
rect 15197 19700 15209 19703
rect 15160 19672 15209 19700
rect 15160 19660 15166 19672
rect 15197 19669 15209 19672
rect 15243 19669 15255 19703
rect 15304 19700 15332 19740
rect 16016 19737 16028 19771
rect 16062 19768 16074 19771
rect 16666 19768 16672 19780
rect 16062 19740 16672 19768
rect 16062 19737 16074 19740
rect 16016 19731 16074 19737
rect 16666 19728 16672 19740
rect 16724 19728 16730 19780
rect 17948 19771 18006 19777
rect 17948 19737 17960 19771
rect 17994 19768 18006 19771
rect 18230 19768 18236 19780
rect 17994 19740 18236 19768
rect 17994 19737 18006 19740
rect 17948 19731 18006 19737
rect 18230 19728 18236 19740
rect 18288 19728 18294 19780
rect 17218 19700 17224 19712
rect 15304 19672 17224 19700
rect 15197 19663 15255 19669
rect 17218 19660 17224 19672
rect 17276 19660 17282 19712
rect 18598 19660 18604 19712
rect 18656 19700 18662 19712
rect 19076 19709 19104 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 19426 19796 19432 19848
rect 19484 19796 19490 19848
rect 19613 19839 19671 19845
rect 19613 19805 19625 19839
rect 19659 19805 19671 19839
rect 19613 19799 19671 19805
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19836 19947 19839
rect 20622 19836 20628 19848
rect 19935 19808 20628 19836
rect 19935 19805 19947 19808
rect 19889 19799 19947 19805
rect 19518 19728 19524 19780
rect 19576 19728 19582 19780
rect 19628 19768 19656 19799
rect 20622 19796 20628 19808
rect 20680 19796 20686 19848
rect 21361 19839 21419 19845
rect 21361 19836 21373 19839
rect 20732 19808 21373 19836
rect 19978 19768 19984 19780
rect 19628 19740 19984 19768
rect 19978 19728 19984 19740
rect 20036 19728 20042 19780
rect 20156 19771 20214 19777
rect 20156 19737 20168 19771
rect 20202 19768 20214 19771
rect 20530 19768 20536 19780
rect 20202 19740 20536 19768
rect 20202 19737 20214 19740
rect 20156 19731 20214 19737
rect 20530 19728 20536 19740
rect 20588 19728 20594 19780
rect 19061 19703 19119 19709
rect 19061 19700 19073 19703
rect 18656 19672 19073 19700
rect 18656 19660 18662 19672
rect 19061 19669 19073 19672
rect 19107 19669 19119 19703
rect 19061 19663 19119 19669
rect 19797 19703 19855 19709
rect 19797 19669 19809 19703
rect 19843 19700 19855 19703
rect 20732 19700 20760 19808
rect 21361 19805 21373 19808
rect 21407 19805 21419 19839
rect 21361 19799 21419 19805
rect 21450 19796 21456 19848
rect 21508 19796 21514 19848
rect 21637 19839 21695 19845
rect 21637 19805 21649 19839
rect 21683 19805 21695 19839
rect 21637 19799 21695 19805
rect 21652 19768 21680 19799
rect 21726 19796 21732 19848
rect 21784 19836 21790 19848
rect 22094 19836 22100 19848
rect 21784 19808 22100 19836
rect 21784 19796 21790 19808
rect 22094 19796 22100 19808
rect 22152 19796 22158 19848
rect 22572 19836 22600 19876
rect 22646 19864 22652 19916
rect 22704 19904 22710 19916
rect 22833 19907 22891 19913
rect 22833 19904 22845 19907
rect 22704 19876 22845 19904
rect 22704 19864 22710 19876
rect 22833 19873 22845 19876
rect 22879 19873 22891 19907
rect 22833 19867 22891 19873
rect 23017 19907 23075 19913
rect 23017 19873 23029 19907
rect 23063 19904 23075 19907
rect 23198 19904 23204 19916
rect 23063 19876 23204 19904
rect 23063 19873 23075 19876
rect 23017 19867 23075 19873
rect 23198 19864 23204 19876
rect 23256 19864 23262 19916
rect 23290 19864 23296 19916
rect 23348 19904 23354 19916
rect 26694 19904 26700 19916
rect 23348 19876 26700 19904
rect 23348 19864 23354 19876
rect 26694 19864 26700 19876
rect 26752 19864 26758 19916
rect 30374 19864 30380 19916
rect 30432 19904 30438 19916
rect 34701 19907 34759 19913
rect 30432 19876 34192 19904
rect 30432 19864 30438 19876
rect 24673 19839 24731 19845
rect 22572 19808 23980 19836
rect 21284 19740 21680 19768
rect 21284 19712 21312 19740
rect 23842 19728 23848 19780
rect 23900 19728 23906 19780
rect 23952 19768 23980 19808
rect 24673 19805 24685 19839
rect 24719 19836 24731 19839
rect 26142 19836 26148 19848
rect 24719 19808 26148 19836
rect 24719 19805 24731 19808
rect 24673 19799 24731 19805
rect 26142 19796 26148 19808
rect 26200 19796 26206 19848
rect 30745 19839 30803 19845
rect 30745 19805 30757 19839
rect 30791 19836 30803 19839
rect 32490 19836 32496 19848
rect 30791 19808 32496 19836
rect 30791 19805 30803 19808
rect 30745 19799 30803 19805
rect 32490 19796 32496 19808
rect 32548 19796 32554 19848
rect 34164 19845 34192 19876
rect 34701 19873 34713 19907
rect 34747 19873 34759 19907
rect 34701 19867 34759 19873
rect 34149 19839 34207 19845
rect 34149 19805 34161 19839
rect 34195 19805 34207 19839
rect 34149 19799 34207 19805
rect 34238 19796 34244 19848
rect 34296 19836 34302 19848
rect 34425 19839 34483 19845
rect 34425 19836 34437 19839
rect 34296 19808 34437 19836
rect 34296 19796 34302 19808
rect 34425 19805 34437 19808
rect 34471 19836 34483 19839
rect 34716 19836 34744 19867
rect 34471 19808 34744 19836
rect 34471 19805 34483 19808
rect 34425 19799 34483 19805
rect 25958 19768 25964 19780
rect 23952 19740 25964 19768
rect 25958 19728 25964 19740
rect 26016 19728 26022 19780
rect 32030 19728 32036 19780
rect 32088 19728 32094 19780
rect 32214 19728 32220 19780
rect 32272 19728 32278 19780
rect 34333 19771 34391 19777
rect 34333 19737 34345 19771
rect 34379 19768 34391 19771
rect 34698 19768 34704 19780
rect 34379 19740 34704 19768
rect 34379 19737 34391 19740
rect 34333 19731 34391 19737
rect 34698 19728 34704 19740
rect 34756 19728 34762 19780
rect 34882 19728 34888 19780
rect 34940 19728 34946 19780
rect 19843 19672 20760 19700
rect 19843 19669 19855 19672
rect 19797 19663 19855 19669
rect 21266 19660 21272 19712
rect 21324 19660 21330 19712
rect 22370 19660 22376 19712
rect 22428 19660 22434 19712
rect 22738 19660 22744 19712
rect 22796 19660 22802 19712
rect 23198 19660 23204 19712
rect 23256 19660 23262 19712
rect 23658 19660 23664 19712
rect 23716 19700 23722 19712
rect 23753 19703 23811 19709
rect 23753 19700 23765 19703
rect 23716 19672 23765 19700
rect 23716 19660 23722 19672
rect 23753 19669 23765 19672
rect 23799 19700 23811 19703
rect 24026 19700 24032 19712
rect 23799 19672 24032 19700
rect 23799 19669 23811 19672
rect 23753 19663 23811 19669
rect 24026 19660 24032 19672
rect 24084 19660 24090 19712
rect 26694 19660 26700 19712
rect 26752 19700 26758 19712
rect 26970 19700 26976 19712
rect 26752 19672 26976 19700
rect 26752 19660 26758 19672
rect 26970 19660 26976 19672
rect 27028 19660 27034 19712
rect 27709 19703 27767 19709
rect 27709 19669 27721 19703
rect 27755 19700 27767 19703
rect 28350 19700 28356 19712
rect 27755 19672 28356 19700
rect 27755 19669 27767 19672
rect 27709 19663 27767 19669
rect 28350 19660 28356 19672
rect 28408 19660 28414 19712
rect 30466 19660 30472 19712
rect 30524 19700 30530 19712
rect 30561 19703 30619 19709
rect 30561 19700 30573 19703
rect 30524 19672 30573 19700
rect 30524 19660 30530 19672
rect 30561 19669 30573 19672
rect 30607 19669 30619 19703
rect 30561 19663 30619 19669
rect 1104 19610 35328 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35328 19610
rect 1104 19536 35328 19558
rect 3789 19499 3847 19505
rect 3789 19465 3801 19499
rect 3835 19465 3847 19499
rect 3789 19459 3847 19465
rect 5169 19499 5227 19505
rect 5169 19465 5181 19499
rect 5215 19465 5227 19499
rect 5169 19459 5227 19465
rect 3510 19428 3516 19440
rect 2332 19400 3516 19428
rect 2332 19369 2360 19400
rect 3510 19388 3516 19400
rect 3568 19388 3574 19440
rect 2317 19363 2375 19369
rect 2317 19329 2329 19363
rect 2363 19329 2375 19363
rect 2317 19323 2375 19329
rect 2584 19363 2642 19369
rect 2584 19329 2596 19363
rect 2630 19360 2642 19363
rect 3804 19360 3832 19459
rect 4154 19388 4160 19440
rect 4212 19428 4218 19440
rect 4212 19400 5120 19428
rect 4212 19388 4218 19400
rect 4617 19363 4675 19369
rect 4617 19360 4629 19363
rect 2630 19332 3832 19360
rect 4264 19332 4629 19360
rect 2630 19329 2642 19332
rect 2584 19323 2642 19329
rect 4264 19301 4292 19332
rect 4617 19329 4629 19332
rect 4663 19329 4675 19363
rect 4617 19323 4675 19329
rect 4801 19363 4859 19369
rect 4801 19329 4813 19363
rect 4847 19329 4859 19363
rect 4801 19323 4859 19329
rect 4249 19295 4307 19301
rect 4249 19261 4261 19295
rect 4295 19261 4307 19295
rect 4249 19255 4307 19261
rect 3697 19227 3755 19233
rect 3697 19193 3709 19227
rect 3743 19224 3755 19227
rect 4264 19224 4292 19255
rect 4430 19252 4436 19304
rect 4488 19252 4494 19304
rect 3743 19196 4292 19224
rect 4816 19224 4844 19323
rect 4890 19320 4896 19372
rect 4948 19320 4954 19372
rect 4982 19320 4988 19372
rect 5040 19320 5046 19372
rect 5092 19292 5120 19400
rect 5184 19360 5212 19459
rect 5350 19456 5356 19508
rect 5408 19456 5414 19508
rect 5442 19456 5448 19508
rect 5500 19496 5506 19508
rect 5813 19499 5871 19505
rect 5813 19496 5825 19499
rect 5500 19468 5825 19496
rect 5500 19456 5506 19468
rect 5813 19465 5825 19468
rect 5859 19465 5871 19499
rect 5813 19459 5871 19465
rect 10505 19499 10563 19505
rect 10505 19465 10517 19499
rect 10551 19496 10563 19499
rect 12802 19496 12808 19508
rect 10551 19468 12808 19496
rect 10551 19465 10563 19468
rect 10505 19459 10563 19465
rect 12802 19456 12808 19468
rect 12860 19456 12866 19508
rect 12897 19499 12955 19505
rect 12897 19465 12909 19499
rect 12943 19465 12955 19499
rect 12897 19459 12955 19465
rect 14093 19499 14151 19505
rect 14093 19465 14105 19499
rect 14139 19496 14151 19499
rect 14274 19496 14280 19508
rect 14139 19468 14280 19496
rect 14139 19465 14151 19468
rect 14093 19459 14151 19465
rect 5721 19431 5779 19437
rect 5721 19397 5733 19431
rect 5767 19428 5779 19431
rect 6178 19428 6184 19440
rect 5767 19400 6184 19428
rect 5767 19397 5779 19400
rect 5721 19391 5779 19397
rect 6178 19388 6184 19400
rect 6236 19428 6242 19440
rect 6236 19400 6500 19428
rect 6236 19388 6242 19400
rect 6472 19369 6500 19400
rect 6638 19388 6644 19440
rect 6696 19388 6702 19440
rect 6733 19431 6791 19437
rect 6733 19397 6745 19431
rect 6779 19428 6791 19431
rect 7006 19428 7012 19440
rect 6779 19400 7012 19428
rect 6779 19397 6791 19400
rect 6733 19391 6791 19397
rect 7006 19388 7012 19400
rect 7064 19388 7070 19440
rect 10045 19431 10103 19437
rect 7576 19400 9352 19428
rect 6365 19363 6423 19369
rect 6365 19360 6377 19363
rect 5184 19332 6377 19360
rect 6365 19329 6377 19332
rect 6411 19329 6423 19363
rect 6365 19323 6423 19329
rect 6458 19363 6516 19369
rect 6458 19329 6470 19363
rect 6504 19329 6516 19363
rect 6458 19323 6516 19329
rect 6871 19363 6929 19369
rect 6871 19329 6883 19363
rect 6917 19329 6929 19363
rect 7576 19360 7604 19400
rect 6871 19323 6929 19329
rect 7024 19332 7604 19360
rect 7644 19363 7702 19369
rect 5442 19292 5448 19304
rect 5092 19264 5448 19292
rect 5442 19252 5448 19264
rect 5500 19252 5506 19304
rect 5994 19252 6000 19304
rect 6052 19252 6058 19304
rect 5350 19224 5356 19236
rect 4816 19196 5356 19224
rect 3743 19193 3755 19196
rect 3697 19187 3755 19193
rect 5350 19184 5356 19196
rect 5408 19184 5414 19236
rect 6886 19156 6914 19323
rect 7024 19233 7052 19332
rect 7644 19329 7656 19363
rect 7690 19360 7702 19363
rect 7926 19360 7932 19372
rect 7690 19332 7932 19360
rect 7690 19329 7702 19332
rect 7644 19323 7702 19329
rect 7926 19320 7932 19332
rect 7984 19320 7990 19372
rect 8849 19363 8907 19369
rect 8849 19360 8861 19363
rect 8772 19332 8861 19360
rect 7374 19252 7380 19304
rect 7432 19252 7438 19304
rect 7009 19227 7067 19233
rect 7009 19193 7021 19227
rect 7055 19193 7067 19227
rect 7009 19187 7067 19193
rect 7285 19159 7343 19165
rect 7285 19156 7297 19159
rect 6886 19128 7297 19156
rect 7285 19125 7297 19128
rect 7331 19156 7343 19159
rect 8110 19156 8116 19168
rect 7331 19128 8116 19156
rect 7331 19125 7343 19128
rect 7285 19119 7343 19125
rect 8110 19116 8116 19128
rect 8168 19116 8174 19168
rect 8294 19116 8300 19168
rect 8352 19156 8358 19168
rect 8772 19165 8800 19332
rect 8849 19329 8861 19332
rect 8895 19329 8907 19363
rect 8849 19323 8907 19329
rect 9030 19320 9036 19372
rect 9088 19320 9094 19372
rect 9122 19320 9128 19372
rect 9180 19320 9186 19372
rect 9217 19363 9275 19369
rect 9217 19329 9229 19363
rect 9263 19329 9275 19363
rect 9324 19360 9352 19400
rect 10045 19397 10057 19431
rect 10091 19428 10103 19431
rect 10597 19431 10655 19437
rect 10597 19428 10609 19431
rect 10091 19400 10609 19428
rect 10091 19397 10103 19400
rect 10045 19391 10103 19397
rect 10597 19397 10609 19400
rect 10643 19397 10655 19431
rect 10597 19391 10655 19397
rect 10686 19388 10692 19440
rect 10744 19428 10750 19440
rect 12912 19428 12940 19459
rect 14274 19456 14280 19468
rect 14332 19496 14338 19508
rect 15105 19499 15163 19505
rect 14332 19468 15056 19496
rect 14332 19456 14338 19468
rect 13173 19431 13231 19437
rect 13173 19428 13185 19431
rect 10744 19400 11008 19428
rect 10744 19388 10750 19400
rect 9324 19332 10180 19360
rect 9217 19323 9275 19329
rect 9232 19292 9260 19323
rect 9858 19292 9864 19304
rect 9232 19264 9864 19292
rect 9858 19252 9864 19264
rect 9916 19252 9922 19304
rect 10152 19301 10180 19332
rect 10226 19320 10232 19372
rect 10284 19360 10290 19372
rect 10796 19369 10824 19400
rect 10321 19363 10379 19369
rect 10321 19360 10333 19363
rect 10284 19332 10333 19360
rect 10284 19320 10290 19332
rect 10321 19329 10333 19332
rect 10367 19329 10379 19363
rect 10321 19323 10379 19329
rect 10781 19363 10839 19369
rect 10781 19329 10793 19363
rect 10827 19329 10839 19363
rect 10781 19323 10839 19329
rect 10873 19363 10931 19369
rect 10873 19329 10885 19363
rect 10919 19329 10931 19363
rect 10873 19323 10931 19329
rect 10137 19295 10195 19301
rect 10137 19261 10149 19295
rect 10183 19261 10195 19295
rect 10137 19255 10195 19261
rect 10686 19252 10692 19304
rect 10744 19292 10750 19304
rect 10888 19292 10916 19323
rect 10744 19264 10916 19292
rect 10744 19252 10750 19264
rect 9401 19227 9459 19233
rect 9401 19193 9413 19227
rect 9447 19224 9459 19227
rect 9447 19196 10088 19224
rect 9447 19193 9459 19196
rect 9401 19187 9459 19193
rect 8757 19159 8815 19165
rect 8757 19156 8769 19159
rect 8352 19128 8769 19156
rect 8352 19116 8358 19128
rect 8757 19125 8769 19128
rect 8803 19125 8815 19159
rect 8757 19119 8815 19125
rect 9030 19116 9036 19168
rect 9088 19156 9094 19168
rect 9493 19159 9551 19165
rect 9493 19156 9505 19159
rect 9088 19128 9505 19156
rect 9088 19116 9094 19128
rect 9493 19125 9505 19128
rect 9539 19125 9551 19159
rect 9493 19119 9551 19125
rect 9769 19159 9827 19165
rect 9769 19125 9781 19159
rect 9815 19156 9827 19159
rect 9858 19156 9864 19168
rect 9815 19128 9864 19156
rect 9815 19125 9827 19128
rect 9769 19119 9827 19125
rect 9858 19116 9864 19128
rect 9916 19116 9922 19168
rect 10060 19165 10088 19196
rect 10045 19159 10103 19165
rect 10045 19125 10057 19159
rect 10091 19125 10103 19159
rect 10980 19156 11008 19400
rect 11072 19400 12940 19428
rect 13004 19400 13185 19428
rect 11072 19369 11100 19400
rect 11057 19363 11115 19369
rect 11057 19329 11069 19363
rect 11103 19329 11115 19363
rect 11057 19323 11115 19329
rect 11149 19363 11207 19369
rect 11149 19329 11161 19363
rect 11195 19360 11207 19363
rect 11238 19360 11244 19372
rect 11195 19332 11244 19360
rect 11195 19329 11207 19332
rect 11149 19323 11207 19329
rect 11238 19320 11244 19332
rect 11296 19360 11302 19372
rect 11517 19363 11575 19369
rect 11517 19360 11529 19363
rect 11296 19332 11529 19360
rect 11296 19320 11302 19332
rect 11517 19329 11529 19332
rect 11563 19329 11575 19363
rect 11517 19323 11575 19329
rect 12434 19320 12440 19372
rect 12492 19320 12498 19372
rect 12529 19363 12587 19369
rect 12529 19329 12541 19363
rect 12575 19360 12587 19363
rect 12894 19360 12900 19372
rect 12575 19332 12900 19360
rect 12575 19329 12587 19332
rect 12529 19323 12587 19329
rect 12894 19320 12900 19332
rect 12952 19360 12958 19372
rect 13004 19360 13032 19400
rect 13173 19397 13185 19400
rect 13219 19397 13231 19431
rect 13173 19391 13231 19397
rect 13265 19431 13323 19437
rect 13265 19397 13277 19431
rect 13311 19428 13323 19431
rect 13722 19428 13728 19440
rect 13311 19400 13728 19428
rect 13311 19397 13323 19400
rect 13265 19391 13323 19397
rect 13722 19388 13728 19400
rect 13780 19388 13786 19440
rect 13906 19388 13912 19440
rect 13964 19428 13970 19440
rect 14734 19428 14740 19440
rect 13964 19400 14740 19428
rect 13964 19388 13970 19400
rect 14734 19388 14740 19400
rect 14792 19388 14798 19440
rect 14826 19388 14832 19440
rect 14884 19388 14890 19440
rect 15028 19428 15056 19468
rect 15105 19465 15117 19499
rect 15151 19496 15163 19499
rect 16666 19496 16672 19508
rect 15151 19468 16672 19496
rect 15151 19465 15163 19468
rect 15105 19459 15163 19465
rect 16666 19456 16672 19468
rect 16724 19456 16730 19508
rect 17497 19499 17555 19505
rect 17497 19496 17509 19499
rect 16960 19468 17509 19496
rect 15930 19428 15936 19440
rect 15028 19400 15936 19428
rect 15930 19388 15936 19400
rect 15988 19388 15994 19440
rect 16960 19437 16988 19468
rect 17497 19465 17509 19468
rect 17543 19496 17555 19499
rect 17586 19496 17592 19508
rect 17543 19468 17592 19496
rect 17543 19465 17555 19468
rect 17497 19459 17555 19465
rect 17586 19456 17592 19468
rect 17644 19456 17650 19508
rect 20530 19456 20536 19508
rect 20588 19496 20594 19508
rect 20809 19499 20867 19505
rect 20809 19496 20821 19499
rect 20588 19468 20821 19496
rect 20588 19456 20594 19468
rect 20809 19465 20821 19468
rect 20855 19465 20867 19499
rect 20809 19459 20867 19465
rect 21266 19456 21272 19508
rect 21324 19456 21330 19508
rect 21358 19456 21364 19508
rect 21416 19496 21422 19508
rect 21910 19496 21916 19508
rect 21416 19468 21916 19496
rect 21416 19456 21422 19468
rect 21910 19456 21916 19468
rect 21968 19456 21974 19508
rect 22738 19456 22744 19508
rect 22796 19496 22802 19508
rect 23201 19499 23259 19505
rect 23201 19496 23213 19499
rect 22796 19468 23213 19496
rect 22796 19456 22802 19468
rect 23201 19465 23213 19468
rect 23247 19465 23259 19499
rect 23201 19459 23259 19465
rect 24029 19499 24087 19505
rect 24029 19465 24041 19499
rect 24075 19496 24087 19499
rect 24118 19496 24124 19508
rect 24075 19468 24124 19496
rect 24075 19465 24087 19468
rect 24029 19459 24087 19465
rect 16945 19431 17003 19437
rect 16316 19400 16804 19428
rect 16316 19372 16344 19400
rect 12952 19332 13032 19360
rect 13081 19363 13139 19369
rect 12952 19320 12958 19332
rect 13081 19329 13093 19363
rect 13127 19329 13139 19363
rect 13081 19323 13139 19329
rect 12710 19252 12716 19304
rect 12768 19252 12774 19304
rect 12986 19184 12992 19236
rect 13044 19224 13050 19236
rect 13096 19224 13124 19323
rect 13446 19320 13452 19372
rect 13504 19320 13510 19372
rect 14001 19363 14059 19369
rect 14001 19329 14013 19363
rect 14047 19360 14059 19363
rect 14458 19360 14464 19372
rect 14047 19332 14464 19360
rect 14047 19329 14059 19332
rect 14001 19323 14059 19329
rect 14458 19320 14464 19332
rect 14516 19360 14522 19372
rect 14553 19363 14611 19369
rect 14553 19360 14565 19363
rect 14516 19332 14565 19360
rect 14516 19320 14522 19332
rect 14553 19329 14565 19332
rect 14599 19329 14611 19363
rect 14553 19323 14611 19329
rect 14642 19320 14648 19372
rect 14700 19360 14706 19372
rect 14921 19363 14979 19369
rect 14921 19360 14933 19363
rect 14700 19332 14933 19360
rect 14700 19320 14706 19332
rect 14921 19329 14933 19332
rect 14967 19360 14979 19363
rect 15102 19360 15108 19372
rect 14967 19332 15108 19360
rect 14967 19329 14979 19332
rect 14921 19323 14979 19329
rect 15102 19320 15108 19332
rect 15160 19320 15166 19372
rect 15841 19363 15899 19369
rect 15841 19329 15853 19363
rect 15887 19360 15899 19363
rect 16298 19360 16304 19372
rect 15887 19332 16304 19360
rect 15887 19329 15899 19332
rect 15841 19323 15899 19329
rect 16298 19320 16304 19332
rect 16356 19320 16362 19372
rect 16666 19320 16672 19372
rect 16724 19320 16730 19372
rect 16776 19369 16804 19400
rect 16945 19397 16957 19431
rect 16991 19397 17003 19431
rect 16945 19391 17003 19397
rect 17034 19388 17040 19440
rect 17092 19388 17098 19440
rect 18690 19388 18696 19440
rect 18748 19428 18754 19440
rect 20070 19428 20076 19440
rect 18748 19400 20076 19428
rect 18748 19388 18754 19400
rect 20070 19388 20076 19400
rect 20128 19428 20134 19440
rect 20257 19431 20315 19437
rect 20257 19428 20269 19431
rect 20128 19400 20269 19428
rect 20128 19388 20134 19400
rect 20257 19397 20269 19400
rect 20303 19428 20315 19431
rect 20303 19400 20576 19428
rect 20303 19397 20315 19400
rect 20257 19391 20315 19397
rect 16762 19363 16820 19369
rect 16762 19329 16774 19363
rect 16808 19329 16820 19363
rect 16762 19323 16820 19329
rect 17175 19363 17233 19369
rect 17175 19329 17187 19363
rect 17221 19360 17233 19363
rect 17494 19360 17500 19372
rect 17221 19332 17500 19360
rect 17221 19329 17233 19332
rect 17175 19323 17233 19329
rect 17494 19320 17500 19332
rect 17552 19320 17558 19372
rect 18138 19320 18144 19372
rect 18196 19320 18202 19372
rect 19518 19320 19524 19372
rect 19576 19360 19582 19372
rect 20349 19363 20407 19369
rect 20349 19360 20361 19363
rect 19576 19332 20361 19360
rect 19576 19320 19582 19332
rect 20349 19329 20361 19332
rect 20395 19329 20407 19363
rect 20548 19360 20576 19400
rect 20622 19388 20628 19440
rect 20680 19428 20686 19440
rect 22088 19431 22146 19437
rect 20680 19400 21763 19428
rect 20680 19388 20686 19400
rect 21177 19363 21235 19369
rect 21177 19360 21189 19363
rect 20548 19332 21189 19360
rect 20349 19323 20407 19329
rect 21177 19329 21189 19332
rect 21223 19360 21235 19363
rect 21358 19360 21364 19372
rect 21223 19332 21364 19360
rect 21223 19329 21235 19332
rect 21177 19323 21235 19329
rect 21358 19320 21364 19332
rect 21416 19320 21422 19372
rect 21735 19334 21763 19400
rect 22088 19397 22100 19431
rect 22134 19428 22146 19431
rect 22370 19428 22376 19440
rect 22134 19400 22376 19428
rect 22134 19397 22146 19400
rect 22088 19391 22146 19397
rect 22370 19388 22376 19400
rect 22428 19388 22434 19440
rect 23216 19360 23244 19459
rect 24118 19456 24124 19468
rect 24176 19456 24182 19508
rect 24397 19499 24455 19505
rect 24397 19465 24409 19499
rect 24443 19496 24455 19499
rect 24854 19496 24860 19508
rect 24443 19468 24860 19496
rect 24443 19465 24455 19468
rect 24397 19459 24455 19465
rect 23658 19388 23664 19440
rect 23716 19388 23722 19440
rect 23477 19363 23535 19369
rect 23477 19360 23489 19363
rect 21735 19306 21772 19334
rect 23216 19332 23489 19360
rect 23477 19329 23489 19332
rect 23523 19329 23535 19363
rect 23477 19323 23535 19329
rect 23750 19320 23756 19372
rect 23808 19320 23814 19372
rect 23845 19363 23903 19369
rect 23845 19329 23857 19363
rect 23891 19360 23903 19363
rect 24412 19360 24440 19459
rect 24854 19456 24860 19468
rect 24912 19456 24918 19508
rect 25041 19499 25099 19505
rect 25041 19465 25053 19499
rect 25087 19496 25099 19499
rect 25961 19499 26019 19505
rect 25961 19496 25973 19499
rect 25087 19468 25973 19496
rect 25087 19465 25099 19468
rect 25041 19459 25099 19465
rect 25961 19465 25973 19468
rect 26007 19496 26019 19499
rect 26234 19496 26240 19508
rect 26007 19468 26240 19496
rect 26007 19465 26019 19468
rect 25961 19459 26019 19465
rect 26234 19456 26240 19468
rect 26292 19456 26298 19508
rect 26329 19499 26387 19505
rect 26329 19465 26341 19499
rect 26375 19496 26387 19499
rect 28074 19496 28080 19508
rect 26375 19468 28080 19496
rect 26375 19465 26387 19468
rect 26329 19459 26387 19465
rect 28074 19456 28080 19468
rect 28132 19456 28138 19508
rect 28718 19456 28724 19508
rect 28776 19496 28782 19508
rect 29086 19496 29092 19508
rect 28776 19468 29092 19496
rect 28776 19456 28782 19468
rect 29086 19456 29092 19468
rect 29144 19456 29150 19508
rect 29365 19499 29423 19505
rect 29365 19465 29377 19499
rect 29411 19496 29423 19499
rect 29914 19496 29920 19508
rect 29411 19468 29920 19496
rect 29411 19465 29423 19468
rect 29365 19459 29423 19465
rect 29914 19456 29920 19468
rect 29972 19456 29978 19508
rect 31202 19456 31208 19508
rect 31260 19496 31266 19508
rect 32309 19499 32367 19505
rect 32309 19496 32321 19499
rect 31260 19468 32321 19496
rect 31260 19456 31266 19468
rect 32309 19465 32321 19468
rect 32355 19465 32367 19499
rect 32309 19459 32367 19465
rect 25501 19431 25559 19437
rect 25501 19397 25513 19431
rect 25547 19397 25559 19431
rect 25501 19391 25559 19397
rect 26053 19431 26111 19437
rect 26053 19397 26065 19431
rect 26099 19428 26111 19431
rect 26418 19428 26424 19440
rect 26099 19400 26424 19428
rect 26099 19397 26111 19400
rect 26053 19391 26111 19397
rect 23891 19332 24440 19360
rect 24949 19363 25007 19369
rect 23891 19329 23903 19332
rect 23845 19323 23903 19329
rect 24949 19329 24961 19363
rect 24995 19360 25007 19363
rect 24995 19332 25360 19360
rect 24995 19329 25007 19332
rect 24949 19323 25007 19329
rect 13630 19252 13636 19304
rect 13688 19252 13694 19304
rect 14277 19295 14335 19301
rect 14277 19261 14289 19295
rect 14323 19292 14335 19295
rect 14366 19292 14372 19304
rect 14323 19264 14372 19292
rect 14323 19261 14335 19264
rect 14277 19255 14335 19261
rect 14366 19252 14372 19264
rect 14424 19252 14430 19304
rect 14734 19252 14740 19304
rect 14792 19292 14798 19304
rect 15289 19295 15347 19301
rect 15289 19292 15301 19295
rect 14792 19264 15301 19292
rect 14792 19252 14798 19264
rect 15289 19261 15301 19264
rect 15335 19261 15347 19295
rect 15289 19255 15347 19261
rect 16022 19252 16028 19304
rect 16080 19252 16086 19304
rect 16206 19252 16212 19304
rect 16264 19292 16270 19304
rect 20165 19295 20223 19301
rect 20165 19292 20177 19295
rect 16264 19264 20177 19292
rect 16264 19252 16270 19264
rect 20165 19261 20177 19264
rect 20211 19292 20223 19295
rect 20438 19292 20444 19304
rect 20211 19264 20444 19292
rect 20211 19261 20223 19264
rect 20165 19255 20223 19261
rect 20438 19252 20444 19264
rect 20496 19252 20502 19304
rect 21453 19295 21511 19301
rect 21453 19261 21465 19295
rect 21499 19292 21511 19295
rect 21634 19292 21640 19304
rect 21499 19264 21640 19292
rect 21499 19261 21511 19264
rect 21453 19255 21511 19261
rect 21634 19252 21640 19264
rect 21692 19252 21698 19304
rect 21744 19292 21772 19306
rect 21821 19295 21879 19301
rect 21821 19292 21833 19295
rect 21744 19264 21833 19292
rect 21821 19261 21833 19264
rect 21867 19261 21879 19295
rect 21821 19255 21879 19261
rect 13044 19196 13124 19224
rect 13648 19224 13676 19252
rect 13648 19196 19334 19224
rect 13044 19184 13050 19196
rect 11054 19156 11060 19168
rect 10980 19128 11060 19156
rect 10045 19119 10103 19125
rect 11054 19116 11060 19128
rect 11112 19156 11118 19168
rect 11241 19159 11299 19165
rect 11241 19156 11253 19159
rect 11112 19128 11253 19156
rect 11112 19116 11118 19128
rect 11241 19125 11253 19128
rect 11287 19125 11299 19159
rect 11241 19119 11299 19125
rect 12066 19116 12072 19168
rect 12124 19116 12130 19168
rect 13354 19116 13360 19168
rect 13412 19156 13418 19168
rect 13633 19159 13691 19165
rect 13633 19156 13645 19159
rect 13412 19128 13645 19156
rect 13412 19116 13418 19128
rect 13633 19125 13645 19128
rect 13679 19125 13691 19159
rect 13633 19119 13691 19125
rect 15470 19116 15476 19168
rect 15528 19116 15534 19168
rect 16022 19116 16028 19168
rect 16080 19156 16086 19168
rect 16301 19159 16359 19165
rect 16301 19156 16313 19159
rect 16080 19128 16313 19156
rect 16080 19116 16086 19128
rect 16301 19125 16313 19128
rect 16347 19125 16359 19159
rect 16301 19119 16359 19125
rect 17126 19116 17132 19168
rect 17184 19156 17190 19168
rect 17313 19159 17371 19165
rect 17313 19156 17325 19159
rect 17184 19128 17325 19156
rect 17184 19116 17190 19128
rect 17313 19125 17325 19128
rect 17359 19125 17371 19159
rect 17313 19119 17371 19125
rect 17494 19116 17500 19168
rect 17552 19156 17558 19168
rect 17589 19159 17647 19165
rect 17589 19156 17601 19159
rect 17552 19128 17601 19156
rect 17552 19116 17558 19128
rect 17589 19125 17601 19128
rect 17635 19125 17647 19159
rect 17589 19119 17647 19125
rect 18049 19159 18107 19165
rect 18049 19125 18061 19159
rect 18095 19156 18107 19159
rect 18138 19156 18144 19168
rect 18095 19128 18144 19156
rect 18095 19125 18107 19128
rect 18049 19119 18107 19125
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 19306 19156 19334 19196
rect 19610 19156 19616 19168
rect 19306 19128 19616 19156
rect 19610 19116 19616 19128
rect 19668 19116 19674 19168
rect 20530 19116 20536 19168
rect 20588 19156 20594 19168
rect 20717 19159 20775 19165
rect 20717 19156 20729 19159
rect 20588 19128 20729 19156
rect 20588 19116 20594 19128
rect 20717 19125 20729 19128
rect 20763 19125 20775 19159
rect 21836 19156 21864 19255
rect 23106 19252 23112 19304
rect 23164 19292 23170 19304
rect 23860 19292 23888 19323
rect 23164 19264 23888 19292
rect 25332 19292 25360 19332
rect 25406 19320 25412 19372
rect 25464 19360 25470 19372
rect 25516 19360 25544 19391
rect 25685 19363 25743 19369
rect 25685 19360 25697 19363
rect 25464 19332 25697 19360
rect 25464 19320 25470 19332
rect 25685 19329 25697 19332
rect 25731 19329 25743 19363
rect 26068 19360 26096 19391
rect 26418 19388 26424 19400
rect 26476 19388 26482 19440
rect 28258 19388 28264 19440
rect 28316 19428 28322 19440
rect 28997 19431 29055 19437
rect 28316 19400 28396 19428
rect 28316 19388 28322 19400
rect 25685 19323 25743 19329
rect 25792 19332 26096 19360
rect 26170 19363 26228 19369
rect 26579 19364 26637 19369
rect 25792 19292 25820 19332
rect 26170 19329 26182 19363
rect 26216 19360 26228 19363
rect 26528 19363 26648 19364
rect 26528 19360 26591 19363
rect 26216 19332 26591 19360
rect 26625 19346 26648 19363
rect 26216 19329 26228 19332
rect 26170 19323 26228 19329
rect 26579 19329 26591 19332
rect 26579 19323 26608 19329
rect 25332 19264 25820 19292
rect 23164 19252 23170 19264
rect 25958 19252 25964 19304
rect 26016 19292 26022 19304
rect 26602 19294 26608 19323
rect 26660 19294 26666 19346
rect 26786 19320 26792 19372
rect 26844 19360 26850 19372
rect 28368 19369 28396 19400
rect 28997 19397 29009 19431
rect 29043 19428 29055 19431
rect 29178 19428 29184 19440
rect 29043 19400 29184 19428
rect 29043 19397 29055 19400
rect 28997 19391 29055 19397
rect 29178 19388 29184 19400
rect 29236 19428 29242 19440
rect 29236 19400 30052 19428
rect 29236 19388 29242 19400
rect 27525 19363 27583 19369
rect 27525 19360 27537 19363
rect 26844 19332 27537 19360
rect 26844 19320 26850 19332
rect 27525 19329 27537 19332
rect 27571 19360 27583 19363
rect 28353 19363 28411 19369
rect 27571 19332 28304 19360
rect 27571 19329 27583 19332
rect 27525 19323 27583 19329
rect 26016 19264 26556 19292
rect 26016 19252 26022 19264
rect 24026 19184 24032 19236
rect 24084 19224 24090 19236
rect 24213 19227 24271 19233
rect 24213 19224 24225 19227
rect 24084 19196 24225 19224
rect 24084 19184 24090 19196
rect 24213 19193 24225 19196
rect 24259 19224 24271 19227
rect 24259 19196 25176 19224
rect 24259 19193 24271 19196
rect 24213 19187 24271 19193
rect 22186 19156 22192 19168
rect 21836 19128 22192 19156
rect 20717 19119 20775 19125
rect 22186 19116 22192 19128
rect 22244 19116 22250 19168
rect 24394 19116 24400 19168
rect 24452 19156 24458 19168
rect 24765 19159 24823 19165
rect 24765 19156 24777 19159
rect 24452 19128 24777 19156
rect 24452 19116 24458 19128
rect 24765 19125 24777 19128
rect 24811 19125 24823 19159
rect 25148 19156 25176 19196
rect 25222 19184 25228 19236
rect 25280 19224 25286 19236
rect 25501 19227 25559 19233
rect 25501 19224 25513 19227
rect 25280 19196 25513 19224
rect 25280 19184 25286 19196
rect 25501 19193 25513 19196
rect 25547 19224 25559 19227
rect 26528 19224 26556 19264
rect 27798 19224 27804 19236
rect 25547 19196 26464 19224
rect 26528 19196 27804 19224
rect 25547 19193 25559 19196
rect 25501 19187 25559 19193
rect 26436 19168 26464 19196
rect 27798 19184 27804 19196
rect 27856 19184 27862 19236
rect 25682 19156 25688 19168
rect 25148 19128 25688 19156
rect 24765 19119 24823 19125
rect 25682 19116 25688 19128
rect 25740 19116 25746 19168
rect 25866 19116 25872 19168
rect 25924 19156 25930 19168
rect 26326 19156 26332 19168
rect 25924 19128 26332 19156
rect 25924 19116 25930 19128
rect 26326 19116 26332 19128
rect 26384 19116 26390 19168
rect 26418 19116 26424 19168
rect 26476 19116 26482 19168
rect 27338 19116 27344 19168
rect 27396 19116 27402 19168
rect 27890 19116 27896 19168
rect 27948 19156 27954 19168
rect 28169 19159 28227 19165
rect 28169 19156 28181 19159
rect 27948 19128 28181 19156
rect 27948 19116 27954 19128
rect 28169 19125 28181 19128
rect 28215 19125 28227 19159
rect 28276 19156 28304 19332
rect 28353 19329 28365 19363
rect 28399 19329 28411 19363
rect 28353 19323 28411 19329
rect 28644 19332 29224 19360
rect 28534 19252 28540 19304
rect 28592 19292 28598 19304
rect 28644 19292 28672 19332
rect 28592 19264 28672 19292
rect 28721 19295 28779 19301
rect 28592 19252 28598 19264
rect 28721 19261 28733 19295
rect 28767 19292 28779 19295
rect 28994 19292 29000 19304
rect 28767 19264 29000 19292
rect 28767 19261 28779 19264
rect 28721 19255 28779 19261
rect 28994 19252 29000 19264
rect 29052 19252 29058 19304
rect 29196 19301 29224 19332
rect 29638 19320 29644 19372
rect 29696 19320 29702 19372
rect 30024 19369 30052 19400
rect 30009 19363 30067 19369
rect 30009 19329 30021 19363
rect 30055 19360 30067 19363
rect 30745 19363 30803 19369
rect 30745 19360 30757 19363
rect 30055 19332 30757 19360
rect 30055 19329 30067 19332
rect 30009 19323 30067 19329
rect 30745 19329 30757 19332
rect 30791 19329 30803 19363
rect 30745 19323 30803 19329
rect 32122 19320 32128 19372
rect 32180 19320 32186 19372
rect 32324 19360 32352 19459
rect 32401 19363 32459 19369
rect 32401 19360 32413 19363
rect 32324 19332 32413 19360
rect 32401 19329 32413 19332
rect 32447 19329 32459 19363
rect 32401 19323 32459 19329
rect 29196 19295 29264 19301
rect 29196 19264 29218 19295
rect 29206 19261 29218 19264
rect 29252 19292 29264 19295
rect 29822 19292 29828 19304
rect 29252 19264 29828 19292
rect 29252 19261 29264 19264
rect 29206 19255 29264 19261
rect 29822 19252 29828 19264
rect 29880 19252 29886 19304
rect 30101 19295 30159 19301
rect 30101 19261 30113 19295
rect 30147 19261 30159 19295
rect 30101 19255 30159 19261
rect 29086 19184 29092 19236
rect 29144 19224 29150 19236
rect 29457 19227 29515 19233
rect 29457 19224 29469 19227
rect 29144 19196 29469 19224
rect 29144 19184 29150 19196
rect 29457 19193 29469 19196
rect 29503 19193 29515 19227
rect 30116 19224 30144 19255
rect 30466 19252 30472 19304
rect 30524 19252 30530 19304
rect 32858 19252 32864 19304
rect 32916 19292 32922 19304
rect 34517 19295 34575 19301
rect 34517 19292 34529 19295
rect 32916 19264 34529 19292
rect 32916 19252 32922 19264
rect 34517 19261 34529 19264
rect 34563 19292 34575 19295
rect 34882 19292 34888 19304
rect 34563 19264 34888 19292
rect 34563 19261 34575 19264
rect 34517 19255 34575 19261
rect 34882 19252 34888 19264
rect 34940 19252 34946 19304
rect 30558 19224 30564 19236
rect 30116 19196 30564 19224
rect 29457 19187 29515 19193
rect 30558 19184 30564 19196
rect 30616 19184 30622 19236
rect 29362 19156 29368 19168
rect 28276 19128 29368 19156
rect 28169 19119 28227 19125
rect 29362 19116 29368 19128
rect 29420 19116 29426 19168
rect 30377 19159 30435 19165
rect 30377 19125 30389 19159
rect 30423 19156 30435 19159
rect 31018 19156 31024 19168
rect 30423 19128 31024 19156
rect 30423 19125 30435 19128
rect 30377 19119 30435 19125
rect 31018 19116 31024 19128
rect 31076 19116 31082 19168
rect 32585 19159 32643 19165
rect 32585 19125 32597 19159
rect 32631 19156 32643 19159
rect 32766 19156 32772 19168
rect 32631 19128 32772 19156
rect 32631 19125 32643 19128
rect 32585 19119 32643 19125
rect 32766 19116 32772 19128
rect 32824 19116 32830 19168
rect 1104 19066 35328 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 35328 19066
rect 1104 18992 35328 19014
rect 5442 18912 5448 18964
rect 5500 18952 5506 18964
rect 5500 18924 6592 18952
rect 5500 18912 5506 18924
rect 6564 18884 6592 18924
rect 7006 18912 7012 18964
rect 7064 18912 7070 18964
rect 7926 18912 7932 18964
rect 7984 18912 7990 18964
rect 9600 18924 12848 18952
rect 6564 18856 9444 18884
rect 7576 18825 7604 18856
rect 9416 18828 9444 18856
rect 9600 18828 9628 18924
rect 12820 18884 12848 18924
rect 12894 18912 12900 18964
rect 12952 18912 12958 18964
rect 14274 18912 14280 18964
rect 14332 18912 14338 18964
rect 14366 18912 14372 18964
rect 14424 18952 14430 18964
rect 14461 18955 14519 18961
rect 14461 18952 14473 18955
rect 14424 18924 14473 18952
rect 14424 18912 14430 18924
rect 14461 18921 14473 18924
rect 14507 18921 14519 18955
rect 16206 18952 16212 18964
rect 14461 18915 14519 18921
rect 14936 18924 16212 18952
rect 14936 18884 14964 18924
rect 16206 18912 16212 18924
rect 16264 18912 16270 18964
rect 16298 18912 16304 18964
rect 16356 18912 16362 18964
rect 18230 18912 18236 18964
rect 18288 18912 18294 18964
rect 19245 18955 19303 18961
rect 19245 18921 19257 18955
rect 19291 18952 19303 18955
rect 19518 18952 19524 18964
rect 19291 18924 19524 18952
rect 19291 18921 19303 18924
rect 19245 18915 19303 18921
rect 19518 18912 19524 18924
rect 19576 18912 19582 18964
rect 20438 18912 20444 18964
rect 20496 18952 20502 18964
rect 20993 18955 21051 18961
rect 20993 18952 21005 18955
rect 20496 18924 21005 18952
rect 20496 18912 20502 18924
rect 20993 18921 21005 18924
rect 21039 18952 21051 18955
rect 21361 18955 21419 18961
rect 21361 18952 21373 18955
rect 21039 18924 21373 18952
rect 21039 18921 21051 18924
rect 20993 18915 21051 18921
rect 21361 18921 21373 18924
rect 21407 18952 21419 18955
rect 21818 18952 21824 18964
rect 21407 18924 21824 18952
rect 21407 18921 21419 18924
rect 21361 18915 21419 18921
rect 21818 18912 21824 18924
rect 21876 18912 21882 18964
rect 21910 18912 21916 18964
rect 21968 18952 21974 18964
rect 23658 18952 23664 18964
rect 21968 18924 23664 18952
rect 21968 18912 21974 18924
rect 23658 18912 23664 18924
rect 23716 18912 23722 18964
rect 23750 18912 23756 18964
rect 23808 18952 23814 18964
rect 24029 18955 24087 18961
rect 24029 18952 24041 18955
rect 23808 18924 24041 18952
rect 23808 18912 23814 18924
rect 24029 18921 24041 18924
rect 24075 18921 24087 18955
rect 24029 18915 24087 18921
rect 25406 18912 25412 18964
rect 25464 18912 25470 18964
rect 26234 18912 26240 18964
rect 26292 18912 26298 18964
rect 26326 18912 26332 18964
rect 26384 18952 26390 18964
rect 27338 18952 27344 18964
rect 26384 18924 27344 18952
rect 26384 18912 26390 18924
rect 27338 18912 27344 18924
rect 27396 18912 27402 18964
rect 27430 18912 27436 18964
rect 27488 18912 27494 18964
rect 28994 18912 29000 18964
rect 29052 18952 29058 18964
rect 30190 18952 30196 18964
rect 29052 18924 30196 18952
rect 29052 18912 29058 18924
rect 30190 18912 30196 18924
rect 30248 18952 30254 18964
rect 30248 18924 30512 18952
rect 30248 18912 30254 18924
rect 12820 18856 14964 18884
rect 16022 18844 16028 18896
rect 16080 18884 16086 18896
rect 19334 18884 19340 18896
rect 16080 18856 19340 18884
rect 16080 18844 16086 18856
rect 19334 18844 19340 18856
rect 19392 18844 19398 18896
rect 22373 18887 22431 18893
rect 22373 18853 22385 18887
rect 22419 18884 22431 18887
rect 22646 18884 22652 18896
rect 22419 18856 22652 18884
rect 22419 18853 22431 18856
rect 22373 18847 22431 18853
rect 22646 18844 22652 18856
rect 22704 18844 22710 18896
rect 23842 18844 23848 18896
rect 23900 18884 23906 18896
rect 26973 18887 27031 18893
rect 26973 18884 26985 18887
rect 23900 18856 26985 18884
rect 23900 18844 23906 18856
rect 26973 18853 26985 18856
rect 27019 18853 27031 18887
rect 26973 18847 27031 18853
rect 27249 18887 27307 18893
rect 27249 18853 27261 18887
rect 27295 18853 27307 18887
rect 29178 18884 29184 18896
rect 27249 18847 27307 18853
rect 28092 18856 29184 18884
rect 7561 18819 7619 18825
rect 7561 18785 7573 18819
rect 7607 18785 7619 18819
rect 7561 18779 7619 18785
rect 7745 18819 7803 18825
rect 7745 18785 7757 18819
rect 7791 18816 7803 18819
rect 7926 18816 7932 18828
rect 7791 18788 7932 18816
rect 7791 18785 7803 18788
rect 7745 18779 7803 18785
rect 7926 18776 7932 18788
rect 7984 18776 7990 18828
rect 8573 18819 8631 18825
rect 8573 18785 8585 18819
rect 8619 18816 8631 18819
rect 9306 18816 9312 18828
rect 8619 18788 9312 18816
rect 8619 18785 8631 18788
rect 8573 18779 8631 18785
rect 9306 18776 9312 18788
rect 9364 18776 9370 18828
rect 9398 18776 9404 18828
rect 9456 18776 9462 18828
rect 9582 18776 9588 18828
rect 9640 18776 9646 18828
rect 14918 18776 14924 18828
rect 14976 18776 14982 18828
rect 17218 18776 17224 18828
rect 17276 18776 17282 18828
rect 17313 18819 17371 18825
rect 17313 18785 17325 18819
rect 17359 18816 17371 18819
rect 17359 18788 18092 18816
rect 17359 18785 17371 18788
rect 17313 18779 17371 18785
rect 1302 18708 1308 18760
rect 1360 18748 1366 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 1360 18720 1409 18748
rect 1360 18708 1366 18720
rect 1397 18717 1409 18720
rect 1443 18748 1455 18751
rect 1857 18751 1915 18757
rect 1857 18748 1869 18751
rect 1443 18720 1869 18748
rect 1443 18717 1455 18720
rect 1397 18711 1455 18717
rect 1857 18717 1869 18720
rect 1903 18717 1915 18751
rect 1857 18711 1915 18717
rect 3510 18708 3516 18760
rect 3568 18748 3574 18760
rect 3789 18751 3847 18757
rect 3789 18748 3801 18751
rect 3568 18720 3801 18748
rect 3568 18708 3574 18720
rect 3789 18717 3801 18720
rect 3835 18748 3847 18751
rect 5629 18751 5687 18757
rect 5629 18748 5641 18751
rect 3835 18720 5641 18748
rect 3835 18717 3847 18720
rect 3789 18711 3847 18717
rect 5629 18717 5641 18720
rect 5675 18717 5687 18751
rect 5629 18711 5687 18717
rect 7006 18708 7012 18760
rect 7064 18748 7070 18760
rect 9769 18751 9827 18757
rect 7064 18720 7236 18748
rect 7064 18708 7070 18720
rect 3878 18640 3884 18692
rect 3936 18680 3942 18692
rect 4034 18683 4092 18689
rect 4034 18680 4046 18683
rect 3936 18652 4046 18680
rect 3936 18640 3942 18652
rect 4034 18649 4046 18652
rect 4080 18649 4092 18683
rect 4034 18643 4092 18649
rect 5896 18683 5954 18689
rect 5896 18649 5908 18683
rect 5942 18680 5954 18683
rect 7208 18680 7236 18720
rect 9769 18717 9781 18751
rect 9815 18748 9827 18751
rect 11517 18751 11575 18757
rect 11517 18748 11529 18751
rect 9815 18720 11529 18748
rect 9815 18717 9827 18720
rect 9769 18711 9827 18717
rect 11517 18717 11529 18720
rect 11563 18717 11575 18751
rect 11517 18711 11575 18717
rect 11784 18751 11842 18757
rect 11784 18717 11796 18751
rect 11830 18748 11842 18751
rect 12066 18748 12072 18760
rect 11830 18720 12072 18748
rect 11830 18717 11842 18720
rect 11784 18711 11842 18717
rect 7469 18683 7527 18689
rect 7469 18680 7481 18683
rect 5942 18652 7144 18680
rect 7208 18652 7481 18680
rect 5942 18649 5954 18652
rect 5896 18643 5954 18649
rect 1581 18615 1639 18621
rect 1581 18581 1593 18615
rect 1627 18612 1639 18615
rect 1762 18612 1768 18624
rect 1627 18584 1768 18612
rect 1627 18581 1639 18584
rect 1581 18575 1639 18581
rect 1762 18572 1768 18584
rect 1820 18572 1826 18624
rect 4154 18572 4160 18624
rect 4212 18612 4218 18624
rect 4890 18612 4896 18624
rect 4212 18584 4896 18612
rect 4212 18572 4218 18584
rect 4890 18572 4896 18584
rect 4948 18612 4954 18624
rect 5169 18615 5227 18621
rect 5169 18612 5181 18615
rect 4948 18584 5181 18612
rect 4948 18572 4954 18584
rect 5169 18581 5181 18584
rect 5215 18581 5227 18615
rect 5169 18575 5227 18581
rect 5350 18572 5356 18624
rect 5408 18572 5414 18624
rect 7116 18621 7144 18652
rect 7469 18649 7481 18652
rect 7515 18649 7527 18683
rect 7469 18643 7527 18649
rect 8294 18640 8300 18692
rect 8352 18640 8358 18692
rect 8389 18683 8447 18689
rect 8389 18649 8401 18683
rect 8435 18680 8447 18683
rect 8435 18652 9076 18680
rect 8435 18649 8447 18652
rect 8389 18643 8447 18649
rect 7101 18615 7159 18621
rect 7101 18581 7113 18615
rect 7147 18581 7159 18615
rect 7101 18575 7159 18581
rect 8938 18572 8944 18624
rect 8996 18572 9002 18624
rect 9048 18612 9076 18652
rect 9122 18640 9128 18692
rect 9180 18680 9186 18692
rect 9309 18683 9367 18689
rect 9309 18680 9321 18683
rect 9180 18652 9321 18680
rect 9180 18640 9186 18652
rect 9309 18649 9321 18652
rect 9355 18649 9367 18683
rect 9309 18643 9367 18649
rect 9398 18640 9404 18692
rect 9456 18680 9462 18692
rect 9784 18680 9812 18711
rect 12066 18708 12072 18720
rect 12124 18708 12130 18760
rect 12342 18708 12348 18760
rect 12400 18748 12406 18760
rect 14093 18751 14151 18757
rect 14093 18748 14105 18751
rect 12400 18720 14105 18748
rect 12400 18708 12406 18720
rect 14093 18717 14105 18720
rect 14139 18717 14151 18751
rect 14093 18711 14151 18717
rect 15188 18751 15246 18757
rect 15188 18717 15200 18751
rect 15234 18748 15246 18751
rect 15470 18748 15476 18760
rect 15234 18720 15476 18748
rect 15234 18717 15246 18720
rect 15188 18711 15246 18717
rect 15470 18708 15476 18720
rect 15528 18708 15534 18760
rect 16945 18751 17003 18757
rect 16945 18717 16957 18751
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 9456 18652 9812 18680
rect 10036 18683 10094 18689
rect 9456 18640 9462 18652
rect 10036 18649 10048 18683
rect 10082 18680 10094 18683
rect 10318 18680 10324 18692
rect 10082 18652 10324 18680
rect 10082 18649 10094 18652
rect 10036 18643 10094 18649
rect 10318 18640 10324 18652
rect 10376 18640 10382 18692
rect 12360 18680 12388 18708
rect 10428 18652 12388 18680
rect 9674 18612 9680 18624
rect 9048 18584 9680 18612
rect 9674 18572 9680 18584
rect 9732 18612 9738 18624
rect 10428 18612 10456 18652
rect 12986 18640 12992 18692
rect 13044 18680 13050 18692
rect 13817 18683 13875 18689
rect 13817 18680 13829 18683
rect 13044 18652 13829 18680
rect 13044 18640 13050 18652
rect 13817 18649 13829 18652
rect 13863 18649 13875 18683
rect 13817 18643 13875 18649
rect 9732 18584 10456 18612
rect 9732 18572 9738 18584
rect 10686 18572 10692 18624
rect 10744 18612 10750 18624
rect 11149 18615 11207 18621
rect 11149 18612 11161 18615
rect 10744 18584 11161 18612
rect 10744 18572 10750 18584
rect 11149 18581 11161 18584
rect 11195 18581 11207 18615
rect 11149 18575 11207 18581
rect 13633 18615 13691 18621
rect 13633 18581 13645 18615
rect 13679 18612 13691 18615
rect 13722 18612 13728 18624
rect 13679 18584 13728 18612
rect 13679 18581 13691 18584
rect 13633 18575 13691 18581
rect 13722 18572 13728 18584
rect 13780 18572 13786 18624
rect 15838 18572 15844 18624
rect 15896 18612 15902 18624
rect 16960 18612 16988 18711
rect 17126 18708 17132 18760
rect 17184 18708 17190 18760
rect 17402 18708 17408 18760
rect 17460 18748 17466 18760
rect 17497 18751 17555 18757
rect 17497 18748 17509 18751
rect 17460 18720 17509 18748
rect 17460 18708 17466 18720
rect 17497 18717 17509 18720
rect 17543 18717 17555 18751
rect 17497 18711 17555 18717
rect 17678 18640 17684 18692
rect 17736 18640 17742 18692
rect 17954 18640 17960 18692
rect 18012 18680 18018 18692
rect 18064 18689 18092 18788
rect 18690 18776 18696 18828
rect 18748 18776 18754 18828
rect 18874 18776 18880 18828
rect 18932 18776 18938 18828
rect 25958 18816 25964 18828
rect 21744 18788 22784 18816
rect 18598 18708 18604 18760
rect 18656 18708 18662 18760
rect 20369 18751 20427 18757
rect 20369 18717 20381 18751
rect 20415 18748 20427 18751
rect 20530 18748 20536 18760
rect 20415 18720 20536 18748
rect 20415 18717 20427 18720
rect 20369 18711 20427 18717
rect 20530 18708 20536 18720
rect 20588 18708 20594 18760
rect 20622 18708 20628 18760
rect 20680 18708 20686 18760
rect 21085 18751 21143 18757
rect 21085 18717 21097 18751
rect 21131 18748 21143 18751
rect 21542 18748 21548 18760
rect 21131 18720 21548 18748
rect 21131 18717 21143 18720
rect 21085 18711 21143 18717
rect 21542 18708 21548 18720
rect 21600 18708 21606 18760
rect 21744 18748 21772 18788
rect 21652 18720 21772 18748
rect 18049 18683 18107 18689
rect 18049 18680 18061 18683
rect 18012 18652 18061 18680
rect 18012 18640 18018 18652
rect 18049 18649 18061 18652
rect 18095 18680 18107 18683
rect 21652 18680 21680 18720
rect 18095 18652 21680 18680
rect 21729 18683 21787 18689
rect 18095 18649 18107 18652
rect 18049 18643 18107 18649
rect 21729 18649 21741 18683
rect 21775 18680 21787 18683
rect 22020 18686 22140 18714
rect 22186 18708 22192 18760
rect 22244 18708 22250 18760
rect 22278 18708 22284 18760
rect 22336 18748 22342 18760
rect 22649 18751 22707 18757
rect 22649 18748 22661 18751
rect 22336 18720 22661 18748
rect 22336 18708 22342 18720
rect 22649 18717 22661 18720
rect 22695 18717 22707 18751
rect 22756 18748 22784 18788
rect 25516 18788 25964 18816
rect 25516 18748 25544 18788
rect 25958 18776 25964 18788
rect 26016 18776 26022 18828
rect 26418 18776 26424 18828
rect 26476 18776 26482 18828
rect 26786 18816 26792 18828
rect 26620 18788 26792 18816
rect 22756 18720 25544 18748
rect 25593 18751 25651 18757
rect 22649 18711 22707 18717
rect 25593 18717 25605 18751
rect 25639 18748 25651 18751
rect 26620 18748 26648 18788
rect 26786 18776 26792 18788
rect 26844 18776 26850 18828
rect 27264 18816 27292 18847
rect 26988 18788 27292 18816
rect 25639 18720 26648 18748
rect 25639 18717 25651 18720
rect 25593 18711 25651 18717
rect 26694 18708 26700 18760
rect 26752 18708 26758 18760
rect 26988 18757 27016 18788
rect 27338 18776 27344 18828
rect 27396 18816 27402 18828
rect 27396 18788 27844 18816
rect 27396 18776 27402 18788
rect 26881 18751 26939 18757
rect 26881 18717 26893 18751
rect 26927 18748 26939 18751
rect 26973 18751 27031 18757
rect 26973 18748 26985 18751
rect 26927 18720 26985 18748
rect 26927 18717 26939 18720
rect 26881 18711 26939 18717
rect 26973 18717 26985 18720
rect 27019 18717 27031 18751
rect 26973 18711 27031 18717
rect 27157 18751 27215 18757
rect 27157 18717 27169 18751
rect 27203 18717 27215 18751
rect 27157 18711 27215 18717
rect 22020 18680 22048 18686
rect 21775 18652 22048 18680
rect 21775 18649 21787 18652
rect 21729 18643 21787 18649
rect 17773 18615 17831 18621
rect 17773 18612 17785 18615
rect 15896 18584 17785 18612
rect 15896 18572 15902 18584
rect 17773 18581 17785 18584
rect 17819 18581 17831 18615
rect 17773 18575 17831 18581
rect 21542 18572 21548 18624
rect 21600 18572 21606 18624
rect 21634 18572 21640 18624
rect 21692 18612 21698 18624
rect 21744 18612 21772 18643
rect 21692 18584 21772 18612
rect 22112 18612 22140 18686
rect 22916 18683 22974 18689
rect 22916 18649 22928 18683
rect 22962 18680 22974 18683
rect 23290 18680 23296 18692
rect 22962 18652 23296 18680
rect 22962 18649 22974 18652
rect 22916 18643 22974 18649
rect 23290 18640 23296 18652
rect 23348 18640 23354 18692
rect 26050 18640 26056 18692
rect 26108 18640 26114 18692
rect 26234 18640 26240 18692
rect 26292 18680 26298 18692
rect 27172 18680 27200 18711
rect 27430 18708 27436 18760
rect 27488 18708 27494 18760
rect 27816 18757 27844 18788
rect 28092 18757 28120 18856
rect 29178 18844 29184 18856
rect 29236 18844 29242 18896
rect 30374 18884 30380 18896
rect 30300 18856 30380 18884
rect 29638 18816 29644 18828
rect 28184 18788 29644 18816
rect 28184 18757 28212 18788
rect 29638 18776 29644 18788
rect 29696 18776 29702 18828
rect 27801 18751 27859 18757
rect 27801 18717 27813 18751
rect 27847 18717 27859 18751
rect 27801 18711 27859 18717
rect 28077 18751 28135 18757
rect 28077 18717 28089 18751
rect 28123 18717 28135 18751
rect 28077 18711 28135 18717
rect 28169 18751 28227 18757
rect 28169 18717 28181 18751
rect 28215 18717 28227 18751
rect 28169 18711 28227 18717
rect 28261 18751 28319 18757
rect 28261 18717 28273 18751
rect 28307 18748 28319 18751
rect 28534 18748 28540 18760
rect 28307 18720 28540 18748
rect 28307 18717 28319 18720
rect 28261 18711 28319 18717
rect 28534 18708 28540 18720
rect 28592 18708 28598 18760
rect 28813 18751 28871 18757
rect 28813 18717 28825 18751
rect 28859 18748 28871 18751
rect 29178 18748 29184 18760
rect 28859 18720 29184 18748
rect 28859 18717 28871 18720
rect 28813 18711 28871 18717
rect 29178 18708 29184 18720
rect 29236 18708 29242 18760
rect 30300 18748 30328 18856
rect 30374 18844 30380 18856
rect 30432 18844 30438 18896
rect 30484 18816 30512 18924
rect 32490 18912 32496 18964
rect 32548 18912 32554 18964
rect 30392 18788 30604 18816
rect 30392 18757 30420 18788
rect 29288 18720 30328 18748
rect 30377 18751 30435 18757
rect 26292 18652 27200 18680
rect 27448 18680 27476 18708
rect 27890 18680 27896 18692
rect 27448 18652 27896 18680
rect 26292 18640 26298 18652
rect 22557 18615 22615 18621
rect 22557 18612 22569 18615
rect 22112 18584 22569 18612
rect 21692 18572 21698 18584
rect 22557 18581 22569 18584
rect 22603 18612 22615 18615
rect 23014 18612 23020 18624
rect 22603 18584 23020 18612
rect 22603 18581 22615 18584
rect 22557 18575 22615 18581
rect 23014 18572 23020 18584
rect 23072 18612 23078 18624
rect 25958 18612 25964 18624
rect 23072 18584 25964 18612
rect 23072 18572 23078 18584
rect 25958 18572 25964 18584
rect 26016 18572 26022 18624
rect 26145 18615 26203 18621
rect 26145 18581 26157 18615
rect 26191 18612 26203 18615
rect 26510 18612 26516 18624
rect 26191 18584 26516 18612
rect 26191 18581 26203 18584
rect 26145 18575 26203 18581
rect 26510 18572 26516 18584
rect 26568 18572 26574 18624
rect 26786 18572 26792 18624
rect 26844 18572 26850 18624
rect 27172 18612 27200 18652
rect 27890 18640 27896 18652
rect 27948 18640 27954 18692
rect 28718 18680 28724 18692
rect 28368 18652 28724 18680
rect 28368 18612 28396 18652
rect 28718 18640 28724 18652
rect 28776 18680 28782 18692
rect 29022 18683 29080 18689
rect 29022 18680 29034 18683
rect 28776 18652 29034 18680
rect 28776 18640 28782 18652
rect 29022 18649 29034 18652
rect 29068 18649 29080 18683
rect 29288 18680 29316 18720
rect 30377 18717 30389 18751
rect 30423 18717 30435 18751
rect 30377 18711 30435 18717
rect 30466 18708 30472 18760
rect 30524 18708 30530 18760
rect 29022 18643 29080 18649
rect 29196 18652 29316 18680
rect 27172 18584 28396 18612
rect 28442 18572 28448 18624
rect 28500 18572 28506 18624
rect 28902 18572 28908 18624
rect 28960 18572 28966 18624
rect 29196 18621 29224 18652
rect 29362 18640 29368 18692
rect 29420 18680 29426 18692
rect 29641 18683 29699 18689
rect 29641 18680 29653 18683
rect 29420 18652 29653 18680
rect 29420 18640 29426 18652
rect 29641 18649 29653 18652
rect 29687 18680 29699 18683
rect 30484 18680 30512 18708
rect 29687 18652 30512 18680
rect 29687 18649 29699 18652
rect 29641 18643 29699 18649
rect 29181 18615 29239 18621
rect 29181 18581 29193 18615
rect 29227 18581 29239 18615
rect 29181 18575 29239 18581
rect 29546 18572 29552 18624
rect 29604 18612 29610 18624
rect 29733 18615 29791 18621
rect 29733 18612 29745 18615
rect 29604 18584 29745 18612
rect 29604 18572 29610 18584
rect 29733 18581 29745 18584
rect 29779 18581 29791 18615
rect 29733 18575 29791 18581
rect 29825 18615 29883 18621
rect 29825 18581 29837 18615
rect 29871 18612 29883 18615
rect 30006 18612 30012 18624
rect 29871 18584 30012 18612
rect 29871 18581 29883 18584
rect 29825 18575 29883 18581
rect 30006 18572 30012 18584
rect 30064 18572 30070 18624
rect 30098 18572 30104 18624
rect 30156 18612 30162 18624
rect 30193 18615 30251 18621
rect 30193 18612 30205 18615
rect 30156 18584 30205 18612
rect 30156 18572 30162 18584
rect 30193 18581 30205 18584
rect 30239 18612 30251 18615
rect 30282 18612 30288 18624
rect 30239 18584 30288 18612
rect 30239 18581 30251 18584
rect 30193 18575 30251 18581
rect 30282 18572 30288 18584
rect 30340 18612 30346 18624
rect 30469 18615 30527 18621
rect 30469 18612 30481 18615
rect 30340 18584 30481 18612
rect 30340 18572 30346 18584
rect 30469 18581 30481 18584
rect 30515 18581 30527 18615
rect 30576 18612 30604 18788
rect 31018 18776 31024 18828
rect 31076 18776 31082 18828
rect 32214 18776 32220 18828
rect 32272 18776 32278 18828
rect 32582 18776 32588 18828
rect 32640 18816 32646 18828
rect 32677 18819 32735 18825
rect 32677 18816 32689 18819
rect 32640 18788 32689 18816
rect 32640 18776 32646 18788
rect 32677 18785 32689 18788
rect 32723 18816 32735 18819
rect 32723 18788 34468 18816
rect 32723 18785 32735 18788
rect 32677 18779 32735 18785
rect 30742 18708 30748 18760
rect 30800 18708 30806 18760
rect 32232 18748 32260 18776
rect 32154 18720 32260 18748
rect 32766 18708 32772 18760
rect 32824 18708 32830 18760
rect 34146 18708 34152 18760
rect 34204 18708 34210 18760
rect 34440 18757 34468 18788
rect 34425 18751 34483 18757
rect 34425 18717 34437 18751
rect 34471 18717 34483 18751
rect 34425 18711 34483 18717
rect 31754 18612 31760 18624
rect 30576 18584 31760 18612
rect 30469 18575 30527 18581
rect 31754 18572 31760 18584
rect 31812 18572 31818 18624
rect 33137 18615 33195 18621
rect 33137 18581 33149 18615
rect 33183 18612 33195 18615
rect 33686 18612 33692 18624
rect 33183 18584 33692 18612
rect 33183 18581 33195 18584
rect 33137 18575 33195 18581
rect 33686 18572 33692 18584
rect 33744 18572 33750 18624
rect 33778 18572 33784 18624
rect 33836 18612 33842 18624
rect 33965 18615 34023 18621
rect 33965 18612 33977 18615
rect 33836 18584 33977 18612
rect 33836 18572 33842 18584
rect 33965 18581 33977 18584
rect 34011 18581 34023 18615
rect 33965 18575 34023 18581
rect 34333 18615 34391 18621
rect 34333 18581 34345 18615
rect 34379 18612 34391 18615
rect 34514 18612 34520 18624
rect 34379 18584 34520 18612
rect 34379 18581 34391 18584
rect 34333 18575 34391 18581
rect 34514 18572 34520 18584
rect 34572 18572 34578 18624
rect 1104 18522 35328 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35328 18522
rect 1104 18448 35328 18470
rect 3789 18411 3847 18417
rect 3789 18377 3801 18411
rect 3835 18408 3847 18411
rect 3878 18408 3884 18420
rect 3835 18380 3884 18408
rect 3835 18377 3847 18380
rect 3789 18371 3847 18377
rect 3878 18368 3884 18380
rect 3936 18368 3942 18420
rect 4154 18368 4160 18420
rect 4212 18368 4218 18420
rect 4249 18411 4307 18417
rect 4249 18377 4261 18411
rect 4295 18408 4307 18411
rect 5442 18408 5448 18420
rect 4295 18380 5448 18408
rect 4295 18377 4307 18380
rect 4249 18371 4307 18377
rect 5442 18368 5448 18380
rect 5500 18368 5506 18420
rect 7098 18368 7104 18420
rect 7156 18408 7162 18420
rect 7156 18380 9076 18408
rect 7156 18368 7162 18380
rect 5994 18300 6000 18352
rect 6052 18340 6058 18352
rect 8012 18343 8070 18349
rect 6052 18312 7880 18340
rect 6052 18300 6058 18312
rect 7374 18232 7380 18284
rect 7432 18272 7438 18284
rect 7745 18275 7803 18281
rect 7745 18272 7757 18275
rect 7432 18244 7757 18272
rect 7432 18232 7438 18244
rect 7745 18241 7757 18244
rect 7791 18241 7803 18275
rect 7852 18272 7880 18312
rect 8012 18309 8024 18343
rect 8058 18340 8070 18343
rect 8938 18340 8944 18352
rect 8058 18312 8944 18340
rect 8058 18309 8070 18312
rect 8012 18303 8070 18309
rect 8938 18300 8944 18312
rect 8996 18300 9002 18352
rect 9048 18340 9076 18380
rect 9122 18368 9128 18420
rect 9180 18368 9186 18420
rect 9582 18368 9588 18420
rect 9640 18408 9646 18420
rect 9769 18411 9827 18417
rect 9769 18408 9781 18411
rect 9640 18380 9781 18408
rect 9640 18368 9646 18380
rect 9769 18377 9781 18380
rect 9815 18377 9827 18411
rect 9769 18371 9827 18377
rect 10318 18368 10324 18420
rect 10376 18368 10382 18420
rect 10686 18368 10692 18420
rect 10744 18368 10750 18420
rect 10778 18368 10784 18420
rect 10836 18368 10842 18420
rect 12710 18368 12716 18420
rect 12768 18408 12774 18420
rect 12768 18380 14136 18408
rect 12768 18368 12774 18380
rect 10410 18340 10416 18352
rect 9048 18312 10416 18340
rect 10410 18300 10416 18312
rect 10468 18340 10474 18352
rect 13354 18349 13360 18352
rect 13348 18340 13360 18349
rect 10468 18312 10916 18340
rect 13315 18312 13360 18340
rect 10468 18300 10474 18312
rect 10318 18272 10324 18284
rect 7852 18244 10324 18272
rect 7745 18235 7803 18241
rect 10318 18232 10324 18244
rect 10376 18232 10382 18284
rect 4433 18207 4491 18213
rect 4433 18173 4445 18207
rect 4479 18204 4491 18207
rect 4706 18204 4712 18216
rect 4479 18176 4712 18204
rect 4479 18173 4491 18176
rect 4433 18167 4491 18173
rect 4706 18164 4712 18176
rect 4764 18204 4770 18216
rect 5258 18204 5264 18216
rect 4764 18176 5264 18204
rect 4764 18164 4770 18176
rect 5258 18164 5264 18176
rect 5316 18164 5322 18216
rect 10888 18213 10916 18312
rect 13348 18303 13360 18312
rect 13354 18300 13360 18303
rect 13412 18300 13418 18352
rect 13998 18300 14004 18352
rect 14056 18300 14062 18352
rect 14108 18340 14136 18380
rect 14458 18368 14464 18420
rect 14516 18368 14522 18420
rect 21542 18368 21548 18420
rect 21600 18408 21606 18420
rect 22005 18411 22063 18417
rect 22005 18408 22017 18411
rect 21600 18380 22017 18408
rect 21600 18368 21606 18380
rect 22005 18377 22017 18380
rect 22051 18377 22063 18411
rect 22005 18371 22063 18377
rect 22186 18368 22192 18420
rect 22244 18408 22250 18420
rect 22462 18408 22468 18420
rect 22244 18380 22468 18408
rect 22244 18368 22250 18380
rect 22462 18368 22468 18380
rect 22520 18368 22526 18420
rect 22646 18368 22652 18420
rect 22704 18368 22710 18420
rect 23198 18368 23204 18420
rect 23256 18368 23262 18420
rect 23290 18368 23296 18420
rect 23348 18368 23354 18420
rect 23658 18368 23664 18420
rect 23716 18368 23722 18420
rect 23750 18368 23756 18420
rect 23808 18368 23814 18420
rect 24765 18411 24823 18417
rect 24765 18377 24777 18411
rect 24811 18408 24823 18411
rect 25406 18408 25412 18420
rect 24811 18380 25412 18408
rect 24811 18377 24823 18380
rect 24765 18371 24823 18377
rect 25406 18368 25412 18380
rect 25464 18368 25470 18420
rect 25682 18368 25688 18420
rect 25740 18408 25746 18420
rect 25740 18380 26188 18408
rect 25740 18368 25746 18380
rect 14108 18312 19334 18340
rect 14016 18272 14044 18300
rect 14553 18275 14611 18281
rect 14553 18272 14565 18275
rect 14016 18244 14565 18272
rect 14553 18241 14565 18244
rect 14599 18272 14611 18275
rect 14599 18244 15240 18272
rect 14599 18241 14611 18244
rect 14553 18235 14611 18241
rect 10873 18207 10931 18213
rect 10873 18173 10885 18207
rect 10919 18204 10931 18207
rect 11149 18207 11207 18213
rect 11149 18204 11161 18207
rect 10919 18176 11161 18204
rect 10919 18173 10931 18176
rect 10873 18167 10931 18173
rect 11149 18173 11161 18176
rect 11195 18204 11207 18207
rect 12066 18204 12072 18216
rect 11195 18176 12072 18204
rect 11195 18173 11207 18176
rect 11149 18167 11207 18173
rect 12066 18164 12072 18176
rect 12124 18164 12130 18216
rect 13078 18164 13084 18216
rect 13136 18164 13142 18216
rect 15102 18204 15108 18216
rect 14936 18176 15108 18204
rect 9858 18096 9864 18148
rect 9916 18136 9922 18148
rect 9916 18108 12434 18136
rect 9916 18096 9922 18108
rect 7653 18071 7711 18077
rect 7653 18037 7665 18071
rect 7699 18068 7711 18071
rect 7926 18068 7932 18080
rect 7699 18040 7932 18068
rect 7699 18037 7711 18040
rect 7653 18031 7711 18037
rect 7926 18028 7932 18040
rect 7984 18028 7990 18080
rect 9306 18028 9312 18080
rect 9364 18068 9370 18080
rect 9582 18068 9588 18080
rect 9364 18040 9588 18068
rect 9364 18028 9370 18040
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 12406 18068 12434 18108
rect 14090 18096 14096 18148
rect 14148 18136 14154 18148
rect 14366 18136 14372 18148
rect 14148 18108 14372 18136
rect 14148 18096 14154 18108
rect 14366 18096 14372 18108
rect 14424 18136 14430 18148
rect 14936 18145 14964 18176
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 14737 18139 14795 18145
rect 14737 18136 14749 18139
rect 14424 18108 14749 18136
rect 14424 18096 14430 18108
rect 14737 18105 14749 18108
rect 14783 18136 14795 18139
rect 14921 18139 14979 18145
rect 14921 18136 14933 18139
rect 14783 18108 14933 18136
rect 14783 18105 14795 18108
rect 14737 18099 14795 18105
rect 14921 18105 14933 18108
rect 14967 18105 14979 18139
rect 14921 18099 14979 18105
rect 13998 18068 14004 18080
rect 12406 18040 14004 18068
rect 13998 18028 14004 18040
rect 14056 18028 14062 18080
rect 15212 18077 15240 18244
rect 16574 18232 16580 18284
rect 16632 18272 16638 18284
rect 16942 18281 16948 18284
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 16632 18244 16681 18272
rect 16632 18232 16638 18244
rect 16669 18241 16681 18244
rect 16715 18241 16727 18275
rect 16669 18235 16727 18241
rect 16936 18235 16948 18281
rect 16942 18232 16948 18235
rect 17000 18232 17006 18284
rect 19306 18272 19334 18312
rect 21726 18300 21732 18352
rect 21784 18340 21790 18352
rect 21913 18343 21971 18349
rect 21913 18340 21925 18343
rect 21784 18312 21925 18340
rect 21784 18300 21790 18312
rect 21913 18309 21925 18312
rect 21959 18309 21971 18343
rect 21913 18303 21971 18309
rect 22922 18300 22928 18352
rect 22980 18340 22986 18352
rect 24581 18343 24639 18349
rect 22980 18312 24256 18340
rect 22980 18300 22986 18312
rect 22572 18272 22784 18276
rect 19306 18248 23888 18272
rect 19306 18244 22600 18248
rect 22756 18244 23888 18248
rect 21542 18164 21548 18216
rect 21600 18164 21606 18216
rect 22738 18164 22744 18216
rect 22796 18164 22802 18216
rect 22925 18207 22983 18213
rect 22925 18173 22937 18207
rect 22971 18204 22983 18207
rect 23014 18204 23020 18216
rect 22971 18176 23020 18204
rect 22971 18173 22983 18176
rect 22925 18167 22983 18173
rect 23014 18164 23020 18176
rect 23072 18164 23078 18216
rect 23860 18213 23888 18244
rect 23845 18207 23903 18213
rect 23845 18173 23857 18207
rect 23891 18204 23903 18207
rect 24121 18207 24179 18213
rect 24121 18204 24133 18207
rect 23891 18176 24133 18204
rect 23891 18173 23903 18176
rect 23845 18167 23903 18173
rect 24121 18173 24133 18176
rect 24167 18173 24179 18207
rect 24228 18204 24256 18312
rect 24581 18309 24593 18343
rect 24627 18340 24639 18343
rect 25130 18340 25136 18352
rect 24627 18312 25136 18340
rect 24627 18309 24639 18312
rect 24581 18303 24639 18309
rect 25130 18300 25136 18312
rect 25188 18340 25194 18352
rect 25777 18343 25835 18349
rect 25777 18340 25789 18343
rect 25188 18312 25789 18340
rect 25188 18300 25194 18312
rect 25777 18309 25789 18312
rect 25823 18340 25835 18343
rect 26050 18340 26056 18352
rect 25823 18312 26056 18340
rect 25823 18309 25835 18312
rect 25777 18303 25835 18309
rect 24673 18275 24731 18281
rect 24673 18241 24685 18275
rect 24719 18272 24731 18275
rect 24854 18272 24860 18284
rect 24719 18244 24860 18272
rect 24719 18241 24731 18244
rect 24673 18235 24731 18241
rect 24854 18232 24860 18244
rect 24912 18232 24918 18284
rect 24949 18275 25007 18281
rect 24949 18241 24961 18275
rect 24995 18272 25007 18275
rect 25222 18272 25228 18284
rect 24995 18244 25228 18272
rect 24995 18241 25007 18244
rect 24949 18235 25007 18241
rect 25222 18232 25228 18244
rect 25280 18232 25286 18284
rect 25976 18281 26004 18312
rect 26050 18300 26056 18312
rect 26108 18300 26114 18352
rect 26160 18340 26188 18380
rect 26326 18368 26332 18420
rect 26384 18368 26390 18420
rect 28905 18411 28963 18417
rect 28905 18377 28917 18411
rect 28951 18408 28963 18411
rect 29086 18408 29092 18420
rect 28951 18380 29092 18408
rect 28951 18377 28963 18380
rect 28905 18371 28963 18377
rect 29086 18368 29092 18380
rect 29144 18368 29150 18420
rect 29181 18411 29239 18417
rect 29181 18377 29193 18411
rect 29227 18408 29239 18411
rect 29638 18408 29644 18420
rect 29227 18380 29644 18408
rect 29227 18377 29239 18380
rect 29181 18371 29239 18377
rect 26446 18343 26504 18349
rect 26160 18312 26372 18340
rect 25961 18275 26019 18281
rect 25961 18241 25973 18275
rect 26007 18241 26019 18275
rect 25961 18235 26019 18241
rect 25041 18207 25099 18213
rect 25041 18204 25053 18207
rect 24228 18176 25053 18204
rect 24121 18167 24179 18173
rect 25041 18173 25053 18176
rect 25087 18173 25099 18207
rect 25041 18167 25099 18173
rect 25314 18164 25320 18216
rect 25372 18204 25378 18216
rect 26237 18207 26295 18213
rect 25372 18176 25912 18204
rect 25372 18164 25378 18176
rect 19610 18096 19616 18148
rect 19668 18136 19674 18148
rect 20073 18139 20131 18145
rect 20073 18136 20085 18139
rect 19668 18108 20085 18136
rect 19668 18096 19674 18108
rect 20073 18105 20085 18108
rect 20119 18136 20131 18139
rect 24762 18136 24768 18148
rect 20119 18108 24768 18136
rect 20119 18105 20131 18108
rect 20073 18099 20131 18105
rect 24762 18096 24768 18108
rect 24820 18096 24826 18148
rect 24854 18096 24860 18148
rect 24912 18136 24918 18148
rect 25332 18136 25360 18164
rect 25884 18148 25912 18176
rect 26237 18173 26249 18207
rect 26283 18173 26295 18207
rect 26344 18204 26372 18312
rect 26446 18309 26458 18343
rect 26492 18340 26504 18343
rect 26602 18340 26608 18352
rect 26492 18312 26608 18340
rect 26492 18309 26504 18312
rect 26446 18303 26504 18309
rect 26602 18300 26608 18312
rect 26660 18340 26666 18352
rect 27062 18340 27068 18352
rect 26660 18312 27068 18340
rect 26660 18300 26666 18312
rect 27062 18300 27068 18312
rect 27120 18340 27126 18352
rect 27430 18340 27436 18352
rect 27120 18312 27436 18340
rect 27120 18300 27126 18312
rect 27430 18300 27436 18312
rect 27488 18300 27494 18352
rect 28721 18343 28779 18349
rect 28721 18309 28733 18343
rect 28767 18340 28779 18343
rect 29196 18340 29224 18371
rect 29638 18368 29644 18380
rect 29696 18368 29702 18420
rect 31481 18411 31539 18417
rect 31481 18408 31493 18411
rect 30208 18380 31493 18408
rect 28767 18312 29224 18340
rect 28767 18309 28779 18312
rect 28721 18303 28779 18309
rect 29546 18300 29552 18352
rect 29604 18340 29610 18352
rect 30208 18340 30236 18380
rect 29604 18312 30236 18340
rect 29604 18300 29610 18312
rect 30926 18300 30932 18352
rect 30984 18340 30990 18352
rect 31173 18343 31231 18349
rect 31173 18340 31185 18343
rect 30984 18312 31185 18340
rect 30984 18300 30990 18312
rect 31173 18309 31185 18312
rect 31219 18309 31231 18343
rect 31173 18303 31231 18309
rect 27614 18232 27620 18284
rect 27672 18272 27678 18284
rect 28902 18272 28908 18284
rect 27672 18244 28908 18272
rect 27672 18232 27678 18244
rect 28902 18232 28908 18244
rect 28960 18232 28966 18284
rect 28997 18265 29055 18271
rect 28997 18231 29009 18265
rect 29043 18231 29055 18265
rect 29086 18232 29092 18284
rect 29144 18272 29150 18284
rect 29273 18275 29331 18281
rect 29273 18272 29285 18275
rect 29144 18244 29285 18272
rect 29144 18232 29150 18244
rect 29273 18241 29285 18244
rect 29319 18272 29331 18275
rect 30006 18272 30012 18284
rect 29319 18244 30012 18272
rect 29319 18241 29331 18244
rect 29273 18235 29331 18241
rect 30006 18232 30012 18244
rect 30064 18272 30070 18284
rect 30377 18275 30435 18281
rect 30377 18272 30389 18275
rect 30064 18244 30389 18272
rect 30064 18232 30070 18244
rect 30377 18241 30389 18244
rect 30423 18241 30435 18275
rect 30377 18235 30435 18241
rect 28997 18225 29055 18231
rect 28534 18204 28540 18216
rect 26344 18176 28540 18204
rect 26237 18167 26295 18173
rect 24912 18108 25360 18136
rect 24912 18096 24918 18108
rect 25406 18096 25412 18148
rect 25464 18136 25470 18148
rect 25777 18139 25835 18145
rect 25777 18136 25789 18139
rect 25464 18108 25789 18136
rect 25464 18096 25470 18108
rect 25777 18105 25789 18108
rect 25823 18105 25835 18139
rect 25777 18099 25835 18105
rect 25866 18096 25872 18148
rect 25924 18136 25930 18148
rect 26252 18136 26280 18167
rect 28534 18164 28540 18176
rect 28592 18164 28598 18216
rect 26694 18136 26700 18148
rect 25924 18108 26700 18136
rect 25924 18096 25930 18108
rect 26694 18096 26700 18108
rect 26752 18136 26758 18148
rect 27433 18139 27491 18145
rect 27433 18136 27445 18139
rect 26752 18108 27445 18136
rect 26752 18096 26758 18108
rect 27433 18105 27445 18108
rect 27479 18105 27491 18139
rect 29012 18136 29040 18225
rect 30098 18164 30104 18216
rect 30156 18164 30162 18216
rect 31312 18204 31340 18380
rect 31481 18377 31493 18380
rect 31527 18377 31539 18411
rect 31481 18371 31539 18377
rect 32122 18368 32128 18420
rect 32180 18408 32186 18420
rect 32217 18411 32275 18417
rect 32217 18408 32229 18411
rect 32180 18380 32229 18408
rect 32180 18368 32186 18380
rect 32217 18377 32229 18380
rect 32263 18377 32275 18411
rect 32766 18408 32772 18420
rect 32217 18371 32275 18377
rect 32324 18380 32772 18408
rect 31389 18343 31447 18349
rect 31389 18309 31401 18343
rect 31435 18340 31447 18343
rect 31754 18340 31760 18352
rect 31435 18312 31760 18340
rect 31435 18309 31447 18312
rect 31389 18303 31447 18309
rect 31754 18300 31760 18312
rect 31812 18340 31818 18352
rect 32324 18340 32352 18380
rect 32766 18368 32772 18380
rect 32824 18368 32830 18420
rect 31812 18312 32352 18340
rect 31812 18300 31818 18312
rect 33134 18300 33140 18352
rect 33192 18300 33198 18352
rect 33686 18300 33692 18352
rect 33744 18300 33750 18352
rect 31662 18232 31668 18284
rect 31720 18232 31726 18284
rect 31941 18275 31999 18281
rect 31941 18241 31953 18275
rect 31987 18241 31999 18275
rect 31941 18235 31999 18241
rect 31956 18204 31984 18235
rect 34514 18232 34520 18284
rect 34572 18232 34578 18284
rect 34790 18232 34796 18284
rect 34848 18232 34854 18284
rect 31312 18176 31984 18204
rect 33965 18207 34023 18213
rect 33965 18173 33977 18207
rect 34011 18173 34023 18207
rect 33965 18167 34023 18173
rect 30558 18136 30564 18148
rect 29012 18108 30564 18136
rect 27433 18099 27491 18105
rect 30558 18096 30564 18108
rect 30616 18136 30622 18148
rect 31021 18139 31079 18145
rect 31021 18136 31033 18139
rect 30616 18108 31033 18136
rect 30616 18096 30622 18108
rect 31021 18105 31033 18108
rect 31067 18136 31079 18139
rect 31570 18136 31576 18148
rect 31067 18108 31576 18136
rect 31067 18105 31079 18108
rect 31021 18099 31079 18105
rect 31570 18096 31576 18108
rect 31628 18096 31634 18148
rect 15197 18071 15255 18077
rect 15197 18037 15209 18071
rect 15243 18068 15255 18071
rect 16298 18068 16304 18080
rect 15243 18040 16304 18068
rect 15243 18037 15255 18040
rect 15197 18031 15255 18037
rect 16298 18028 16304 18040
rect 16356 18028 16362 18080
rect 17310 18028 17316 18080
rect 17368 18068 17374 18080
rect 18049 18071 18107 18077
rect 18049 18068 18061 18071
rect 17368 18040 18061 18068
rect 17368 18028 17374 18040
rect 18049 18037 18061 18040
rect 18095 18037 18107 18071
rect 18049 18031 18107 18037
rect 18874 18028 18880 18080
rect 18932 18068 18938 18080
rect 19153 18071 19211 18077
rect 19153 18068 19165 18071
rect 18932 18040 19165 18068
rect 18932 18028 18938 18040
rect 19153 18037 19165 18040
rect 19199 18068 19211 18071
rect 22094 18068 22100 18080
rect 19199 18040 22100 18068
rect 19199 18037 19211 18040
rect 19153 18031 19211 18037
rect 22094 18028 22100 18040
rect 22152 18028 22158 18080
rect 22186 18028 22192 18080
rect 22244 18068 22250 18080
rect 22281 18071 22339 18077
rect 22281 18068 22293 18071
rect 22244 18040 22293 18068
rect 22244 18028 22250 18040
rect 22281 18037 22293 18040
rect 22327 18037 22339 18071
rect 22281 18031 22339 18037
rect 24397 18071 24455 18077
rect 24397 18037 24409 18071
rect 24443 18068 24455 18071
rect 24578 18068 24584 18080
rect 24443 18040 24584 18068
rect 24443 18037 24455 18040
rect 24397 18031 24455 18037
rect 24578 18028 24584 18040
rect 24636 18028 24642 18080
rect 24670 18028 24676 18080
rect 24728 18068 24734 18080
rect 26605 18071 26663 18077
rect 26605 18068 26617 18071
rect 24728 18040 26617 18068
rect 24728 18028 24734 18040
rect 26605 18037 26617 18040
rect 26651 18037 26663 18071
rect 26605 18031 26663 18037
rect 28718 18028 28724 18080
rect 28776 18028 28782 18080
rect 29270 18028 29276 18080
rect 29328 18068 29334 18080
rect 29457 18071 29515 18077
rect 29457 18068 29469 18071
rect 29328 18040 29469 18068
rect 29328 18028 29334 18040
rect 29457 18037 29469 18040
rect 29503 18068 29515 18071
rect 29638 18068 29644 18080
rect 29503 18040 29644 18068
rect 29503 18037 29515 18040
rect 29457 18031 29515 18037
rect 29638 18028 29644 18040
rect 29696 18028 29702 18080
rect 29822 18028 29828 18080
rect 29880 18068 29886 18080
rect 31205 18071 31263 18077
rect 31205 18068 31217 18071
rect 29880 18040 31217 18068
rect 29880 18028 29886 18040
rect 31205 18037 31217 18040
rect 31251 18068 31263 18071
rect 31294 18068 31300 18080
rect 31251 18040 31300 18068
rect 31251 18037 31263 18040
rect 31205 18031 31263 18037
rect 31294 18028 31300 18040
rect 31352 18068 31358 18080
rect 31757 18071 31815 18077
rect 31757 18068 31769 18071
rect 31352 18040 31769 18068
rect 31352 18028 31358 18040
rect 31757 18037 31769 18040
rect 31803 18037 31815 18071
rect 31757 18031 31815 18037
rect 32674 18028 32680 18080
rect 32732 18068 32738 18080
rect 33980 18068 34008 18167
rect 32732 18040 34008 18068
rect 32732 18028 32738 18040
rect 1104 17978 35328 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 35328 17978
rect 1104 17904 35328 17926
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 16853 17867 16911 17873
rect 1820 17836 16436 17864
rect 1820 17824 1826 17836
rect 7190 17756 7196 17808
rect 7248 17796 7254 17808
rect 11882 17796 11888 17808
rect 7248 17768 11888 17796
rect 7248 17756 7254 17768
rect 11882 17756 11888 17768
rect 11940 17756 11946 17808
rect 15102 17756 15108 17808
rect 15160 17796 15166 17808
rect 15565 17799 15623 17805
rect 15565 17796 15577 17799
rect 15160 17768 15577 17796
rect 15160 17756 15166 17768
rect 15565 17765 15577 17768
rect 15611 17765 15623 17799
rect 16408 17796 16436 17836
rect 16853 17833 16865 17867
rect 16899 17864 16911 17867
rect 16942 17864 16948 17876
rect 16899 17836 16948 17864
rect 16899 17833 16911 17836
rect 16853 17827 16911 17833
rect 16942 17824 16948 17836
rect 17000 17824 17006 17876
rect 17126 17824 17132 17876
rect 17184 17864 17190 17876
rect 17184 17836 22094 17864
rect 17184 17824 17190 17836
rect 18325 17799 18383 17805
rect 18325 17796 18337 17799
rect 16408 17768 18337 17796
rect 15565 17759 15623 17765
rect 18325 17765 18337 17768
rect 18371 17765 18383 17799
rect 18325 17759 18383 17765
rect 10318 17688 10324 17740
rect 10376 17728 10382 17740
rect 10413 17731 10471 17737
rect 10413 17728 10425 17731
rect 10376 17700 10425 17728
rect 10376 17688 10382 17700
rect 10413 17697 10425 17700
rect 10459 17697 10471 17731
rect 10413 17691 10471 17697
rect 16850 17688 16856 17740
rect 16908 17728 16914 17740
rect 17126 17728 17132 17740
rect 16908 17700 17132 17728
rect 16908 17688 16914 17700
rect 17126 17688 17132 17700
rect 17184 17688 17190 17740
rect 17310 17688 17316 17740
rect 17368 17688 17374 17740
rect 17497 17731 17555 17737
rect 17497 17697 17509 17731
rect 17543 17728 17555 17731
rect 17586 17728 17592 17740
rect 17543 17700 17592 17728
rect 17543 17697 17555 17700
rect 17497 17691 17555 17697
rect 17586 17688 17592 17700
rect 17644 17688 17650 17740
rect 7742 17620 7748 17672
rect 7800 17660 7806 17672
rect 10781 17663 10839 17669
rect 10781 17660 10793 17663
rect 7800 17632 10793 17660
rect 7800 17620 7806 17632
rect 10781 17629 10793 17632
rect 10827 17629 10839 17663
rect 10781 17623 10839 17629
rect 10874 17663 10932 17669
rect 10874 17629 10886 17663
rect 10920 17629 10932 17663
rect 10874 17623 10932 17629
rect 11287 17663 11345 17669
rect 11287 17629 11299 17663
rect 11333 17660 11345 17663
rect 14093 17663 14151 17669
rect 11333 17632 12664 17660
rect 11333 17629 11345 17632
rect 11287 17623 11345 17629
rect 10229 17595 10287 17601
rect 10229 17561 10241 17595
rect 10275 17592 10287 17595
rect 10686 17592 10692 17604
rect 10275 17564 10692 17592
rect 10275 17561 10287 17564
rect 10229 17555 10287 17561
rect 10686 17552 10692 17564
rect 10744 17592 10750 17604
rect 10888 17592 10916 17623
rect 10744 17564 10916 17592
rect 11057 17595 11115 17601
rect 10744 17552 10750 17564
rect 11057 17561 11069 17595
rect 11103 17561 11115 17595
rect 11057 17555 11115 17561
rect 7374 17484 7380 17536
rect 7432 17524 7438 17536
rect 9306 17524 9312 17536
rect 7432 17496 9312 17524
rect 7432 17484 7438 17496
rect 9306 17484 9312 17496
rect 9364 17484 9370 17536
rect 9858 17484 9864 17536
rect 9916 17484 9922 17536
rect 10321 17527 10379 17533
rect 10321 17493 10333 17527
rect 10367 17524 10379 17527
rect 10870 17524 10876 17536
rect 10367 17496 10876 17524
rect 10367 17493 10379 17496
rect 10321 17487 10379 17493
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 11072 17524 11100 17555
rect 11146 17552 11152 17604
rect 11204 17552 11210 17604
rect 11793 17595 11851 17601
rect 11256 17564 11652 17592
rect 11256 17524 11284 17564
rect 11624 17536 11652 17564
rect 11793 17561 11805 17595
rect 11839 17561 11851 17595
rect 11793 17555 11851 17561
rect 11072 17496 11284 17524
rect 11422 17484 11428 17536
rect 11480 17484 11486 17536
rect 11606 17484 11612 17536
rect 11664 17484 11670 17536
rect 11808 17524 11836 17555
rect 12434 17524 12440 17536
rect 11808 17496 12440 17524
rect 12434 17484 12440 17496
rect 12492 17524 12498 17536
rect 12636 17533 12664 17632
rect 14093 17629 14105 17663
rect 14139 17660 14151 17663
rect 14918 17660 14924 17672
rect 14139 17632 14924 17660
rect 14139 17629 14151 17632
rect 14093 17623 14151 17629
rect 14918 17620 14924 17632
rect 14976 17620 14982 17672
rect 16758 17620 16764 17672
rect 16816 17660 16822 17672
rect 17221 17663 17279 17669
rect 17221 17660 17233 17663
rect 16816 17632 17233 17660
rect 16816 17620 16822 17632
rect 17221 17629 17233 17632
rect 17267 17629 17279 17663
rect 18340 17660 18368 17759
rect 22066 17728 22094 17836
rect 22370 17824 22376 17876
rect 22428 17864 22434 17876
rect 24857 17867 24915 17873
rect 24857 17864 24869 17867
rect 22428 17836 24869 17864
rect 22428 17824 22434 17836
rect 24857 17833 24869 17836
rect 24903 17833 24915 17867
rect 24857 17827 24915 17833
rect 25406 17824 25412 17876
rect 25464 17864 25470 17876
rect 25685 17867 25743 17873
rect 25685 17864 25697 17867
rect 25464 17836 25697 17864
rect 25464 17824 25470 17836
rect 25222 17796 25228 17808
rect 25056 17768 25228 17796
rect 24854 17728 24860 17740
rect 22066 17700 24860 17728
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 25056 17737 25084 17768
rect 25222 17756 25228 17768
rect 25280 17756 25286 17808
rect 25016 17731 25084 17737
rect 25016 17697 25028 17731
rect 25062 17697 25084 17731
rect 25016 17691 25084 17697
rect 18509 17663 18567 17669
rect 18509 17660 18521 17663
rect 18340 17632 18521 17660
rect 17221 17623 17279 17629
rect 18509 17629 18521 17632
rect 18555 17629 18567 17663
rect 18509 17623 18567 17629
rect 19337 17663 19395 17669
rect 19337 17629 19349 17663
rect 19383 17629 19395 17663
rect 19337 17623 19395 17629
rect 14360 17595 14418 17601
rect 14360 17561 14372 17595
rect 14406 17592 14418 17595
rect 14642 17592 14648 17604
rect 14406 17564 14648 17592
rect 14406 17561 14418 17564
rect 14360 17555 14418 17561
rect 14642 17552 14648 17564
rect 14700 17552 14706 17604
rect 17494 17552 17500 17604
rect 17552 17592 17558 17604
rect 19352 17592 19380 17623
rect 22278 17620 22284 17672
rect 22336 17620 22342 17672
rect 17552 17564 19380 17592
rect 19604 17595 19662 17601
rect 17552 17552 17558 17564
rect 19604 17561 19616 17595
rect 19650 17592 19662 17595
rect 19886 17592 19892 17604
rect 19650 17564 19892 17592
rect 19650 17561 19662 17564
rect 19604 17555 19662 17561
rect 19886 17552 19892 17564
rect 19944 17552 19950 17604
rect 22462 17592 22468 17604
rect 19996 17564 22468 17592
rect 12621 17527 12679 17533
rect 12492 17496 12537 17524
rect 12492 17484 12498 17496
rect 12621 17493 12633 17527
rect 12667 17524 12679 17527
rect 12986 17524 12992 17536
rect 12667 17496 12992 17524
rect 12667 17493 12679 17496
rect 12621 17487 12679 17493
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 14274 17484 14280 17536
rect 14332 17524 14338 17536
rect 14826 17524 14832 17536
rect 14332 17496 14832 17524
rect 14332 17484 14338 17496
rect 14826 17484 14832 17496
rect 14884 17524 14890 17536
rect 15473 17527 15531 17533
rect 15473 17524 15485 17527
rect 14884 17496 15485 17524
rect 14884 17484 14890 17496
rect 15473 17493 15485 17496
rect 15519 17493 15531 17527
rect 15473 17487 15531 17493
rect 17586 17484 17592 17536
rect 17644 17524 17650 17536
rect 17681 17527 17739 17533
rect 17681 17524 17693 17527
rect 17644 17496 17693 17524
rect 17644 17484 17650 17496
rect 17681 17493 17693 17496
rect 17727 17493 17739 17527
rect 17681 17487 17739 17493
rect 18693 17527 18751 17533
rect 18693 17493 18705 17527
rect 18739 17524 18751 17527
rect 18966 17524 18972 17536
rect 18739 17496 18972 17524
rect 18739 17493 18751 17496
rect 18693 17487 18751 17493
rect 18966 17484 18972 17496
rect 19024 17524 19030 17536
rect 19996 17524 20024 17564
rect 22462 17552 22468 17564
rect 22520 17592 22526 17604
rect 24946 17592 24952 17604
rect 22520 17564 24952 17592
rect 22520 17552 22526 17564
rect 24946 17552 24952 17564
rect 25004 17552 25010 17604
rect 25056 17592 25084 17691
rect 25130 17688 25136 17740
rect 25188 17688 25194 17740
rect 25516 17737 25544 17836
rect 25685 17833 25697 17836
rect 25731 17833 25743 17867
rect 25685 17827 25743 17833
rect 25777 17867 25835 17873
rect 25777 17833 25789 17867
rect 25823 17864 25835 17867
rect 25866 17864 25872 17876
rect 25823 17836 25872 17864
rect 25823 17833 25835 17836
rect 25777 17827 25835 17833
rect 25866 17824 25872 17836
rect 25924 17824 25930 17876
rect 25958 17824 25964 17876
rect 26016 17824 26022 17876
rect 26142 17824 26148 17876
rect 26200 17864 26206 17876
rect 26421 17867 26479 17873
rect 26421 17864 26433 17867
rect 26200 17836 26433 17864
rect 26200 17824 26206 17836
rect 26421 17833 26433 17836
rect 26467 17833 26479 17867
rect 26421 17827 26479 17833
rect 29178 17824 29184 17876
rect 29236 17864 29242 17876
rect 29917 17867 29975 17873
rect 29917 17864 29929 17867
rect 29236 17836 29929 17864
rect 29236 17824 29242 17836
rect 29917 17833 29929 17836
rect 29963 17833 29975 17867
rect 29917 17827 29975 17833
rect 34514 17824 34520 17876
rect 34572 17824 34578 17876
rect 26053 17799 26111 17805
rect 26053 17796 26065 17799
rect 25976 17768 26065 17796
rect 25501 17731 25559 17737
rect 25501 17697 25513 17731
rect 25547 17697 25559 17731
rect 25501 17691 25559 17697
rect 25148 17660 25176 17688
rect 25976 17669 26004 17768
rect 26053 17765 26065 17768
rect 26099 17765 26111 17799
rect 28258 17796 28264 17808
rect 26053 17759 26111 17765
rect 26896 17768 28264 17796
rect 26326 17688 26332 17740
rect 26384 17728 26390 17740
rect 26896 17737 26924 17768
rect 28258 17756 28264 17768
rect 28316 17796 28322 17808
rect 31202 17796 31208 17808
rect 28316 17768 31208 17796
rect 28316 17756 28322 17768
rect 26789 17731 26847 17737
rect 26789 17728 26801 17731
rect 26384 17700 26801 17728
rect 26384 17688 26390 17700
rect 26789 17697 26801 17700
rect 26835 17697 26847 17731
rect 26789 17691 26847 17697
rect 26881 17731 26939 17737
rect 26881 17697 26893 17731
rect 26927 17697 26939 17731
rect 26881 17691 26939 17697
rect 27062 17688 27068 17740
rect 27120 17688 27126 17740
rect 27338 17688 27344 17740
rect 27396 17688 27402 17740
rect 27614 17728 27620 17740
rect 27448 17700 27620 17728
rect 25961 17663 26019 17669
rect 25961 17660 25973 17663
rect 25148 17632 25973 17660
rect 25961 17629 25973 17632
rect 26007 17629 26019 17663
rect 25961 17623 26019 17629
rect 26237 17663 26295 17669
rect 26237 17629 26249 17663
rect 26283 17660 26295 17663
rect 26418 17660 26424 17672
rect 26283 17632 26424 17660
rect 26283 17629 26295 17632
rect 26237 17623 26295 17629
rect 26418 17620 26424 17632
rect 26476 17660 26482 17672
rect 26605 17663 26663 17669
rect 26605 17660 26617 17663
rect 26476 17632 26617 17660
rect 26476 17620 26482 17632
rect 26605 17629 26617 17632
rect 26651 17629 26663 17663
rect 26605 17623 26663 17629
rect 26697 17663 26755 17669
rect 26697 17629 26709 17663
rect 26743 17629 26755 17663
rect 26697 17623 26755 17629
rect 25593 17595 25651 17601
rect 25593 17592 25605 17595
rect 25056 17564 25605 17592
rect 25593 17561 25605 17564
rect 25639 17561 25651 17595
rect 25593 17555 25651 17561
rect 19024 17496 20024 17524
rect 19024 17484 19030 17496
rect 20714 17484 20720 17536
rect 20772 17484 20778 17536
rect 22094 17484 22100 17536
rect 22152 17524 22158 17536
rect 22738 17524 22744 17536
rect 22152 17496 22744 17524
rect 22152 17484 22158 17496
rect 22738 17484 22744 17496
rect 22796 17484 22802 17536
rect 23934 17484 23940 17536
rect 23992 17524 23998 17536
rect 24118 17524 24124 17536
rect 23992 17496 24124 17524
rect 23992 17484 23998 17496
rect 24118 17484 24124 17496
rect 24176 17524 24182 17536
rect 25130 17524 25136 17536
rect 24176 17496 25136 17524
rect 24176 17484 24182 17496
rect 25130 17484 25136 17496
rect 25188 17484 25194 17536
rect 25225 17527 25283 17533
rect 25225 17493 25237 17527
rect 25271 17524 25283 17527
rect 25314 17524 25320 17536
rect 25271 17496 25320 17524
rect 25271 17493 25283 17496
rect 25225 17487 25283 17493
rect 25314 17484 25320 17496
rect 25372 17484 25378 17536
rect 26620 17524 26648 17623
rect 26712 17592 26740 17623
rect 27448 17601 27476 17700
rect 27614 17688 27620 17700
rect 27672 17688 27678 17740
rect 29546 17728 29552 17740
rect 28000 17700 29552 17728
rect 27706 17620 27712 17672
rect 27764 17660 27770 17672
rect 28000 17669 28028 17700
rect 29546 17688 29552 17700
rect 29604 17688 29610 17740
rect 30006 17688 30012 17740
rect 30064 17688 30070 17740
rect 27985 17663 28043 17669
rect 27764 17632 27936 17660
rect 27764 17620 27770 17632
rect 27433 17595 27491 17601
rect 27433 17592 27445 17595
rect 26712 17564 27445 17592
rect 27433 17561 27445 17564
rect 27479 17561 27491 17595
rect 27550 17595 27608 17601
rect 27550 17592 27562 17595
rect 27433 17555 27491 17561
rect 27540 17561 27562 17592
rect 27596 17592 27608 17595
rect 27908 17592 27936 17632
rect 27985 17629 27997 17663
rect 28031 17629 28043 17663
rect 27985 17623 28043 17629
rect 28442 17620 28448 17672
rect 28500 17660 28506 17672
rect 29089 17663 29147 17669
rect 29089 17660 29101 17663
rect 28500 17632 29101 17660
rect 28500 17620 28506 17632
rect 29089 17629 29101 17632
rect 29135 17629 29147 17663
rect 29089 17623 29147 17629
rect 29273 17663 29331 17669
rect 29273 17629 29285 17663
rect 29319 17660 29331 17663
rect 29638 17660 29644 17672
rect 29319 17632 29644 17660
rect 29319 17629 29331 17632
rect 29273 17623 29331 17629
rect 28258 17592 28264 17604
rect 27596 17564 27844 17592
rect 27908 17564 28264 17592
rect 27596 17561 27608 17564
rect 27540 17555 27608 17561
rect 27540 17524 27568 17555
rect 26620 17496 27568 17524
rect 27706 17484 27712 17536
rect 27764 17484 27770 17536
rect 27816 17533 27844 17564
rect 28258 17552 28264 17564
rect 28316 17552 28322 17604
rect 28905 17595 28963 17601
rect 28905 17561 28917 17595
rect 28951 17592 28963 17595
rect 29288 17592 29316 17623
rect 29638 17620 29644 17632
rect 29696 17660 29702 17672
rect 29733 17663 29791 17669
rect 29733 17660 29745 17663
rect 29696 17632 29745 17660
rect 29696 17620 29702 17632
rect 29733 17629 29745 17632
rect 29779 17629 29791 17663
rect 29733 17623 29791 17629
rect 29822 17620 29828 17672
rect 29880 17660 29886 17672
rect 29917 17663 29975 17669
rect 29917 17660 29929 17663
rect 29880 17632 29929 17660
rect 29880 17620 29886 17632
rect 29917 17629 29929 17632
rect 29963 17629 29975 17663
rect 29917 17623 29975 17629
rect 30190 17620 30196 17672
rect 30248 17620 30254 17672
rect 30926 17620 30932 17672
rect 30984 17660 30990 17672
rect 31128 17669 31156 17768
rect 31202 17756 31208 17768
rect 31260 17756 31266 17808
rect 31297 17799 31355 17805
rect 31297 17765 31309 17799
rect 31343 17765 31355 17799
rect 31297 17759 31355 17765
rect 31021 17663 31079 17669
rect 31021 17660 31033 17663
rect 30984 17632 31033 17660
rect 30984 17620 30990 17632
rect 31021 17629 31033 17632
rect 31067 17629 31079 17663
rect 31021 17623 31079 17629
rect 31113 17663 31171 17669
rect 31113 17629 31125 17663
rect 31159 17629 31171 17663
rect 31312 17660 31340 17759
rect 33045 17731 33103 17737
rect 33045 17697 33057 17731
rect 33091 17728 33103 17731
rect 33778 17728 33784 17740
rect 33091 17700 33784 17728
rect 33091 17697 33103 17700
rect 33045 17691 33103 17697
rect 33778 17688 33784 17700
rect 33836 17688 33842 17740
rect 31389 17663 31447 17669
rect 31389 17660 31401 17663
rect 31312 17632 31401 17660
rect 31113 17623 31171 17629
rect 31389 17629 31401 17632
rect 31435 17629 31447 17663
rect 31389 17623 31447 17629
rect 31570 17620 31576 17672
rect 31628 17620 31634 17672
rect 32122 17620 32128 17672
rect 32180 17660 32186 17672
rect 32674 17660 32680 17672
rect 32180 17632 32680 17660
rect 32180 17620 32186 17632
rect 32674 17620 32680 17632
rect 32732 17660 32738 17672
rect 32769 17663 32827 17669
rect 32769 17660 32781 17663
rect 32732 17632 32781 17660
rect 32732 17620 32738 17632
rect 32769 17629 32781 17632
rect 32815 17629 32827 17663
rect 32769 17623 32827 17629
rect 28951 17564 29316 17592
rect 28951 17561 28963 17564
rect 28905 17555 28963 17561
rect 31294 17552 31300 17604
rect 31352 17552 31358 17604
rect 33134 17552 33140 17604
rect 33192 17592 33198 17604
rect 33192 17564 33534 17592
rect 33192 17552 33198 17564
rect 27801 17527 27859 17533
rect 27801 17493 27813 17527
rect 27847 17493 27859 17527
rect 27801 17487 27859 17493
rect 28994 17484 29000 17536
rect 29052 17524 29058 17536
rect 29549 17527 29607 17533
rect 29549 17524 29561 17527
rect 29052 17496 29561 17524
rect 29052 17484 29058 17496
rect 29549 17493 29561 17496
rect 29595 17493 29607 17527
rect 29549 17487 29607 17493
rect 30377 17527 30435 17533
rect 30377 17493 30389 17527
rect 30423 17524 30435 17527
rect 31018 17524 31024 17536
rect 30423 17496 31024 17524
rect 30423 17493 30435 17496
rect 30377 17487 30435 17493
rect 31018 17484 31024 17496
rect 31076 17484 31082 17536
rect 31478 17484 31484 17536
rect 31536 17484 31542 17536
rect 1104 17434 35328 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35328 17434
rect 1104 17360 35328 17382
rect 4893 17323 4951 17329
rect 4893 17289 4905 17323
rect 4939 17289 4951 17323
rect 4893 17283 4951 17289
rect 4614 17212 4620 17264
rect 4672 17252 4678 17264
rect 4908 17252 4936 17283
rect 4982 17280 4988 17332
rect 5040 17320 5046 17332
rect 5258 17320 5264 17332
rect 5040 17292 5264 17320
rect 5040 17280 5046 17292
rect 5258 17280 5264 17292
rect 5316 17320 5322 17332
rect 5316 17292 7604 17320
rect 5316 17280 5322 17292
rect 7469 17255 7527 17261
rect 7469 17252 7481 17255
rect 4672 17224 7481 17252
rect 4672 17212 4678 17224
rect 7469 17221 7481 17224
rect 7515 17221 7527 17255
rect 7469 17215 7527 17221
rect 3780 17187 3838 17193
rect 3780 17153 3792 17187
rect 3826 17184 3838 17187
rect 4062 17184 4068 17196
rect 3826 17156 4068 17184
rect 3826 17153 3838 17156
rect 3780 17147 3838 17153
rect 4062 17144 4068 17156
rect 4120 17144 4126 17196
rect 6730 17144 6736 17196
rect 6788 17184 6794 17196
rect 7576 17193 7604 17292
rect 7742 17280 7748 17332
rect 7800 17280 7806 17332
rect 8297 17323 8355 17329
rect 8297 17320 8309 17323
rect 8036 17292 8309 17320
rect 8036 17261 8064 17292
rect 8297 17289 8309 17292
rect 8343 17320 8355 17323
rect 9490 17320 9496 17332
rect 8343 17292 9496 17320
rect 8343 17289 8355 17292
rect 8297 17283 8355 17289
rect 9490 17280 9496 17292
rect 9548 17280 9554 17332
rect 10686 17280 10692 17332
rect 10744 17280 10750 17332
rect 11146 17280 11152 17332
rect 11204 17320 11210 17332
rect 12250 17320 12256 17332
rect 11204 17292 12256 17320
rect 11204 17280 11210 17292
rect 12250 17280 12256 17292
rect 12308 17320 12314 17332
rect 12897 17323 12955 17329
rect 12897 17320 12909 17323
rect 12308 17292 12909 17320
rect 12308 17280 12314 17292
rect 12897 17289 12909 17292
rect 12943 17289 12955 17323
rect 12897 17283 12955 17289
rect 14274 17280 14280 17332
rect 14332 17280 14338 17332
rect 14642 17280 14648 17332
rect 14700 17280 14706 17332
rect 14734 17280 14740 17332
rect 14792 17320 14798 17332
rect 14921 17323 14979 17329
rect 14921 17320 14933 17323
rect 14792 17292 14933 17320
rect 14792 17280 14798 17292
rect 14921 17289 14933 17292
rect 14967 17320 14979 17323
rect 15102 17320 15108 17332
rect 14967 17292 15108 17320
rect 14967 17289 14979 17292
rect 14921 17283 14979 17289
rect 15102 17280 15108 17292
rect 15160 17280 15166 17332
rect 19153 17323 19211 17329
rect 19153 17289 19165 17323
rect 19199 17289 19211 17323
rect 19153 17283 19211 17289
rect 8021 17255 8079 17261
rect 8021 17221 8033 17255
rect 8067 17221 8079 17255
rect 8021 17215 8079 17221
rect 9576 17255 9634 17261
rect 9576 17221 9588 17255
rect 9622 17252 9634 17255
rect 9858 17252 9864 17264
rect 9622 17224 9864 17252
rect 9622 17221 9634 17224
rect 9576 17215 9634 17221
rect 9858 17212 9864 17224
rect 9916 17212 9922 17264
rect 13078 17252 13084 17264
rect 11532 17224 13084 17252
rect 7193 17187 7251 17193
rect 7193 17184 7205 17187
rect 6788 17156 7205 17184
rect 6788 17144 6794 17156
rect 7193 17153 7205 17156
rect 7239 17153 7251 17187
rect 7193 17147 7251 17153
rect 7377 17187 7435 17193
rect 7377 17153 7389 17187
rect 7423 17153 7435 17187
rect 7377 17147 7435 17153
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17184 7619 17187
rect 7837 17187 7895 17193
rect 7837 17184 7849 17187
rect 7607 17156 7849 17184
rect 7607 17153 7619 17156
rect 7561 17147 7619 17153
rect 7837 17153 7849 17156
rect 7883 17153 7895 17187
rect 7837 17147 7895 17153
rect 3510 17076 3516 17128
rect 3568 17076 3574 17128
rect 6822 17076 6828 17128
rect 6880 17076 6886 17128
rect 7006 17076 7012 17128
rect 7064 17076 7070 17128
rect 5718 17008 5724 17060
rect 5776 17048 5782 17060
rect 7392 17048 7420 17147
rect 9306 17144 9312 17196
rect 9364 17144 9370 17196
rect 11532 17128 11560 17224
rect 13078 17212 13084 17224
rect 13136 17212 13142 17264
rect 14182 17212 14188 17264
rect 14240 17252 14246 17264
rect 19168 17252 19196 17283
rect 19886 17280 19892 17332
rect 19944 17280 19950 17332
rect 21542 17280 21548 17332
rect 21600 17320 21606 17332
rect 21600 17292 22232 17320
rect 21600 17280 21606 17292
rect 19334 17252 19340 17264
rect 14240 17224 14780 17252
rect 14240 17212 14246 17224
rect 14752 17196 14780 17224
rect 15028 17224 18920 17252
rect 19168 17224 19340 17252
rect 11790 17193 11796 17196
rect 11784 17147 11796 17193
rect 11790 17144 11796 17147
rect 11848 17144 11854 17196
rect 12066 17144 12072 17196
rect 12124 17184 12130 17196
rect 14642 17184 14648 17196
rect 12124 17156 14648 17184
rect 12124 17144 12130 17156
rect 14642 17144 14648 17156
rect 14700 17144 14706 17196
rect 14734 17144 14740 17196
rect 14792 17144 14798 17196
rect 11514 17076 11520 17128
rect 11572 17076 11578 17128
rect 13814 17076 13820 17128
rect 13872 17116 13878 17128
rect 14090 17116 14096 17128
rect 13872 17088 14096 17116
rect 13872 17076 13878 17088
rect 14090 17076 14096 17088
rect 14148 17076 14154 17128
rect 14182 17076 14188 17128
rect 14240 17076 14246 17128
rect 14550 17076 14556 17128
rect 14608 17116 14614 17128
rect 15028 17116 15056 17224
rect 15372 17187 15430 17193
rect 15372 17153 15384 17187
rect 15418 17184 15430 17187
rect 15746 17184 15752 17196
rect 15418 17156 15752 17184
rect 15418 17153 15430 17156
rect 15372 17147 15430 17153
rect 15746 17144 15752 17156
rect 15804 17144 15810 17196
rect 17494 17144 17500 17196
rect 17552 17144 17558 17196
rect 17764 17187 17822 17193
rect 17764 17153 17776 17187
rect 17810 17184 17822 17187
rect 18046 17184 18052 17196
rect 17810 17156 18052 17184
rect 17810 17153 17822 17156
rect 17764 17147 17822 17153
rect 18046 17144 18052 17156
rect 18104 17144 18110 17196
rect 14608 17088 15056 17116
rect 15105 17119 15163 17125
rect 14608 17076 14614 17088
rect 15105 17085 15117 17119
rect 15151 17085 15163 17119
rect 15105 17079 15163 17085
rect 8478 17048 8484 17060
rect 5776 17020 6500 17048
rect 7392 17020 8484 17048
rect 5776 17008 5782 17020
rect 6362 16940 6368 16992
rect 6420 16940 6426 16992
rect 6472 16980 6500 17020
rect 8478 17008 8484 17020
rect 8536 17048 8542 17060
rect 9030 17048 9036 17060
rect 8536 17020 9036 17048
rect 8536 17008 8542 17020
rect 9030 17008 9036 17020
rect 9088 17008 9094 17060
rect 10244 17020 10916 17048
rect 10244 16980 10272 17020
rect 6472 16952 10272 16980
rect 10318 16940 10324 16992
rect 10376 16980 10382 16992
rect 10781 16983 10839 16989
rect 10781 16980 10793 16983
rect 10376 16952 10793 16980
rect 10376 16940 10382 16952
rect 10781 16949 10793 16952
rect 10827 16949 10839 16983
rect 10888 16980 10916 17020
rect 13078 17008 13084 17060
rect 13136 17048 13142 17060
rect 15120 17048 15148 17079
rect 16574 17048 16580 17060
rect 13136 17020 15148 17048
rect 16408 17020 16580 17048
rect 13136 17008 13142 17020
rect 16408 16980 16436 17020
rect 16574 17008 16580 17020
rect 16632 17008 16638 17060
rect 18892 17048 18920 17224
rect 19334 17212 19340 17224
rect 19392 17252 19398 17264
rect 20257 17255 20315 17261
rect 20257 17252 20269 17255
rect 19392 17224 20269 17252
rect 19392 17212 19398 17224
rect 20257 17221 20269 17224
rect 20303 17252 20315 17255
rect 20530 17252 20536 17264
rect 20303 17224 20536 17252
rect 20303 17221 20315 17224
rect 20257 17215 20315 17221
rect 20530 17212 20536 17224
rect 20588 17252 20594 17264
rect 20588 17224 21956 17252
rect 20588 17212 20594 17224
rect 18966 17144 18972 17196
rect 19024 17144 19030 17196
rect 20349 17187 20407 17193
rect 20349 17153 20361 17187
rect 20395 17184 20407 17187
rect 20714 17184 20720 17196
rect 20395 17156 20720 17184
rect 20395 17153 20407 17156
rect 20349 17147 20407 17153
rect 20714 17144 20720 17156
rect 20772 17184 20778 17196
rect 21821 17187 21879 17193
rect 21821 17184 21833 17187
rect 20772 17156 21833 17184
rect 20772 17144 20778 17156
rect 21821 17153 21833 17156
rect 21867 17153 21879 17187
rect 21821 17147 21879 17153
rect 19794 17076 19800 17128
rect 19852 17116 19858 17128
rect 20441 17119 20499 17125
rect 20441 17116 20453 17119
rect 19852 17088 20453 17116
rect 19852 17076 19858 17088
rect 20441 17085 20453 17088
rect 20487 17116 20499 17119
rect 20809 17119 20867 17125
rect 20809 17116 20821 17119
rect 20487 17088 20821 17116
rect 20487 17085 20499 17088
rect 20441 17079 20499 17085
rect 20809 17085 20821 17088
rect 20855 17085 20867 17119
rect 20809 17079 20867 17085
rect 21542 17048 21548 17060
rect 18892 17020 21548 17048
rect 21542 17008 21548 17020
rect 21600 17008 21606 17060
rect 10888 16952 16436 16980
rect 10781 16943 10839 16949
rect 16482 16940 16488 16992
rect 16540 16940 16546 16992
rect 18874 16940 18880 16992
rect 18932 16940 18938 16992
rect 20162 16940 20168 16992
rect 20220 16980 20226 16992
rect 20990 16980 20996 16992
rect 20220 16952 20996 16980
rect 20220 16940 20226 16952
rect 20990 16940 20996 16952
rect 21048 16940 21054 16992
rect 21928 16980 21956 17224
rect 22094 17212 22100 17264
rect 22152 17212 22158 17264
rect 22204 17193 22232 17292
rect 22646 17280 22652 17332
rect 22704 17320 22710 17332
rect 24765 17323 24823 17329
rect 24765 17320 24777 17323
rect 22704 17292 24777 17320
rect 22704 17280 22710 17292
rect 24765 17289 24777 17292
rect 24811 17289 24823 17323
rect 24765 17283 24823 17289
rect 24854 17280 24860 17332
rect 24912 17320 24918 17332
rect 27062 17320 27068 17332
rect 24912 17292 27068 17320
rect 24912 17280 24918 17292
rect 27062 17280 27068 17292
rect 27120 17280 27126 17332
rect 28261 17323 28319 17329
rect 28261 17289 28273 17323
rect 28307 17320 28319 17323
rect 28307 17292 29776 17320
rect 28307 17289 28319 17292
rect 28261 17283 28319 17289
rect 24578 17212 24584 17264
rect 24636 17252 24642 17264
rect 25593 17255 25651 17261
rect 25593 17252 25605 17255
rect 24636 17224 25605 17252
rect 24636 17212 24642 17224
rect 25593 17221 25605 17224
rect 25639 17221 25651 17255
rect 25593 17215 25651 17221
rect 26602 17212 26608 17264
rect 26660 17252 26666 17264
rect 26697 17255 26755 17261
rect 26697 17252 26709 17255
rect 26660 17224 26709 17252
rect 26660 17212 26666 17224
rect 26697 17221 26709 17224
rect 26743 17252 26755 17255
rect 27246 17252 27252 17264
rect 26743 17224 27252 17252
rect 26743 17221 26755 17224
rect 26697 17215 26755 17221
rect 27246 17212 27252 17224
rect 27304 17212 27310 17264
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17184 22063 17187
rect 22189 17187 22247 17193
rect 22051 17156 22140 17184
rect 22051 17153 22063 17156
rect 22005 17147 22063 17153
rect 22112 17116 22140 17156
rect 22189 17153 22201 17187
rect 22235 17153 22247 17187
rect 23106 17184 23112 17196
rect 22189 17147 22247 17153
rect 22296 17156 23112 17184
rect 22296 17116 22324 17156
rect 23106 17144 23112 17156
rect 23164 17144 23170 17196
rect 23382 17144 23388 17196
rect 23440 17144 23446 17196
rect 23845 17187 23903 17193
rect 23845 17153 23857 17187
rect 23891 17153 23903 17187
rect 23845 17147 23903 17153
rect 24673 17187 24731 17193
rect 24673 17153 24685 17187
rect 24719 17153 24731 17187
rect 24673 17147 24731 17153
rect 22112 17088 22324 17116
rect 22370 17076 22376 17128
rect 22428 17116 22434 17128
rect 22557 17119 22615 17125
rect 22557 17116 22569 17119
rect 22428 17088 22569 17116
rect 22428 17076 22434 17088
rect 22557 17085 22569 17088
rect 22603 17085 22615 17119
rect 22557 17079 22615 17085
rect 23860 17048 23888 17147
rect 23934 17076 23940 17128
rect 23992 17076 23998 17128
rect 24026 17076 24032 17128
rect 24084 17076 24090 17128
rect 24578 17076 24584 17128
rect 24636 17116 24642 17128
rect 24688 17116 24716 17147
rect 25130 17144 25136 17196
rect 25188 17184 25194 17196
rect 25869 17187 25927 17193
rect 25869 17184 25881 17187
rect 25188 17156 25881 17184
rect 25188 17144 25194 17156
rect 25869 17153 25881 17156
rect 25915 17153 25927 17187
rect 25869 17147 25927 17153
rect 26326 17144 26332 17196
rect 26384 17184 26390 17196
rect 27157 17187 27215 17193
rect 27157 17184 27169 17187
rect 26384 17156 27169 17184
rect 26384 17144 26390 17156
rect 27157 17153 27169 17156
rect 27203 17184 27215 17187
rect 27203 17156 27476 17184
rect 27203 17153 27215 17156
rect 27157 17147 27215 17153
rect 24636 17088 24716 17116
rect 24857 17119 24915 17125
rect 24636 17076 24642 17088
rect 24857 17085 24869 17119
rect 24903 17085 24915 17119
rect 24857 17079 24915 17085
rect 24872 17048 24900 17079
rect 24946 17076 24952 17128
rect 25004 17116 25010 17128
rect 27338 17116 27344 17128
rect 25004 17088 27344 17116
rect 25004 17076 25010 17088
rect 27338 17076 27344 17088
rect 27396 17076 27402 17128
rect 25317 17051 25375 17057
rect 25317 17048 25329 17051
rect 22103 17020 23888 17048
rect 24228 17020 25329 17048
rect 22103 16980 22131 17020
rect 21928 16952 22131 16980
rect 22370 16940 22376 16992
rect 22428 16940 22434 16992
rect 23474 16940 23480 16992
rect 23532 16940 23538 16992
rect 23842 16940 23848 16992
rect 23900 16980 23906 16992
rect 24228 16980 24256 17020
rect 25317 17017 25329 17020
rect 25363 17048 25375 17051
rect 26053 17051 26111 17057
rect 26053 17048 26065 17051
rect 25363 17020 26065 17048
rect 25363 17017 25375 17020
rect 25317 17011 25375 17017
rect 26053 17017 26065 17020
rect 26099 17048 26111 17051
rect 26237 17051 26295 17057
rect 26237 17048 26249 17051
rect 26099 17020 26249 17048
rect 26099 17017 26111 17020
rect 26053 17011 26111 17017
rect 26237 17017 26249 17020
rect 26283 17017 26295 17051
rect 26237 17011 26295 17017
rect 26878 17008 26884 17060
rect 26936 17048 26942 17060
rect 26973 17051 27031 17057
rect 26973 17048 26985 17051
rect 26936 17020 26985 17048
rect 26936 17008 26942 17020
rect 26973 17017 26985 17020
rect 27019 17017 27031 17051
rect 26973 17011 27031 17017
rect 23900 16952 24256 16980
rect 23900 16940 23906 16952
rect 24302 16940 24308 16992
rect 24360 16940 24366 16992
rect 25590 16940 25596 16992
rect 25648 16980 25654 16992
rect 25685 16983 25743 16989
rect 25685 16980 25697 16983
rect 25648 16952 25697 16980
rect 25648 16940 25654 16952
rect 25685 16949 25697 16952
rect 25731 16980 25743 16983
rect 26421 16983 26479 16989
rect 26421 16980 26433 16983
rect 25731 16952 26433 16980
rect 25731 16949 25743 16952
rect 25685 16943 25743 16949
rect 26421 16949 26433 16952
rect 26467 16949 26479 16983
rect 27448 16980 27476 17156
rect 27798 17076 27804 17128
rect 27856 17116 27862 17128
rect 28353 17119 28411 17125
rect 28353 17116 28365 17119
rect 27856 17088 28365 17116
rect 27856 17076 27862 17088
rect 28353 17085 28365 17088
rect 28399 17085 28411 17119
rect 28353 17079 28411 17085
rect 28626 17076 28632 17128
rect 28684 17076 28690 17128
rect 29748 17116 29776 17292
rect 30098 17280 30104 17332
rect 30156 17280 30162 17332
rect 30926 17280 30932 17332
rect 30984 17320 30990 17332
rect 31294 17320 31300 17332
rect 30984 17292 31300 17320
rect 30984 17280 30990 17292
rect 31294 17280 31300 17292
rect 31352 17280 31358 17332
rect 29822 17116 29828 17128
rect 29748 17088 29828 17116
rect 29822 17076 29828 17088
rect 29880 17076 29886 17128
rect 29270 16980 29276 16992
rect 27448 16952 29276 16980
rect 26421 16943 26479 16949
rect 29270 16940 29276 16952
rect 29328 16940 29334 16992
rect 1104 16890 35328 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 35328 16890
rect 1104 16816 35328 16838
rect 5350 16736 5356 16788
rect 5408 16776 5414 16788
rect 5534 16776 5540 16788
rect 5408 16748 5540 16776
rect 5408 16736 5414 16748
rect 5534 16736 5540 16748
rect 5592 16736 5598 16788
rect 6730 16736 6736 16788
rect 6788 16736 6794 16788
rect 7006 16736 7012 16788
rect 7064 16776 7070 16788
rect 7285 16779 7343 16785
rect 7285 16776 7297 16779
rect 7064 16748 7297 16776
rect 7064 16736 7070 16748
rect 7285 16745 7297 16748
rect 7331 16776 7343 16779
rect 9674 16776 9680 16788
rect 7331 16748 9680 16776
rect 7331 16745 7343 16748
rect 7285 16739 7343 16745
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 12434 16776 12440 16788
rect 11808 16748 12440 16776
rect 5350 16640 5356 16652
rect 4080 16612 5356 16640
rect 1394 16532 1400 16584
rect 1452 16572 1458 16584
rect 1673 16575 1731 16581
rect 1673 16572 1685 16575
rect 1452 16544 1685 16572
rect 1452 16532 1458 16544
rect 1673 16541 1685 16544
rect 1719 16541 1731 16575
rect 1673 16535 1731 16541
rect 2774 16464 2780 16516
rect 2832 16504 2838 16516
rect 3145 16507 3203 16513
rect 3145 16504 3157 16507
rect 2832 16476 3157 16504
rect 2832 16464 2838 16476
rect 3145 16473 3157 16476
rect 3191 16504 3203 16507
rect 3510 16504 3516 16516
rect 3191 16476 3516 16504
rect 3191 16473 3203 16476
rect 3145 16467 3203 16473
rect 3510 16464 3516 16476
rect 3568 16504 3574 16516
rect 4080 16513 4108 16612
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 7374 16600 7380 16652
rect 7432 16600 7438 16652
rect 9306 16600 9312 16652
rect 9364 16640 9370 16652
rect 11149 16643 11207 16649
rect 11149 16640 11161 16643
rect 9364 16612 11161 16640
rect 9364 16600 9370 16612
rect 11149 16609 11161 16612
rect 11195 16640 11207 16643
rect 11514 16640 11520 16652
rect 11195 16612 11520 16640
rect 11195 16609 11207 16612
rect 11149 16603 11207 16609
rect 11514 16600 11520 16612
rect 11572 16600 11578 16652
rect 11808 16649 11836 16748
rect 12434 16736 12440 16748
rect 12492 16776 12498 16788
rect 12492 16748 13952 16776
rect 12492 16736 12498 16748
rect 13630 16668 13636 16720
rect 13688 16668 13694 16720
rect 11793 16643 11851 16649
rect 11793 16609 11805 16643
rect 11839 16609 11851 16643
rect 11793 16603 11851 16609
rect 5620 16575 5678 16581
rect 5620 16541 5632 16575
rect 5666 16572 5678 16575
rect 6362 16572 6368 16584
rect 5666 16544 6368 16572
rect 5666 16541 5678 16544
rect 5620 16535 5678 16541
rect 6362 16532 6368 16544
rect 6420 16532 6426 16584
rect 10413 16575 10471 16581
rect 10413 16572 10425 16575
rect 6472 16544 10425 16572
rect 4065 16507 4123 16513
rect 4065 16504 4077 16507
rect 3568 16476 4077 16504
rect 3568 16464 3574 16476
rect 4065 16473 4077 16476
rect 4111 16473 4123 16507
rect 4065 16467 4123 16473
rect 4893 16507 4951 16513
rect 4893 16473 4905 16507
rect 4939 16473 4951 16507
rect 4893 16467 4951 16473
rect 1578 16396 1584 16448
rect 1636 16396 1642 16448
rect 4908 16436 4936 16467
rect 6472 16448 6500 16544
rect 10413 16541 10425 16544
rect 10459 16572 10471 16575
rect 11425 16575 11483 16581
rect 11425 16572 11437 16575
rect 10459 16544 11437 16572
rect 10459 16541 10471 16544
rect 10413 16535 10471 16541
rect 11425 16541 11437 16544
rect 11471 16572 11483 16575
rect 11808 16572 11836 16603
rect 11882 16600 11888 16652
rect 11940 16640 11946 16652
rect 13814 16640 13820 16652
rect 11940 16612 13820 16640
rect 11940 16600 11946 16612
rect 13814 16600 13820 16612
rect 13872 16600 13878 16652
rect 13924 16649 13952 16748
rect 13998 16736 14004 16788
rect 14056 16776 14062 16788
rect 14369 16779 14427 16785
rect 14369 16776 14381 16779
rect 14056 16748 14381 16776
rect 14056 16736 14062 16748
rect 14369 16745 14381 16748
rect 14415 16776 14427 16779
rect 14550 16776 14556 16788
rect 14415 16748 14556 16776
rect 14415 16745 14427 16748
rect 14369 16739 14427 16745
rect 14550 16736 14556 16748
rect 14608 16736 14614 16788
rect 14642 16736 14648 16788
rect 14700 16776 14706 16788
rect 14700 16748 15424 16776
rect 14700 16736 14706 16748
rect 14182 16668 14188 16720
rect 14240 16708 14246 16720
rect 14277 16711 14335 16717
rect 14277 16708 14289 16711
rect 14240 16680 14289 16708
rect 14240 16668 14246 16680
rect 14277 16677 14289 16680
rect 14323 16708 14335 16711
rect 15010 16708 15016 16720
rect 14323 16680 15016 16708
rect 14323 16677 14335 16680
rect 14277 16671 14335 16677
rect 15010 16668 15016 16680
rect 15068 16668 15074 16720
rect 15286 16668 15292 16720
rect 15344 16668 15350 16720
rect 13909 16643 13967 16649
rect 13909 16609 13921 16643
rect 13955 16640 13967 16643
rect 14734 16640 14740 16652
rect 13955 16612 14740 16640
rect 13955 16609 13967 16612
rect 13909 16603 13967 16609
rect 14734 16600 14740 16612
rect 14792 16600 14798 16652
rect 15396 16640 15424 16748
rect 15746 16736 15752 16788
rect 15804 16736 15810 16788
rect 18046 16736 18052 16788
rect 18104 16736 18110 16788
rect 21450 16776 21456 16788
rect 20548 16748 21456 16776
rect 19334 16708 19340 16720
rect 18524 16680 19340 16708
rect 18524 16649 18552 16680
rect 19334 16668 19340 16680
rect 19392 16668 19398 16720
rect 16301 16643 16359 16649
rect 16301 16640 16313 16643
rect 15396 16612 16313 16640
rect 16301 16609 16313 16612
rect 16347 16640 16359 16643
rect 17313 16643 17371 16649
rect 17313 16640 17325 16643
rect 16347 16612 17325 16640
rect 16347 16609 16359 16612
rect 16301 16603 16359 16609
rect 17313 16609 17325 16612
rect 17359 16609 17371 16643
rect 17313 16603 17371 16609
rect 18509 16643 18567 16649
rect 18509 16609 18521 16643
rect 18555 16609 18567 16643
rect 18509 16603 18567 16609
rect 18693 16643 18751 16649
rect 18693 16609 18705 16643
rect 18739 16640 18751 16643
rect 18969 16643 19027 16649
rect 18969 16640 18981 16643
rect 18739 16612 18981 16640
rect 18739 16609 18751 16612
rect 18693 16603 18751 16609
rect 18969 16609 18981 16612
rect 19015 16640 19027 16643
rect 19150 16640 19156 16652
rect 19015 16612 19156 16640
rect 19015 16609 19027 16612
rect 18969 16603 19027 16609
rect 19150 16600 19156 16612
rect 19208 16640 19214 16652
rect 19886 16640 19892 16652
rect 19208 16612 19892 16640
rect 19208 16600 19214 16612
rect 19886 16600 19892 16612
rect 19944 16600 19950 16652
rect 11471 16544 11836 16572
rect 13541 16575 13599 16581
rect 11471 16541 11483 16544
rect 11425 16535 11483 16541
rect 13541 16541 13553 16575
rect 13587 16572 13599 16575
rect 13630 16572 13636 16584
rect 13587 16544 13636 16572
rect 13587 16541 13599 16544
rect 13541 16535 13599 16541
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 14093 16575 14151 16581
rect 14093 16541 14105 16575
rect 14139 16541 14151 16575
rect 14093 16535 14151 16541
rect 7644 16507 7702 16513
rect 7644 16473 7656 16507
rect 7690 16504 7702 16507
rect 8018 16504 8024 16516
rect 7690 16476 8024 16504
rect 7690 16473 7702 16476
rect 7644 16467 7702 16473
rect 8018 16464 8024 16476
rect 8076 16464 8082 16516
rect 11146 16464 11152 16516
rect 11204 16504 11210 16516
rect 14108 16504 14136 16535
rect 14550 16532 14556 16584
rect 14608 16532 14614 16584
rect 14642 16532 14648 16584
rect 14700 16572 14706 16584
rect 14700 16544 14780 16572
rect 14700 16532 14706 16544
rect 14752 16513 14780 16544
rect 14826 16532 14832 16584
rect 14884 16532 14890 16584
rect 14921 16575 14979 16581
rect 14921 16541 14933 16575
rect 14967 16572 14979 16575
rect 15102 16572 15108 16584
rect 14967 16544 15108 16572
rect 14967 16541 14979 16544
rect 14921 16535 14979 16541
rect 15102 16532 15108 16544
rect 15160 16572 15166 16584
rect 15473 16575 15531 16581
rect 15473 16572 15485 16575
rect 15160 16544 15485 16572
rect 15160 16532 15166 16544
rect 15473 16541 15485 16544
rect 15519 16541 15531 16575
rect 15473 16535 15531 16541
rect 15930 16532 15936 16584
rect 15988 16572 15994 16584
rect 16117 16575 16175 16581
rect 16117 16572 16129 16575
rect 15988 16544 16129 16572
rect 15988 16532 15994 16544
rect 16117 16541 16129 16544
rect 16163 16572 16175 16575
rect 16482 16572 16488 16584
rect 16163 16544 16488 16572
rect 16163 16541 16175 16544
rect 16117 16535 16175 16541
rect 16482 16532 16488 16544
rect 16540 16532 16546 16584
rect 16574 16532 16580 16584
rect 16632 16572 16638 16584
rect 17218 16572 17224 16584
rect 16632 16544 17224 16572
rect 16632 16532 16638 16544
rect 17218 16532 17224 16544
rect 17276 16532 17282 16584
rect 18417 16575 18475 16581
rect 18417 16541 18429 16575
rect 18463 16572 18475 16575
rect 18874 16572 18880 16584
rect 18463 16544 18880 16572
rect 18463 16541 18475 16544
rect 18417 16535 18475 16541
rect 18874 16532 18880 16544
rect 18932 16532 18938 16584
rect 20548 16572 20576 16748
rect 21450 16736 21456 16748
rect 21508 16736 21514 16788
rect 22094 16736 22100 16788
rect 22152 16776 22158 16788
rect 22189 16779 22247 16785
rect 22189 16776 22201 16779
rect 22152 16748 22201 16776
rect 22152 16736 22158 16748
rect 22189 16745 22201 16748
rect 22235 16745 22247 16779
rect 22189 16739 22247 16745
rect 27062 16736 27068 16788
rect 27120 16776 27126 16788
rect 27709 16779 27767 16785
rect 27709 16776 27721 16779
rect 27120 16748 27721 16776
rect 27120 16736 27126 16748
rect 27709 16745 27721 16748
rect 27755 16745 27767 16779
rect 27709 16739 27767 16745
rect 28445 16779 28503 16785
rect 28445 16745 28457 16779
rect 28491 16776 28503 16779
rect 28626 16776 28632 16788
rect 28491 16748 28632 16776
rect 28491 16745 28503 16748
rect 28445 16739 28503 16745
rect 28626 16736 28632 16748
rect 28684 16736 28690 16788
rect 29730 16736 29736 16788
rect 29788 16736 29794 16788
rect 30190 16736 30196 16788
rect 30248 16776 30254 16788
rect 30377 16779 30435 16785
rect 30377 16776 30389 16779
rect 30248 16748 30389 16776
rect 30248 16736 30254 16748
rect 30377 16745 30389 16748
rect 30423 16776 30435 16779
rect 30834 16776 30840 16788
rect 30423 16748 30840 16776
rect 30423 16745 30435 16748
rect 30377 16739 30435 16745
rect 30834 16736 30840 16748
rect 30892 16736 30898 16788
rect 23661 16711 23719 16717
rect 23661 16677 23673 16711
rect 23707 16708 23719 16711
rect 23934 16708 23940 16720
rect 23707 16680 23940 16708
rect 23707 16677 23719 16680
rect 23661 16671 23719 16677
rect 23934 16668 23940 16680
rect 23992 16708 23998 16720
rect 25314 16708 25320 16720
rect 23992 16680 25320 16708
rect 23992 16668 23998 16680
rect 25314 16668 25320 16680
rect 25372 16668 25378 16720
rect 26142 16708 26148 16720
rect 25700 16680 26148 16708
rect 20622 16600 20628 16652
rect 20680 16640 20686 16652
rect 20809 16643 20867 16649
rect 20809 16640 20821 16643
rect 20680 16612 20821 16640
rect 20680 16600 20686 16612
rect 20809 16609 20821 16612
rect 20855 16609 20867 16643
rect 20809 16603 20867 16609
rect 23845 16643 23903 16649
rect 23845 16609 23857 16643
rect 23891 16640 23903 16643
rect 24026 16640 24032 16652
rect 23891 16612 24032 16640
rect 23891 16609 23903 16612
rect 23845 16603 23903 16609
rect 24026 16600 24032 16612
rect 24084 16600 24090 16652
rect 24394 16600 24400 16652
rect 24452 16600 24458 16652
rect 24688 16612 25544 16640
rect 19536 16544 20576 16572
rect 21076 16575 21134 16581
rect 11204 16476 14136 16504
rect 14737 16507 14795 16513
rect 11204 16464 11210 16476
rect 14737 16473 14749 16507
rect 14783 16473 14795 16507
rect 14737 16467 14795 16473
rect 5077 16439 5135 16445
rect 5077 16436 5089 16439
rect 4908 16408 5089 16436
rect 5077 16405 5089 16408
rect 5123 16436 5135 16439
rect 6454 16436 6460 16448
rect 5123 16408 6460 16436
rect 5123 16405 5135 16408
rect 5077 16399 5135 16405
rect 6454 16396 6460 16408
rect 6512 16396 6518 16448
rect 8757 16439 8815 16445
rect 8757 16405 8769 16439
rect 8803 16436 8815 16439
rect 8938 16436 8944 16448
rect 8803 16408 8944 16436
rect 8803 16405 8815 16408
rect 8757 16399 8815 16405
rect 8938 16396 8944 16408
rect 8996 16396 9002 16448
rect 15105 16439 15163 16445
rect 15105 16405 15117 16439
rect 15151 16436 15163 16439
rect 15194 16436 15200 16448
rect 15151 16408 15200 16436
rect 15151 16405 15163 16408
rect 15105 16399 15163 16405
rect 15194 16396 15200 16408
rect 15252 16396 15258 16448
rect 16206 16396 16212 16448
rect 16264 16396 16270 16448
rect 16758 16396 16764 16448
rect 16816 16436 16822 16448
rect 16945 16439 17003 16445
rect 16945 16436 16957 16439
rect 16816 16408 16957 16436
rect 16816 16396 16822 16408
rect 16945 16405 16957 16408
rect 16991 16405 17003 16439
rect 16945 16399 17003 16405
rect 19334 16396 19340 16448
rect 19392 16436 19398 16448
rect 19536 16445 19564 16544
rect 21076 16541 21088 16575
rect 21122 16572 21134 16575
rect 22186 16572 22192 16584
rect 21122 16544 22192 16572
rect 21122 16541 21134 16544
rect 21076 16535 21134 16541
rect 22186 16532 22192 16544
rect 22244 16532 22250 16584
rect 22278 16532 22284 16584
rect 22336 16532 22342 16584
rect 22548 16575 22606 16581
rect 22548 16541 22560 16575
rect 22594 16572 22606 16575
rect 23474 16572 23480 16584
rect 22594 16544 23480 16572
rect 22594 16541 22606 16544
rect 22548 16535 22606 16541
rect 23474 16532 23480 16544
rect 23532 16532 23538 16584
rect 24486 16532 24492 16584
rect 24544 16572 24550 16584
rect 24688 16581 24716 16612
rect 24673 16575 24731 16581
rect 24673 16572 24685 16575
rect 24544 16544 24685 16572
rect 24544 16532 24550 16544
rect 24673 16541 24685 16544
rect 24719 16541 24731 16575
rect 24673 16535 24731 16541
rect 25314 16532 25320 16584
rect 25372 16532 25378 16584
rect 25516 16581 25544 16612
rect 25590 16600 25596 16652
rect 25648 16640 25654 16652
rect 25700 16640 25728 16680
rect 26142 16668 26148 16680
rect 26200 16708 26206 16720
rect 27525 16711 27583 16717
rect 27525 16708 27537 16711
rect 26200 16680 27537 16708
rect 26200 16668 26206 16680
rect 27525 16677 27537 16680
rect 27571 16677 27583 16711
rect 27525 16671 27583 16677
rect 25648 16612 25728 16640
rect 25648 16600 25654 16612
rect 25700 16581 25728 16612
rect 26602 16600 26608 16652
rect 26660 16600 26666 16652
rect 28994 16600 29000 16652
rect 29052 16640 29058 16652
rect 29641 16643 29699 16649
rect 29641 16640 29653 16643
rect 29052 16612 29653 16640
rect 29052 16600 29058 16612
rect 29641 16609 29653 16612
rect 29687 16609 29699 16643
rect 30561 16643 30619 16649
rect 30561 16640 30573 16643
rect 29641 16603 29699 16609
rect 30300 16612 30573 16640
rect 25501 16575 25559 16581
rect 25501 16541 25513 16575
rect 25547 16541 25559 16575
rect 25501 16535 25559 16541
rect 25685 16575 25743 16581
rect 25685 16541 25697 16575
rect 25731 16541 25743 16575
rect 25685 16535 25743 16541
rect 26510 16532 26516 16584
rect 26568 16572 26574 16584
rect 26973 16575 27031 16581
rect 26973 16572 26985 16575
rect 26568 16544 26985 16572
rect 26568 16532 26574 16544
rect 26973 16541 26985 16544
rect 27019 16541 27031 16575
rect 26973 16535 27031 16541
rect 27249 16575 27307 16581
rect 27249 16541 27261 16575
rect 27295 16572 27307 16575
rect 27338 16572 27344 16584
rect 27295 16544 27344 16572
rect 27295 16541 27307 16544
rect 27249 16535 27307 16541
rect 27338 16532 27344 16544
rect 27396 16572 27402 16584
rect 28074 16572 28080 16584
rect 27396 16544 28080 16572
rect 27396 16532 27402 16544
rect 28074 16532 28080 16544
rect 28132 16532 28138 16584
rect 28629 16575 28687 16581
rect 28629 16541 28641 16575
rect 28675 16572 28687 16575
rect 28718 16572 28724 16584
rect 28675 16544 28724 16572
rect 28675 16541 28687 16544
rect 28629 16535 28687 16541
rect 28718 16532 28724 16544
rect 28776 16532 28782 16584
rect 28902 16532 28908 16584
rect 28960 16532 28966 16584
rect 29546 16532 29552 16584
rect 29604 16532 29610 16584
rect 30006 16532 30012 16584
rect 30064 16572 30070 16584
rect 30300 16572 30328 16612
rect 30561 16609 30573 16612
rect 30607 16609 30619 16643
rect 30561 16603 30619 16609
rect 31021 16643 31079 16649
rect 31021 16609 31033 16643
rect 31067 16640 31079 16643
rect 31478 16640 31484 16652
rect 31067 16612 31484 16640
rect 31067 16609 31079 16612
rect 31021 16603 31079 16609
rect 31478 16600 31484 16612
rect 31536 16600 31542 16652
rect 30064 16544 30328 16572
rect 30064 16532 30070 16544
rect 30374 16532 30380 16584
rect 30432 16572 30438 16584
rect 30742 16572 30748 16584
rect 30432 16544 30748 16572
rect 30432 16532 30438 16544
rect 30742 16532 30748 16544
rect 30800 16532 30806 16584
rect 32769 16575 32827 16581
rect 32769 16541 32781 16575
rect 32815 16572 32827 16575
rect 32858 16572 32864 16584
rect 32815 16544 32864 16572
rect 32815 16541 32827 16544
rect 32769 16535 32827 16541
rect 32858 16532 32864 16544
rect 32916 16532 32922 16584
rect 34054 16532 34060 16584
rect 34112 16532 34118 16584
rect 23382 16464 23388 16516
rect 23440 16504 23446 16516
rect 23934 16504 23940 16516
rect 23440 16476 23940 16504
rect 23440 16464 23446 16476
rect 23934 16464 23940 16476
rect 23992 16464 23998 16516
rect 25406 16504 25412 16516
rect 24504 16476 25412 16504
rect 19521 16439 19579 16445
rect 19521 16436 19533 16439
rect 19392 16408 19533 16436
rect 19392 16396 19398 16408
rect 19521 16405 19533 16408
rect 19567 16405 19579 16439
rect 19521 16399 19579 16405
rect 22094 16396 22100 16448
rect 22152 16436 22158 16448
rect 24504 16436 24532 16476
rect 25406 16464 25412 16476
rect 25464 16464 25470 16516
rect 25593 16507 25651 16513
rect 25593 16473 25605 16507
rect 25639 16473 25651 16507
rect 30926 16504 30932 16516
rect 25593 16467 25651 16473
rect 26528 16476 27476 16504
rect 22152 16408 24532 16436
rect 22152 16396 22158 16408
rect 24578 16396 24584 16448
rect 24636 16436 24642 16448
rect 25608 16436 25636 16467
rect 24636 16408 25636 16436
rect 24636 16396 24642 16408
rect 25866 16396 25872 16448
rect 25924 16396 25930 16448
rect 26050 16396 26056 16448
rect 26108 16396 26114 16448
rect 26418 16396 26424 16448
rect 26476 16396 26482 16448
rect 26528 16445 26556 16476
rect 27448 16448 27476 16476
rect 29932 16476 30932 16504
rect 26513 16439 26571 16445
rect 26513 16405 26525 16439
rect 26559 16405 26571 16439
rect 26513 16399 26571 16405
rect 27430 16396 27436 16448
rect 27488 16396 27494 16448
rect 28813 16439 28871 16445
rect 28813 16405 28825 16439
rect 28859 16436 28871 16439
rect 29086 16436 29092 16448
rect 28859 16408 29092 16436
rect 28859 16405 28871 16408
rect 28813 16399 28871 16405
rect 29086 16396 29092 16408
rect 29144 16396 29150 16448
rect 29270 16396 29276 16448
rect 29328 16396 29334 16448
rect 29932 16445 29960 16476
rect 30926 16464 30932 16476
rect 30984 16464 30990 16516
rect 33134 16504 33140 16516
rect 32246 16476 33140 16504
rect 33134 16464 33140 16476
rect 33192 16464 33198 16516
rect 34330 16464 34336 16516
rect 34388 16464 34394 16516
rect 29917 16439 29975 16445
rect 29917 16405 29929 16439
rect 29963 16405 29975 16439
rect 29917 16399 29975 16405
rect 31662 16396 31668 16448
rect 31720 16436 31726 16448
rect 32493 16439 32551 16445
rect 32493 16436 32505 16439
rect 31720 16408 32505 16436
rect 31720 16396 31726 16408
rect 32493 16405 32505 16408
rect 32539 16405 32551 16439
rect 32493 16399 32551 16405
rect 32582 16396 32588 16448
rect 32640 16396 32646 16448
rect 32950 16396 32956 16448
rect 33008 16396 33014 16448
rect 1104 16346 35328 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35328 16346
rect 1104 16272 35328 16294
rect 3605 16235 3663 16241
rect 3605 16201 3617 16235
rect 3651 16232 3663 16235
rect 3651 16204 3740 16232
rect 3651 16201 3663 16204
rect 3605 16195 3663 16201
rect 3712 16164 3740 16204
rect 4062 16192 4068 16244
rect 4120 16192 4126 16244
rect 4433 16235 4491 16241
rect 4433 16201 4445 16235
rect 4479 16232 4491 16235
rect 4614 16232 4620 16244
rect 4479 16204 4620 16232
rect 4479 16201 4491 16204
rect 4433 16195 4491 16201
rect 4614 16192 4620 16204
rect 4672 16192 4678 16244
rect 8018 16192 8024 16244
rect 8076 16192 8082 16244
rect 8481 16235 8539 16241
rect 8481 16232 8493 16235
rect 8128 16204 8493 16232
rect 8128 16164 8156 16204
rect 8481 16201 8493 16204
rect 8527 16232 8539 16235
rect 11146 16232 11152 16244
rect 8527 16204 11152 16232
rect 8527 16201 8539 16204
rect 8481 16195 8539 16201
rect 11146 16192 11152 16204
rect 11204 16192 11210 16244
rect 11790 16192 11796 16244
rect 11848 16192 11854 16244
rect 12250 16192 12256 16244
rect 12308 16192 12314 16244
rect 12710 16192 12716 16244
rect 12768 16192 12774 16244
rect 14553 16235 14611 16241
rect 14553 16201 14565 16235
rect 14599 16201 14611 16235
rect 14553 16195 14611 16201
rect 3712 16136 8156 16164
rect 8389 16167 8447 16173
rect 1578 16056 1584 16108
rect 1636 16096 1642 16108
rect 3712 16105 3740 16136
rect 8389 16133 8401 16167
rect 8435 16164 8447 16167
rect 12161 16167 12219 16173
rect 12161 16164 12173 16167
rect 8435 16136 8984 16164
rect 8435 16133 8447 16136
rect 8389 16127 8447 16133
rect 8956 16108 8984 16136
rect 10888 16136 12173 16164
rect 10888 16108 10916 16136
rect 12161 16133 12173 16136
rect 12207 16133 12219 16167
rect 13348 16167 13406 16173
rect 12161 16127 12219 16133
rect 12406 16136 13308 16164
rect 3421 16099 3479 16105
rect 3421 16096 3433 16099
rect 1636 16068 3433 16096
rect 1636 16056 1642 16068
rect 3421 16065 3433 16068
rect 3467 16065 3479 16099
rect 3421 16059 3479 16065
rect 3697 16099 3755 16105
rect 3697 16065 3709 16099
rect 3743 16065 3755 16099
rect 3697 16059 3755 16065
rect 5350 16056 5356 16108
rect 5408 16096 5414 16108
rect 6638 16105 6644 16108
rect 6365 16099 6423 16105
rect 6365 16096 6377 16099
rect 5408 16068 6377 16096
rect 5408 16056 5414 16068
rect 6365 16065 6377 16068
rect 6411 16065 6423 16099
rect 6365 16059 6423 16065
rect 6632 16059 6644 16105
rect 6638 16056 6644 16059
rect 6696 16056 6702 16108
rect 7558 16056 7564 16108
rect 7616 16096 7622 16108
rect 8849 16099 8907 16105
rect 8849 16096 8861 16099
rect 7616 16068 8861 16096
rect 7616 16056 7622 16068
rect 8849 16065 8861 16068
rect 8895 16065 8907 16099
rect 8849 16059 8907 16065
rect 8938 16056 8944 16108
rect 8996 16096 9002 16108
rect 9125 16099 9183 16105
rect 8996 16068 9041 16096
rect 8996 16056 9002 16068
rect 9125 16065 9137 16099
rect 9171 16065 9183 16099
rect 9125 16059 9183 16065
rect 4525 16031 4583 16037
rect 4525 15997 4537 16031
rect 4571 15997 4583 16031
rect 4525 15991 4583 15997
rect 3881 15895 3939 15901
rect 3881 15861 3893 15895
rect 3927 15892 3939 15895
rect 4062 15892 4068 15904
rect 3927 15864 4068 15892
rect 3927 15861 3939 15864
rect 3881 15855 3939 15861
rect 4062 15852 4068 15864
rect 4120 15892 4126 15904
rect 4540 15892 4568 15991
rect 4706 15988 4712 16040
rect 4764 15988 4770 16040
rect 8665 16031 8723 16037
rect 8665 15997 8677 16031
rect 8711 16028 8723 16031
rect 9030 16028 9036 16040
rect 8711 16000 9036 16028
rect 8711 15997 8723 16000
rect 8665 15991 8723 15997
rect 9030 15988 9036 16000
rect 9088 15988 9094 16040
rect 9140 16028 9168 16059
rect 9214 16056 9220 16108
rect 9272 16056 9278 16108
rect 9398 16105 9404 16108
rect 9355 16099 9404 16105
rect 9355 16065 9367 16099
rect 9401 16065 9404 16099
rect 9355 16059 9404 16065
rect 9398 16056 9404 16059
rect 9456 16096 9462 16108
rect 9769 16099 9827 16105
rect 9769 16096 9781 16099
rect 9456 16068 9781 16096
rect 9456 16056 9462 16068
rect 9769 16065 9781 16068
rect 9815 16065 9827 16099
rect 9769 16059 9827 16065
rect 10870 16056 10876 16108
rect 10928 16056 10934 16108
rect 11146 16056 11152 16108
rect 11204 16056 11210 16108
rect 12406 16096 12434 16136
rect 11624 16068 12434 16096
rect 9140 16000 9260 16028
rect 6730 15892 6736 15904
rect 4120 15864 6736 15892
rect 4120 15852 4126 15864
rect 6730 15852 6736 15864
rect 6788 15852 6794 15904
rect 7742 15852 7748 15904
rect 7800 15852 7806 15904
rect 9232 15892 9260 16000
rect 9493 15963 9551 15969
rect 9493 15929 9505 15963
rect 9539 15960 9551 15963
rect 11330 15960 11336 15972
rect 9539 15932 11336 15960
rect 9539 15929 9551 15932
rect 9493 15923 9551 15929
rect 11330 15920 11336 15932
rect 11388 15920 11394 15972
rect 9677 15895 9735 15901
rect 9677 15892 9689 15895
rect 9232 15864 9689 15892
rect 9677 15861 9689 15864
rect 9723 15892 9735 15895
rect 9766 15892 9772 15904
rect 9723 15864 9772 15892
rect 9723 15861 9735 15864
rect 9677 15855 9735 15861
rect 9766 15852 9772 15864
rect 9824 15892 9830 15904
rect 11624 15892 11652 16068
rect 13078 16056 13084 16108
rect 13136 16056 13142 16108
rect 13280 16096 13308 16136
rect 13348 16133 13360 16167
rect 13394 16164 13406 16167
rect 14568 16164 14596 16195
rect 15102 16192 15108 16244
rect 15160 16232 15166 16244
rect 15381 16235 15439 16241
rect 15381 16232 15393 16235
rect 15160 16204 15393 16232
rect 15160 16192 15166 16204
rect 15381 16201 15393 16204
rect 15427 16201 15439 16235
rect 15381 16195 15439 16201
rect 15654 16192 15660 16244
rect 15712 16232 15718 16244
rect 16114 16232 16120 16244
rect 15712 16204 16120 16232
rect 15712 16192 15718 16204
rect 16114 16192 16120 16204
rect 16172 16232 16178 16244
rect 16301 16235 16359 16241
rect 16301 16232 16313 16235
rect 16172 16204 16313 16232
rect 16172 16192 16178 16204
rect 16301 16201 16313 16204
rect 16347 16201 16359 16235
rect 16301 16195 16359 16201
rect 17589 16235 17647 16241
rect 17589 16201 17601 16235
rect 17635 16232 17647 16235
rect 17954 16232 17960 16244
rect 17635 16204 17960 16232
rect 17635 16201 17647 16204
rect 17589 16195 17647 16201
rect 17954 16192 17960 16204
rect 18012 16192 18018 16244
rect 22094 16232 22100 16244
rect 18892 16204 22100 16232
rect 13394 16136 14596 16164
rect 15672 16164 15700 16192
rect 15841 16167 15899 16173
rect 15841 16164 15853 16167
rect 15672 16136 15853 16164
rect 13394 16133 13406 16136
rect 13348 16127 13406 16133
rect 15841 16133 15853 16136
rect 15887 16133 15899 16167
rect 15841 16127 15899 16133
rect 15930 16124 15936 16176
rect 15988 16124 15994 16176
rect 18892 16173 18920 16204
rect 22094 16192 22100 16204
rect 22152 16192 22158 16244
rect 22370 16232 22376 16244
rect 22204 16204 22376 16232
rect 18877 16167 18935 16173
rect 18877 16133 18889 16167
rect 18923 16133 18935 16167
rect 22204 16164 22232 16204
rect 22370 16192 22376 16204
rect 22428 16192 22434 16244
rect 22462 16192 22468 16244
rect 22520 16232 22526 16244
rect 23017 16235 23075 16241
rect 23017 16232 23029 16235
rect 22520 16204 23029 16232
rect 22520 16192 22526 16204
rect 23017 16201 23029 16204
rect 23063 16201 23075 16235
rect 23017 16195 23075 16201
rect 25406 16192 25412 16244
rect 25464 16232 25470 16244
rect 27617 16235 27675 16241
rect 25464 16204 27568 16232
rect 25464 16192 25470 16204
rect 18877 16127 18935 16133
rect 21928 16136 22232 16164
rect 13722 16096 13728 16108
rect 13280 16068 13728 16096
rect 13722 16056 13728 16068
rect 13780 16096 13786 16108
rect 14090 16096 14096 16108
rect 13780 16068 14096 16096
rect 13780 16056 13786 16068
rect 14090 16056 14096 16068
rect 14148 16056 14154 16108
rect 14550 16096 14556 16108
rect 14476 16068 14556 16096
rect 12437 16031 12495 16037
rect 12437 15997 12449 16031
rect 12483 16028 12495 16031
rect 12710 16028 12716 16040
rect 12483 16000 12716 16028
rect 12483 15997 12495 16000
rect 12437 15991 12495 15997
rect 12710 15988 12716 16000
rect 12768 15988 12774 16040
rect 14476 15969 14504 16068
rect 14550 16056 14556 16068
rect 14608 16096 14614 16108
rect 14921 16099 14979 16105
rect 14921 16096 14933 16099
rect 14608 16068 14933 16096
rect 14608 16056 14614 16068
rect 14921 16065 14933 16068
rect 14967 16065 14979 16099
rect 14921 16059 14979 16065
rect 15194 16056 15200 16108
rect 15252 16096 15258 16108
rect 15565 16099 15623 16105
rect 15565 16096 15577 16099
rect 15252 16068 15577 16096
rect 15252 16056 15258 16068
rect 15565 16065 15577 16068
rect 15611 16065 15623 16099
rect 15565 16059 15623 16065
rect 15654 16056 15660 16108
rect 15712 16056 15718 16108
rect 16030 16099 16088 16105
rect 16030 16096 16042 16099
rect 15764 16068 16042 16096
rect 15010 15988 15016 16040
rect 15068 15988 15074 16040
rect 15102 15988 15108 16040
rect 15160 15988 15166 16040
rect 15378 15988 15384 16040
rect 15436 16028 15442 16040
rect 15764 16028 15792 16068
rect 16030 16065 16042 16068
rect 16076 16096 16088 16099
rect 16669 16099 16727 16105
rect 16669 16096 16681 16099
rect 16076 16068 16681 16096
rect 16076 16065 16088 16068
rect 16030 16059 16088 16065
rect 16669 16065 16681 16068
rect 16715 16096 16727 16099
rect 16758 16096 16764 16108
rect 16715 16068 16764 16096
rect 16715 16065 16727 16068
rect 16669 16059 16727 16065
rect 16758 16056 16764 16068
rect 16816 16056 16822 16108
rect 17313 16099 17371 16105
rect 17313 16065 17325 16099
rect 17359 16096 17371 16099
rect 17494 16096 17500 16108
rect 17359 16068 17500 16096
rect 17359 16065 17371 16068
rect 17313 16059 17371 16065
rect 17494 16056 17500 16068
rect 17552 16056 17558 16108
rect 18782 16105 18788 16108
rect 18601 16099 18659 16105
rect 18601 16065 18613 16099
rect 18647 16065 18659 16099
rect 18601 16059 18659 16065
rect 18749 16099 18788 16105
rect 18749 16065 18761 16099
rect 18749 16059 18788 16065
rect 15436 16000 15792 16028
rect 18616 16028 18644 16059
rect 18782 16056 18788 16059
rect 18840 16056 18846 16108
rect 18966 16056 18972 16108
rect 19024 16056 19030 16108
rect 19107 16099 19165 16105
rect 19107 16065 19119 16099
rect 19153 16096 19165 16099
rect 19242 16096 19248 16108
rect 19153 16068 19248 16096
rect 19153 16065 19165 16068
rect 19107 16059 19165 16065
rect 19242 16056 19248 16068
rect 19300 16056 19306 16108
rect 19788 16099 19846 16105
rect 19788 16065 19800 16099
rect 19834 16096 19846 16099
rect 20070 16096 20076 16108
rect 19834 16068 20076 16096
rect 19834 16065 19846 16068
rect 19788 16059 19846 16065
rect 20070 16056 20076 16068
rect 20128 16056 20134 16108
rect 21450 16056 21456 16108
rect 21508 16096 21514 16108
rect 21928 16105 21956 16136
rect 22278 16124 22284 16176
rect 22336 16164 22342 16176
rect 24670 16164 24676 16176
rect 22336 16136 24676 16164
rect 22336 16124 22342 16136
rect 21821 16099 21879 16105
rect 21821 16096 21833 16099
rect 21508 16068 21833 16096
rect 21508 16056 21514 16068
rect 21821 16065 21833 16068
rect 21867 16065 21879 16099
rect 21821 16059 21879 16065
rect 21913 16099 21971 16105
rect 21913 16065 21925 16099
rect 21959 16065 21971 16099
rect 21913 16059 21971 16065
rect 22097 16099 22155 16105
rect 22097 16065 22109 16099
rect 22143 16065 22155 16099
rect 22097 16059 22155 16065
rect 19334 16028 19340 16040
rect 18616 16000 19340 16028
rect 15436 15988 15442 16000
rect 19334 15988 19340 16000
rect 19392 15988 19398 16040
rect 19426 15988 19432 16040
rect 19484 16028 19490 16040
rect 19521 16031 19579 16037
rect 19521 16028 19533 16031
rect 19484 16000 19533 16028
rect 19484 15988 19490 16000
rect 19521 15997 19533 16000
rect 19567 15997 19579 16031
rect 22112 16028 22140 16059
rect 22186 16056 22192 16108
rect 22244 16096 22250 16108
rect 22462 16096 22468 16108
rect 22244 16068 22468 16096
rect 22244 16056 22250 16068
rect 22462 16056 22468 16068
rect 22520 16056 22526 16108
rect 22649 16099 22707 16105
rect 22649 16065 22661 16099
rect 22695 16096 22707 16099
rect 22922 16096 22928 16108
rect 22695 16068 22928 16096
rect 22695 16065 22707 16068
rect 22649 16059 22707 16065
rect 22922 16056 22928 16068
rect 22980 16056 22986 16108
rect 23308 16105 23336 16136
rect 24670 16124 24676 16136
rect 24728 16124 24734 16176
rect 24762 16124 24768 16176
rect 24820 16164 24826 16176
rect 24857 16167 24915 16173
rect 24857 16164 24869 16167
rect 24820 16136 24869 16164
rect 24820 16124 24826 16136
rect 24857 16133 24869 16136
rect 24903 16164 24915 16167
rect 24949 16167 25007 16173
rect 24949 16164 24961 16167
rect 24903 16136 24961 16164
rect 24903 16133 24915 16136
rect 24857 16127 24915 16133
rect 24949 16133 24961 16136
rect 24995 16133 25007 16167
rect 24949 16127 25007 16133
rect 25866 16124 25872 16176
rect 25924 16164 25930 16176
rect 25924 16136 26832 16164
rect 25924 16124 25930 16136
rect 23293 16099 23351 16105
rect 23293 16065 23305 16099
rect 23339 16065 23351 16099
rect 23293 16059 23351 16065
rect 23560 16099 23618 16105
rect 23560 16065 23572 16099
rect 23606 16096 23618 16099
rect 24302 16096 24308 16108
rect 23606 16068 24308 16096
rect 23606 16065 23618 16068
rect 23560 16059 23618 16065
rect 24302 16056 24308 16068
rect 24360 16056 24366 16108
rect 25314 16056 25320 16108
rect 25372 16096 25378 16108
rect 26326 16096 26332 16108
rect 25372 16068 26332 16096
rect 25372 16056 25378 16068
rect 26326 16056 26332 16068
rect 26384 16096 26390 16108
rect 26513 16099 26571 16105
rect 26513 16096 26525 16099
rect 26384 16068 26525 16096
rect 26384 16056 26390 16068
rect 26513 16065 26525 16068
rect 26559 16065 26571 16099
rect 26804 16096 26832 16136
rect 26878 16124 26884 16176
rect 26936 16164 26942 16176
rect 27249 16167 27307 16173
rect 27249 16164 27261 16167
rect 26936 16136 27261 16164
rect 26936 16124 26942 16136
rect 27249 16133 27261 16136
rect 27295 16133 27307 16167
rect 27540 16164 27568 16204
rect 27617 16201 27629 16235
rect 27663 16232 27675 16235
rect 29546 16232 29552 16244
rect 27663 16204 29552 16232
rect 27663 16201 27675 16204
rect 27617 16195 27675 16201
rect 29546 16192 29552 16204
rect 29604 16192 29610 16244
rect 28902 16164 28908 16176
rect 27540 16136 28908 16164
rect 27249 16127 27307 16133
rect 28902 16124 28908 16136
rect 28960 16124 28966 16176
rect 29270 16124 29276 16176
rect 29328 16164 29334 16176
rect 31202 16164 31208 16176
rect 29328 16136 31208 16164
rect 29328 16124 29334 16136
rect 31202 16124 31208 16136
rect 31260 16124 31266 16176
rect 33134 16124 33140 16176
rect 33192 16124 33198 16176
rect 26973 16099 27031 16105
rect 26973 16096 26985 16099
rect 26804 16068 26985 16096
rect 26513 16059 26571 16065
rect 26973 16065 26985 16068
rect 27019 16065 27031 16099
rect 26973 16059 27031 16065
rect 27062 16056 27068 16108
rect 27120 16056 27126 16108
rect 27341 16099 27399 16105
rect 27341 16065 27353 16099
rect 27387 16065 27399 16099
rect 27341 16059 27399 16065
rect 27438 16099 27496 16105
rect 27438 16065 27450 16099
rect 27484 16065 27496 16099
rect 27438 16059 27496 16065
rect 28068 16099 28126 16105
rect 28068 16065 28080 16099
rect 28114 16096 28126 16099
rect 28442 16096 28448 16108
rect 28114 16068 28448 16096
rect 28114 16065 28126 16068
rect 28068 16059 28126 16065
rect 22554 16028 22560 16040
rect 22112 16000 22560 16028
rect 19521 15991 19579 15997
rect 22554 15988 22560 16000
rect 22612 15988 22618 16040
rect 26418 15988 26424 16040
rect 26476 16028 26482 16040
rect 27356 16028 27384 16059
rect 26476 16000 27384 16028
rect 26476 15988 26482 16000
rect 14461 15963 14519 15969
rect 14461 15929 14473 15963
rect 14507 15929 14519 15963
rect 14461 15923 14519 15929
rect 19245 15963 19303 15969
rect 19245 15929 19257 15963
rect 19291 15960 19303 15963
rect 22373 15963 22431 15969
rect 19291 15932 19564 15960
rect 19291 15929 19303 15932
rect 19245 15923 19303 15929
rect 19536 15904 19564 15932
rect 22373 15929 22385 15963
rect 22419 15960 22431 15963
rect 22419 15932 23336 15960
rect 22419 15929 22431 15932
rect 22373 15923 22431 15929
rect 9824 15864 11652 15892
rect 9824 15852 9830 15864
rect 11698 15852 11704 15904
rect 11756 15892 11762 15904
rect 14274 15892 14280 15904
rect 11756 15864 14280 15892
rect 11756 15852 11762 15864
rect 14274 15852 14280 15864
rect 14332 15852 14338 15904
rect 15838 15852 15844 15904
rect 15896 15892 15902 15904
rect 16209 15895 16267 15901
rect 16209 15892 16221 15895
rect 15896 15864 16221 15892
rect 15896 15852 15902 15864
rect 16209 15861 16221 15864
rect 16255 15861 16267 15895
rect 16209 15855 16267 15861
rect 19334 15852 19340 15904
rect 19392 15852 19398 15904
rect 19518 15852 19524 15904
rect 19576 15852 19582 15904
rect 20714 15852 20720 15904
rect 20772 15892 20778 15904
rect 20901 15895 20959 15901
rect 20901 15892 20913 15895
rect 20772 15864 20913 15892
rect 20772 15852 20778 15864
rect 20901 15861 20913 15864
rect 20947 15861 20959 15895
rect 20901 15855 20959 15861
rect 22925 15895 22983 15901
rect 22925 15861 22937 15895
rect 22971 15892 22983 15895
rect 23106 15892 23112 15904
rect 22971 15864 23112 15892
rect 22971 15861 22983 15864
rect 22925 15855 22983 15861
rect 23106 15852 23112 15864
rect 23164 15852 23170 15904
rect 23308 15892 23336 15932
rect 24578 15920 24584 15972
rect 24636 15960 24642 15972
rect 24673 15963 24731 15969
rect 24673 15960 24685 15963
rect 24636 15932 24685 15960
rect 24636 15920 24642 15932
rect 24673 15929 24685 15932
rect 24719 15929 24731 15963
rect 24673 15923 24731 15929
rect 25774 15920 25780 15972
rect 25832 15960 25838 15972
rect 27246 15960 27252 15972
rect 25832 15932 27252 15960
rect 25832 15920 25838 15932
rect 27246 15920 27252 15932
rect 27304 15960 27310 15972
rect 27448 15960 27476 16059
rect 28442 16056 28448 16068
rect 28500 16056 28506 16108
rect 30834 16056 30840 16108
rect 30892 16096 30898 16108
rect 30929 16099 30987 16105
rect 30929 16096 30941 16099
rect 30892 16068 30941 16096
rect 30892 16056 30898 16068
rect 30929 16065 30941 16068
rect 30975 16065 30987 16099
rect 30929 16059 30987 16065
rect 31021 16099 31079 16105
rect 31021 16065 31033 16099
rect 31067 16096 31079 16099
rect 31386 16096 31392 16108
rect 31067 16068 31392 16096
rect 31067 16065 31079 16068
rect 31021 16059 31079 16065
rect 31386 16056 31392 16068
rect 31444 16056 31450 16108
rect 31605 16099 31663 16105
rect 31605 16096 31617 16099
rect 31588 16065 31617 16096
rect 31651 16065 31663 16099
rect 31588 16059 31663 16065
rect 27798 15988 27804 16040
rect 27856 15988 27862 16040
rect 30101 16031 30159 16037
rect 30101 15997 30113 16031
rect 30147 16028 30159 16031
rect 30374 16028 30380 16040
rect 30147 16000 30380 16028
rect 30147 15997 30159 16000
rect 30101 15991 30159 15997
rect 30374 15988 30380 16000
rect 30432 15988 30438 16040
rect 30469 16031 30527 16037
rect 30469 15997 30481 16031
rect 30515 16028 30527 16031
rect 30558 16028 30564 16040
rect 30515 16000 30564 16028
rect 30515 15997 30527 16000
rect 30469 15991 30527 15997
rect 30558 15988 30564 16000
rect 30616 16028 30622 16040
rect 31110 16028 31116 16040
rect 30616 16000 31116 16028
rect 30616 15988 30622 16000
rect 31110 15988 31116 16000
rect 31168 15988 31174 16040
rect 27304 15932 27476 15960
rect 27304 15920 27310 15932
rect 29086 15920 29092 15972
rect 29144 15960 29150 15972
rect 29454 15960 29460 15972
rect 29144 15932 29460 15960
rect 29144 15920 29150 15932
rect 29454 15920 29460 15932
rect 29512 15960 29518 15972
rect 31588 15960 31616 16059
rect 32122 15988 32128 16040
rect 32180 16028 32186 16040
rect 32401 16031 32459 16037
rect 32401 16028 32413 16031
rect 32180 16000 32413 16028
rect 32180 15988 32186 16000
rect 32401 15997 32413 16000
rect 32447 15997 32459 16031
rect 32401 15991 32459 15997
rect 32674 15988 32680 16040
rect 32732 15988 32738 16040
rect 29512 15932 31984 15960
rect 29512 15920 29518 15932
rect 31956 15904 31984 15932
rect 28994 15892 29000 15904
rect 23308 15864 29000 15892
rect 28994 15852 29000 15864
rect 29052 15852 29058 15904
rect 29178 15852 29184 15904
rect 29236 15852 29242 15904
rect 30561 15895 30619 15901
rect 30561 15861 30573 15895
rect 30607 15892 30619 15895
rect 30650 15892 30656 15904
rect 30607 15864 30656 15892
rect 30607 15861 30619 15864
rect 30561 15855 30619 15861
rect 30650 15852 30656 15864
rect 30708 15852 30714 15904
rect 31478 15852 31484 15904
rect 31536 15852 31542 15904
rect 31846 15852 31852 15904
rect 31904 15852 31910 15904
rect 31938 15852 31944 15904
rect 31996 15892 32002 15904
rect 32125 15895 32183 15901
rect 32125 15892 32137 15895
rect 31996 15864 32137 15892
rect 31996 15852 32002 15864
rect 32125 15861 32137 15864
rect 32171 15861 32183 15895
rect 32125 15855 32183 15861
rect 33410 15852 33416 15904
rect 33468 15892 33474 15904
rect 34054 15892 34060 15904
rect 33468 15864 34060 15892
rect 33468 15852 33474 15864
rect 34054 15852 34060 15864
rect 34112 15892 34118 15904
rect 34149 15895 34207 15901
rect 34149 15892 34161 15895
rect 34112 15864 34161 15892
rect 34112 15852 34118 15864
rect 34149 15861 34161 15864
rect 34195 15861 34207 15895
rect 34149 15855 34207 15861
rect 1104 15802 35328 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 35328 15802
rect 1104 15728 35328 15750
rect 6638 15648 6644 15700
rect 6696 15688 6702 15700
rect 6825 15691 6883 15697
rect 6825 15688 6837 15691
rect 6696 15660 6837 15688
rect 6696 15648 6702 15660
rect 6825 15657 6837 15660
rect 6871 15657 6883 15691
rect 6825 15651 6883 15657
rect 7558 15648 7564 15700
rect 7616 15648 7622 15700
rect 7650 15648 7656 15700
rect 7708 15648 7714 15700
rect 8110 15648 8116 15700
rect 8168 15688 8174 15700
rect 12894 15688 12900 15700
rect 8168 15660 12900 15688
rect 8168 15648 8174 15660
rect 5813 15623 5871 15629
rect 5813 15589 5825 15623
rect 5859 15620 5871 15623
rect 5859 15592 8432 15620
rect 5859 15589 5871 15592
rect 5813 15583 5871 15589
rect 5442 15512 5448 15564
rect 5500 15552 5506 15564
rect 5500 15524 5672 15552
rect 5500 15512 5506 15524
rect 2225 15487 2283 15493
rect 2225 15453 2237 15487
rect 2271 15484 2283 15487
rect 2774 15484 2780 15496
rect 2271 15456 2780 15484
rect 2271 15453 2283 15456
rect 2225 15447 2283 15453
rect 2774 15444 2780 15456
rect 2832 15484 2838 15496
rect 3789 15487 3847 15493
rect 3789 15484 3801 15487
rect 2832 15456 3801 15484
rect 2832 15444 2838 15456
rect 3789 15453 3801 15456
rect 3835 15453 3847 15487
rect 5261 15487 5319 15493
rect 5261 15484 5273 15487
rect 3789 15447 3847 15453
rect 3988 15456 5273 15484
rect 2492 15419 2550 15425
rect 2492 15385 2504 15419
rect 2538 15416 2550 15419
rect 2866 15416 2872 15428
rect 2538 15388 2872 15416
rect 2538 15385 2550 15388
rect 2492 15379 2550 15385
rect 2866 15376 2872 15388
rect 2924 15376 2930 15428
rect 3234 15308 3240 15360
rect 3292 15348 3298 15360
rect 3605 15351 3663 15357
rect 3605 15348 3617 15351
rect 3292 15320 3617 15348
rect 3292 15308 3298 15320
rect 3605 15317 3617 15320
rect 3651 15348 3663 15351
rect 3988 15348 4016 15456
rect 5261 15453 5273 15456
rect 5307 15453 5319 15487
rect 5261 15447 5319 15453
rect 5534 15444 5540 15496
rect 5592 15444 5598 15496
rect 5644 15493 5672 15524
rect 6270 15512 6276 15564
rect 6328 15512 6334 15564
rect 7193 15555 7251 15561
rect 7193 15552 7205 15555
rect 6472 15524 7205 15552
rect 5629 15487 5687 15493
rect 5629 15453 5641 15487
rect 5675 15453 5687 15487
rect 5629 15447 5687 15453
rect 4056 15419 4114 15425
rect 4056 15385 4068 15419
rect 4102 15416 4114 15419
rect 4154 15416 4160 15428
rect 4102 15388 4160 15416
rect 4102 15385 4114 15388
rect 4056 15379 4114 15385
rect 4154 15376 4160 15388
rect 4212 15376 4218 15428
rect 5350 15376 5356 15428
rect 5408 15416 5414 15428
rect 5445 15419 5503 15425
rect 5445 15416 5457 15419
rect 5408 15388 5457 15416
rect 5408 15376 5414 15388
rect 5445 15385 5457 15388
rect 5491 15416 5503 15419
rect 5905 15419 5963 15425
rect 5905 15416 5917 15419
rect 5491 15388 5917 15416
rect 5491 15385 5503 15388
rect 5445 15379 5503 15385
rect 5644 15360 5672 15388
rect 5905 15385 5917 15388
rect 5951 15385 5963 15419
rect 5905 15379 5963 15385
rect 3651 15320 4016 15348
rect 3651 15317 3663 15320
rect 3605 15311 3663 15317
rect 4614 15308 4620 15360
rect 4672 15348 4678 15360
rect 5169 15351 5227 15357
rect 5169 15348 5181 15351
rect 4672 15320 5181 15348
rect 4672 15308 4678 15320
rect 5169 15317 5181 15320
rect 5215 15348 5227 15351
rect 5534 15348 5540 15360
rect 5215 15320 5540 15348
rect 5215 15317 5227 15320
rect 5169 15311 5227 15317
rect 5534 15308 5540 15320
rect 5592 15308 5598 15360
rect 5626 15308 5632 15360
rect 5684 15308 5690 15360
rect 6288 15348 6316 15512
rect 6472 15493 6500 15524
rect 7193 15521 7205 15524
rect 7239 15552 7251 15555
rect 7742 15552 7748 15564
rect 7239 15524 7748 15552
rect 7239 15521 7251 15524
rect 7193 15515 7251 15521
rect 7742 15512 7748 15524
rect 7800 15512 7806 15564
rect 6457 15487 6515 15493
rect 6457 15453 6469 15487
rect 6503 15453 6515 15487
rect 6457 15447 6515 15453
rect 7377 15487 7435 15493
rect 7377 15453 7389 15487
rect 7423 15484 7435 15487
rect 7650 15484 7656 15496
rect 7423 15456 7656 15484
rect 7423 15453 7435 15456
rect 7377 15447 7435 15453
rect 7650 15444 7656 15456
rect 7708 15444 7714 15496
rect 8404 15484 8432 15592
rect 8573 15555 8631 15561
rect 8573 15521 8585 15555
rect 8619 15552 8631 15555
rect 9122 15552 9128 15564
rect 8619 15524 9128 15552
rect 8619 15521 8631 15524
rect 8573 15515 8631 15521
rect 9122 15512 9128 15524
rect 9180 15512 9186 15564
rect 9306 15512 9312 15564
rect 9364 15552 9370 15564
rect 9401 15555 9459 15561
rect 9401 15552 9413 15555
rect 9364 15524 9413 15552
rect 9364 15512 9370 15524
rect 9401 15521 9413 15524
rect 9447 15521 9459 15555
rect 9401 15515 9459 15521
rect 10873 15487 10931 15493
rect 10873 15484 10885 15487
rect 8404 15456 10885 15484
rect 10873 15453 10885 15456
rect 10919 15453 10931 15487
rect 10873 15447 10931 15453
rect 10966 15487 11024 15493
rect 10966 15453 10978 15487
rect 11012 15453 11024 15487
rect 11072 15484 11100 15660
rect 12894 15648 12900 15660
rect 12952 15688 12958 15700
rect 18877 15691 18935 15697
rect 12952 15660 18460 15688
rect 12952 15648 12958 15660
rect 15102 15580 15108 15632
rect 15160 15620 15166 15632
rect 15381 15623 15439 15629
rect 15381 15620 15393 15623
rect 15160 15592 15393 15620
rect 15160 15580 15166 15592
rect 15381 15589 15393 15592
rect 15427 15620 15439 15623
rect 16482 15620 16488 15632
rect 15427 15592 16488 15620
rect 15427 15589 15439 15592
rect 15381 15583 15439 15589
rect 16482 15580 16488 15592
rect 16540 15580 16546 15632
rect 18432 15620 18460 15660
rect 18877 15657 18889 15691
rect 18923 15688 18935 15691
rect 18966 15688 18972 15700
rect 18923 15660 18972 15688
rect 18923 15657 18935 15660
rect 18877 15651 18935 15657
rect 18966 15648 18972 15660
rect 19024 15648 19030 15700
rect 20070 15648 20076 15700
rect 20128 15648 20134 15700
rect 22554 15648 22560 15700
rect 22612 15688 22618 15700
rect 22649 15691 22707 15697
rect 22649 15688 22661 15691
rect 22612 15660 22661 15688
rect 22612 15648 22618 15660
rect 22649 15657 22661 15660
rect 22695 15657 22707 15691
rect 22649 15651 22707 15657
rect 23566 15648 23572 15700
rect 23624 15688 23630 15700
rect 23845 15691 23903 15697
rect 23845 15688 23857 15691
rect 23624 15660 23857 15688
rect 23624 15648 23630 15660
rect 23845 15657 23857 15660
rect 23891 15688 23903 15691
rect 24118 15688 24124 15700
rect 23891 15660 24124 15688
rect 23891 15657 23903 15660
rect 23845 15651 23903 15657
rect 24118 15648 24124 15660
rect 24176 15648 24182 15700
rect 24210 15648 24216 15700
rect 24268 15688 24274 15700
rect 24397 15691 24455 15697
rect 24397 15688 24409 15691
rect 24268 15660 24409 15688
rect 24268 15648 24274 15660
rect 24397 15657 24409 15660
rect 24443 15688 24455 15691
rect 24673 15691 24731 15697
rect 24673 15688 24685 15691
rect 24443 15660 24685 15688
rect 24443 15657 24455 15660
rect 24397 15651 24455 15657
rect 24673 15657 24685 15660
rect 24719 15657 24731 15691
rect 24673 15651 24731 15657
rect 26418 15648 26424 15700
rect 26476 15688 26482 15700
rect 26789 15691 26847 15697
rect 26789 15688 26801 15691
rect 26476 15660 26801 15688
rect 26476 15648 26482 15660
rect 26789 15657 26801 15660
rect 26835 15657 26847 15691
rect 26789 15651 26847 15657
rect 26878 15648 26884 15700
rect 26936 15648 26942 15700
rect 28442 15648 28448 15700
rect 28500 15648 28506 15700
rect 30190 15648 30196 15700
rect 30248 15648 30254 15700
rect 31386 15648 31392 15700
rect 31444 15688 31450 15700
rect 31757 15691 31815 15697
rect 31757 15688 31769 15691
rect 31444 15660 31769 15688
rect 31444 15648 31450 15660
rect 31757 15657 31769 15660
rect 31803 15657 31815 15691
rect 31757 15651 31815 15657
rect 19334 15620 19340 15632
rect 18432 15592 19340 15620
rect 19334 15580 19340 15592
rect 19392 15620 19398 15632
rect 19429 15623 19487 15629
rect 19429 15620 19441 15623
rect 19392 15592 19441 15620
rect 19392 15580 19398 15592
rect 19429 15589 19441 15592
rect 19475 15620 19487 15623
rect 19613 15623 19671 15629
rect 19613 15620 19625 15623
rect 19475 15592 19625 15620
rect 19475 15589 19487 15592
rect 19429 15583 19487 15589
rect 19613 15589 19625 15592
rect 19659 15589 19671 15623
rect 19613 15583 19671 15589
rect 22462 15580 22468 15632
rect 22520 15620 22526 15632
rect 22833 15623 22891 15629
rect 22833 15620 22845 15623
rect 22520 15592 22845 15620
rect 22520 15580 22526 15592
rect 22833 15589 22845 15592
rect 22879 15589 22891 15623
rect 22833 15583 22891 15589
rect 13078 15512 13084 15564
rect 13136 15512 13142 15564
rect 13722 15512 13728 15564
rect 13780 15552 13786 15564
rect 15933 15555 15991 15561
rect 15933 15552 15945 15555
rect 13780 15524 15945 15552
rect 13780 15512 13786 15524
rect 15933 15521 15945 15524
rect 15979 15521 15991 15555
rect 15933 15515 15991 15521
rect 16025 15555 16083 15561
rect 16025 15521 16037 15555
rect 16071 15552 16083 15555
rect 17313 15555 17371 15561
rect 16071 15524 17264 15552
rect 16071 15521 16083 15524
rect 16025 15515 16083 15521
rect 11149 15487 11207 15493
rect 11149 15484 11161 15487
rect 11072 15456 11161 15484
rect 10966 15447 11024 15453
rect 11149 15453 11161 15456
rect 11195 15453 11207 15487
rect 11149 15447 11207 15453
rect 11379 15487 11437 15493
rect 11379 15453 11391 15487
rect 11425 15484 11437 15487
rect 11698 15484 11704 15496
rect 11425 15456 11704 15484
rect 11425 15453 11437 15456
rect 11379 15447 11437 15453
rect 6365 15419 6423 15425
rect 6365 15385 6377 15419
rect 6411 15416 6423 15419
rect 6822 15416 6828 15428
rect 6411 15388 6828 15416
rect 6411 15385 6423 15388
rect 6365 15379 6423 15385
rect 6822 15376 6828 15388
rect 6880 15416 6886 15428
rect 8297 15419 8355 15425
rect 6880 15388 8064 15416
rect 6880 15376 6886 15388
rect 7006 15348 7012 15360
rect 6288 15320 7012 15348
rect 7006 15308 7012 15320
rect 7064 15308 7070 15360
rect 7926 15308 7932 15360
rect 7984 15308 7990 15360
rect 8036 15348 8064 15388
rect 8297 15385 8309 15419
rect 8343 15416 8355 15419
rect 9214 15416 9220 15428
rect 8343 15388 9220 15416
rect 8343 15385 8355 15388
rect 8297 15379 8355 15385
rect 9214 15376 9220 15388
rect 9272 15376 9278 15428
rect 9668 15419 9726 15425
rect 9668 15385 9680 15419
rect 9714 15416 9726 15419
rect 9950 15416 9956 15428
rect 9714 15388 9956 15416
rect 9714 15385 9726 15388
rect 9668 15379 9726 15385
rect 9950 15376 9956 15388
rect 10008 15376 10014 15428
rect 10980 15416 11008 15447
rect 11698 15444 11704 15456
rect 11756 15444 11762 15496
rect 12250 15444 12256 15496
rect 12308 15484 12314 15496
rect 15378 15484 15384 15496
rect 12308 15456 15384 15484
rect 12308 15444 12314 15456
rect 15378 15444 15384 15456
rect 15436 15444 15442 15496
rect 15657 15487 15715 15493
rect 15657 15453 15669 15487
rect 15703 15484 15715 15487
rect 15746 15484 15752 15496
rect 15703 15456 15752 15484
rect 15703 15453 15715 15456
rect 15657 15447 15715 15453
rect 15746 15444 15752 15456
rect 15804 15444 15810 15496
rect 15838 15444 15844 15496
rect 15896 15444 15902 15496
rect 16114 15444 16120 15496
rect 16172 15484 16178 15496
rect 16209 15487 16267 15493
rect 16209 15484 16221 15487
rect 16172 15456 16221 15484
rect 16172 15444 16178 15456
rect 16209 15453 16221 15456
rect 16255 15453 16267 15487
rect 17236 15484 17264 15524
rect 17313 15521 17325 15555
rect 17359 15552 17371 15555
rect 17494 15552 17500 15564
rect 17359 15524 17500 15552
rect 17359 15521 17371 15524
rect 17313 15515 17371 15521
rect 17494 15512 17500 15524
rect 17552 15512 17558 15564
rect 20530 15512 20536 15564
rect 20588 15512 20594 15564
rect 20717 15555 20775 15561
rect 20717 15521 20729 15555
rect 20763 15552 20775 15555
rect 20990 15552 20996 15564
rect 20763 15524 20996 15552
rect 20763 15521 20775 15524
rect 20717 15515 20775 15521
rect 20990 15512 20996 15524
rect 21048 15512 21054 15564
rect 22922 15512 22928 15564
rect 22980 15552 22986 15564
rect 23934 15552 23940 15564
rect 22980 15524 23940 15552
rect 22980 15512 22986 15524
rect 23934 15512 23940 15524
rect 23992 15512 23998 15564
rect 24026 15512 24032 15564
rect 24084 15512 24090 15564
rect 24136 15552 24164 15648
rect 26510 15580 26516 15632
rect 26568 15620 26574 15632
rect 26896 15620 26924 15648
rect 27801 15623 27859 15629
rect 27801 15620 27813 15623
rect 26568 15592 26924 15620
rect 27264 15592 27813 15620
rect 26568 15580 26574 15592
rect 27264 15564 27292 15592
rect 27801 15589 27813 15592
rect 27847 15620 27859 15623
rect 27985 15623 28043 15629
rect 27985 15620 27997 15623
rect 27847 15592 27997 15620
rect 27847 15589 27859 15592
rect 27801 15583 27859 15589
rect 27985 15589 27997 15592
rect 28031 15589 28043 15623
rect 27985 15583 28043 15589
rect 28920 15592 29224 15620
rect 24394 15552 24400 15564
rect 24136 15524 24400 15552
rect 24394 15512 24400 15524
rect 24452 15512 24458 15564
rect 26786 15512 26792 15564
rect 26844 15552 26850 15564
rect 26881 15555 26939 15561
rect 26881 15552 26893 15555
rect 26844 15524 26893 15552
rect 26844 15512 26850 15524
rect 26881 15521 26893 15524
rect 26927 15521 26939 15555
rect 26881 15515 26939 15521
rect 27157 15555 27215 15561
rect 27157 15521 27169 15555
rect 27203 15552 27215 15555
rect 27246 15552 27252 15564
rect 27203 15524 27252 15552
rect 27203 15521 27215 15524
rect 27157 15515 27215 15521
rect 27246 15512 27252 15524
rect 27304 15512 27310 15564
rect 27430 15512 27436 15564
rect 27488 15552 27494 15564
rect 28920 15561 28948 15592
rect 28905 15555 28963 15561
rect 28905 15552 28917 15555
rect 27488 15524 28917 15552
rect 27488 15512 27494 15524
rect 28905 15521 28917 15524
rect 28951 15521 28963 15555
rect 28905 15515 28963 15521
rect 29086 15512 29092 15564
rect 29144 15512 29150 15564
rect 29196 15552 29224 15592
rect 29196 15524 30512 15552
rect 18046 15484 18052 15496
rect 17236 15456 18052 15484
rect 16209 15447 16267 15453
rect 18046 15444 18052 15456
rect 18104 15484 18110 15496
rect 19058 15484 19064 15496
rect 18104 15456 19064 15484
rect 18104 15444 18110 15456
rect 19058 15444 19064 15456
rect 19116 15444 19122 15496
rect 19245 15487 19303 15493
rect 19245 15453 19257 15487
rect 19291 15453 19303 15487
rect 19245 15447 19303 15453
rect 10796 15388 11008 15416
rect 11241 15419 11299 15425
rect 10796 15360 10824 15388
rect 11241 15385 11253 15419
rect 11287 15416 11299 15419
rect 11287 15388 11744 15416
rect 11287 15385 11299 15388
rect 11241 15379 11299 15385
rect 8389 15351 8447 15357
rect 8389 15348 8401 15351
rect 8036 15320 8401 15348
rect 8389 15317 8401 15320
rect 8435 15317 8447 15351
rect 8389 15311 8447 15317
rect 9030 15308 9036 15360
rect 9088 15308 9094 15360
rect 10778 15308 10784 15360
rect 10836 15308 10842 15360
rect 11514 15308 11520 15360
rect 11572 15308 11578 15360
rect 11716 15357 11744 15388
rect 12618 15376 12624 15428
rect 12676 15416 12682 15428
rect 12814 15419 12872 15425
rect 12814 15416 12826 15419
rect 12676 15388 12826 15416
rect 12676 15376 12682 15388
rect 12814 15385 12826 15388
rect 12860 15385 12872 15419
rect 12814 15379 12872 15385
rect 14734 15376 14740 15428
rect 14792 15416 14798 15428
rect 15473 15419 15531 15425
rect 15473 15416 15485 15419
rect 14792 15388 15485 15416
rect 14792 15376 14798 15388
rect 15473 15385 15485 15388
rect 15519 15416 15531 15419
rect 16485 15419 16543 15425
rect 16485 15416 16497 15419
rect 15519 15388 16497 15416
rect 15519 15385 15531 15388
rect 15473 15379 15531 15385
rect 16485 15385 16497 15388
rect 16531 15385 16543 15419
rect 16485 15379 16543 15385
rect 17764 15419 17822 15425
rect 17764 15385 17776 15419
rect 17810 15416 17822 15419
rect 17954 15416 17960 15428
rect 17810 15388 17960 15416
rect 17810 15385 17822 15388
rect 17764 15379 17822 15385
rect 17954 15376 17960 15388
rect 18012 15376 18018 15428
rect 19260 15416 19288 15447
rect 19426 15444 19432 15496
rect 19484 15484 19490 15496
rect 21269 15487 21327 15493
rect 21269 15484 21281 15487
rect 19484 15456 21281 15484
rect 19484 15444 19490 15456
rect 21269 15453 21281 15456
rect 21315 15453 21327 15487
rect 21269 15447 21327 15453
rect 21358 15444 21364 15496
rect 21416 15484 21422 15496
rect 24044 15484 24072 15512
rect 21416 15456 24072 15484
rect 21416 15444 21422 15456
rect 24670 15444 24676 15496
rect 24728 15484 24734 15496
rect 25409 15487 25467 15493
rect 25409 15484 25421 15487
rect 24728 15456 25421 15484
rect 24728 15444 24734 15456
rect 25409 15453 25421 15456
rect 25455 15453 25467 15487
rect 25409 15447 25467 15453
rect 27798 15444 27804 15496
rect 27856 15484 27862 15496
rect 29549 15487 29607 15493
rect 29549 15484 29561 15487
rect 27856 15456 29561 15484
rect 27856 15444 27862 15456
rect 29549 15453 29561 15456
rect 29595 15484 29607 15487
rect 30374 15484 30380 15496
rect 29595 15456 30380 15484
rect 29595 15453 29607 15456
rect 29549 15447 29607 15453
rect 30374 15444 30380 15456
rect 30432 15444 30438 15496
rect 20441 15419 20499 15425
rect 19260 15388 19932 15416
rect 11701 15351 11759 15357
rect 11701 15317 11713 15351
rect 11747 15348 11759 15351
rect 12434 15348 12440 15360
rect 11747 15320 12440 15348
rect 11747 15317 11759 15320
rect 11701 15311 11759 15317
rect 12434 15308 12440 15320
rect 12492 15308 12498 15360
rect 12894 15308 12900 15360
rect 12952 15348 12958 15360
rect 13173 15351 13231 15357
rect 13173 15348 13185 15351
rect 12952 15320 13185 15348
rect 12952 15308 12958 15320
rect 13173 15317 13185 15320
rect 13219 15317 13231 15351
rect 13173 15311 13231 15317
rect 16390 15308 16396 15360
rect 16448 15308 16454 15360
rect 19904 15357 19932 15388
rect 20441 15385 20453 15419
rect 20487 15416 20499 15419
rect 20714 15416 20720 15428
rect 20487 15388 20720 15416
rect 20487 15385 20499 15388
rect 20441 15379 20499 15385
rect 20714 15376 20720 15388
rect 20772 15376 20778 15428
rect 21536 15419 21594 15425
rect 21536 15385 21548 15419
rect 21582 15416 21594 15419
rect 21818 15416 21824 15428
rect 21582 15388 21824 15416
rect 21582 15385 21594 15388
rect 21536 15379 21594 15385
rect 21818 15376 21824 15388
rect 21876 15376 21882 15428
rect 23934 15376 23940 15428
rect 23992 15416 23998 15428
rect 24857 15419 24915 15425
rect 24857 15416 24869 15419
rect 23992 15388 24869 15416
rect 23992 15376 23998 15388
rect 24857 15385 24869 15388
rect 24903 15416 24915 15419
rect 25314 15416 25320 15428
rect 24903 15388 25320 15416
rect 24903 15385 24915 15388
rect 24857 15379 24915 15385
rect 25314 15376 25320 15388
rect 25372 15376 25378 15428
rect 25676 15419 25734 15425
rect 25676 15385 25688 15419
rect 25722 15416 25734 15419
rect 26050 15416 26056 15428
rect 25722 15388 26056 15416
rect 25722 15385 25734 15388
rect 25676 15379 25734 15385
rect 26050 15376 26056 15388
rect 26108 15376 26114 15428
rect 28813 15419 28871 15425
rect 28813 15385 28825 15419
rect 28859 15416 28871 15419
rect 29178 15416 29184 15428
rect 28859 15388 29184 15416
rect 28859 15385 28871 15388
rect 28813 15379 28871 15385
rect 29178 15376 29184 15388
rect 29236 15376 29242 15428
rect 30484 15416 30512 15524
rect 30650 15493 30656 15496
rect 30644 15484 30656 15493
rect 30611 15456 30656 15484
rect 30644 15447 30656 15456
rect 30650 15444 30656 15447
rect 30708 15444 30714 15496
rect 33413 15487 33471 15493
rect 33413 15453 33425 15487
rect 33459 15453 33471 15487
rect 33413 15447 33471 15453
rect 34517 15487 34575 15493
rect 34517 15453 34529 15487
rect 34563 15484 34575 15487
rect 34790 15484 34796 15496
rect 34563 15456 34796 15484
rect 34563 15453 34575 15456
rect 34517 15447 34575 15453
rect 30834 15416 30840 15428
rect 30484 15388 30840 15416
rect 30834 15376 30840 15388
rect 30892 15376 30898 15428
rect 31202 15376 31208 15428
rect 31260 15416 31266 15428
rect 31941 15419 31999 15425
rect 31941 15416 31953 15419
rect 31260 15388 31953 15416
rect 31260 15376 31266 15388
rect 31941 15385 31953 15388
rect 31987 15416 31999 15419
rect 32309 15419 32367 15425
rect 32309 15416 32321 15419
rect 31987 15388 32321 15416
rect 31987 15385 31999 15388
rect 31941 15379 31999 15385
rect 32309 15385 32321 15388
rect 32355 15385 32367 15419
rect 32309 15379 32367 15385
rect 33042 15376 33048 15428
rect 33100 15416 33106 15428
rect 33428 15416 33456 15447
rect 34790 15444 34796 15456
rect 34848 15444 34854 15496
rect 33100 15388 33456 15416
rect 34241 15419 34299 15425
rect 33100 15376 33106 15388
rect 34241 15385 34253 15419
rect 34287 15416 34299 15419
rect 34698 15416 34704 15428
rect 34287 15388 34704 15416
rect 34287 15385 34299 15388
rect 34241 15379 34299 15385
rect 34698 15376 34704 15388
rect 34756 15376 34762 15428
rect 19889 15351 19947 15357
rect 19889 15317 19901 15351
rect 19935 15348 19947 15351
rect 20806 15348 20812 15360
rect 19935 15320 20812 15348
rect 19935 15317 19947 15320
rect 19889 15311 19947 15317
rect 20806 15308 20812 15320
rect 20864 15308 20870 15360
rect 20990 15308 20996 15360
rect 21048 15348 21054 15360
rect 21910 15348 21916 15360
rect 21048 15320 21916 15348
rect 21048 15308 21054 15320
rect 21910 15308 21916 15320
rect 21968 15308 21974 15360
rect 24118 15308 24124 15360
rect 24176 15348 24182 15360
rect 24213 15351 24271 15357
rect 24213 15348 24225 15351
rect 24176 15320 24225 15348
rect 24176 15308 24182 15320
rect 24213 15317 24225 15320
rect 24259 15348 24271 15351
rect 24762 15348 24768 15360
rect 24259 15320 24768 15348
rect 24259 15317 24271 15320
rect 24213 15311 24271 15317
rect 24762 15308 24768 15320
rect 24820 15348 24826 15360
rect 25498 15348 25504 15360
rect 24820 15320 25504 15348
rect 24820 15308 24826 15320
rect 25498 15308 25504 15320
rect 25556 15308 25562 15360
rect 29270 15308 29276 15360
rect 29328 15308 29334 15360
rect 30374 15308 30380 15360
rect 30432 15348 30438 15360
rect 30558 15348 30564 15360
rect 30432 15320 30564 15348
rect 30432 15308 30438 15320
rect 30558 15308 30564 15320
rect 30616 15308 30622 15360
rect 31478 15308 31484 15360
rect 31536 15348 31542 15360
rect 32125 15351 32183 15357
rect 32125 15348 32137 15351
rect 31536 15320 32137 15348
rect 31536 15308 31542 15320
rect 32125 15317 32137 15320
rect 32171 15317 32183 15351
rect 32125 15311 32183 15317
rect 1104 15258 35328 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35328 15258
rect 1104 15184 35328 15206
rect 2866 15104 2872 15156
rect 2924 15104 2930 15156
rect 3234 15104 3240 15156
rect 3292 15104 3298 15156
rect 3694 15104 3700 15156
rect 3752 15104 3758 15156
rect 4154 15104 4160 15156
rect 4212 15104 4218 15156
rect 4614 15104 4620 15156
rect 4672 15104 4678 15156
rect 8757 15147 8815 15153
rect 8757 15113 8769 15147
rect 8803 15144 8815 15147
rect 9214 15144 9220 15156
rect 8803 15116 9220 15144
rect 8803 15113 8815 15116
rect 8757 15107 8815 15113
rect 9214 15104 9220 15116
rect 9272 15104 9278 15156
rect 9950 15104 9956 15156
rect 10008 15104 10014 15156
rect 10321 15147 10379 15153
rect 10321 15113 10333 15147
rect 10367 15144 10379 15147
rect 10778 15144 10784 15156
rect 10367 15116 10784 15144
rect 10367 15113 10379 15116
rect 10321 15107 10379 15113
rect 10778 15104 10784 15116
rect 10836 15104 10842 15156
rect 12161 15147 12219 15153
rect 10888 15116 11928 15144
rect 10888 15088 10916 15116
rect 3329 15079 3387 15085
rect 3329 15045 3341 15079
rect 3375 15076 3387 15079
rect 4062 15076 4068 15088
rect 3375 15048 4068 15076
rect 3375 15045 3387 15048
rect 3329 15039 3387 15045
rect 4062 15036 4068 15048
rect 4120 15076 4126 15088
rect 4525 15079 4583 15085
rect 4525 15076 4537 15079
rect 4120 15048 4537 15076
rect 4120 15036 4126 15048
rect 4525 15045 4537 15048
rect 4571 15045 4583 15079
rect 9306 15076 9312 15088
rect 4525 15039 4583 15045
rect 7392 15048 9312 15076
rect 1302 14968 1308 15020
rect 1360 15008 1366 15020
rect 7392 15017 7420 15048
rect 9306 15036 9312 15048
rect 9364 15036 9370 15088
rect 10413 15079 10471 15085
rect 10413 15045 10425 15079
rect 10459 15076 10471 15079
rect 10870 15076 10876 15088
rect 10459 15048 10876 15076
rect 10459 15045 10471 15048
rect 10413 15039 10471 15045
rect 10870 15036 10876 15048
rect 10928 15036 10934 15088
rect 11330 15036 11336 15088
rect 11388 15076 11394 15088
rect 11517 15079 11575 15085
rect 11517 15076 11529 15079
rect 11388 15048 11529 15076
rect 11388 15036 11394 15048
rect 11517 15045 11529 15048
rect 11563 15045 11575 15079
rect 11517 15039 11575 15045
rect 1397 15011 1455 15017
rect 1397 15008 1409 15011
rect 1360 14980 1409 15008
rect 1360 14968 1366 14980
rect 1397 14977 1409 14980
rect 1443 15008 1455 15011
rect 1857 15011 1915 15017
rect 1857 15008 1869 15011
rect 1443 14980 1869 15008
rect 1443 14977 1455 14980
rect 1397 14971 1455 14977
rect 1857 14977 1869 14980
rect 1903 14977 1915 15011
rect 1857 14971 1915 14977
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 7644 15011 7702 15017
rect 7644 14977 7656 15011
rect 7690 15008 7702 15011
rect 7926 15008 7932 15020
rect 7690 14980 7932 15008
rect 7690 14977 7702 14980
rect 7644 14971 7702 14977
rect 7926 14968 7932 14980
rect 7984 14968 7990 15020
rect 8018 14968 8024 15020
rect 8076 15008 8082 15020
rect 8076 14980 10548 15008
rect 8076 14968 8082 14980
rect 3513 14943 3571 14949
rect 3513 14909 3525 14943
rect 3559 14940 3571 14943
rect 3694 14940 3700 14952
rect 3559 14912 3700 14940
rect 3559 14909 3571 14912
rect 3513 14903 3571 14909
rect 3694 14900 3700 14912
rect 3752 14900 3758 14952
rect 4801 14943 4859 14949
rect 4801 14909 4813 14943
rect 4847 14940 4859 14943
rect 5350 14940 5356 14952
rect 4847 14912 5356 14940
rect 4847 14909 4859 14912
rect 4801 14903 4859 14909
rect 5350 14900 5356 14912
rect 5408 14900 5414 14952
rect 10520 14949 10548 14980
rect 11238 14968 11244 15020
rect 11296 15008 11302 15020
rect 11793 15011 11851 15017
rect 11793 15008 11805 15011
rect 11296 14980 11805 15008
rect 11296 14968 11302 14980
rect 11793 14977 11805 14980
rect 11839 14977 11851 15011
rect 11900 15008 11928 15116
rect 12161 15113 12173 15147
rect 12207 15144 12219 15147
rect 12618 15144 12624 15156
rect 12207 15116 12624 15144
rect 12207 15113 12219 15116
rect 12161 15107 12219 15113
rect 12618 15104 12624 15116
rect 12676 15104 12682 15156
rect 12802 15104 12808 15156
rect 12860 15144 12866 15156
rect 13081 15147 13139 15153
rect 13081 15144 13093 15147
rect 12860 15116 13093 15144
rect 12860 15104 12866 15116
rect 13081 15113 13093 15116
rect 13127 15144 13139 15147
rect 14918 15144 14924 15156
rect 13127 15116 14924 15144
rect 13127 15113 13139 15116
rect 13081 15107 13139 15113
rect 14918 15104 14924 15116
rect 14976 15104 14982 15156
rect 15473 15147 15531 15153
rect 15473 15113 15485 15147
rect 15519 15144 15531 15147
rect 15654 15144 15660 15156
rect 15519 15116 15660 15144
rect 15519 15113 15531 15116
rect 15473 15107 15531 15113
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 16206 15104 16212 15156
rect 16264 15144 16270 15156
rect 17037 15147 17095 15153
rect 17037 15144 17049 15147
rect 16264 15116 17049 15144
rect 16264 15104 16270 15116
rect 17037 15113 17049 15116
rect 17083 15113 17095 15147
rect 17037 15107 17095 15113
rect 17954 15104 17960 15156
rect 18012 15104 18018 15156
rect 18325 15147 18383 15153
rect 18325 15113 18337 15147
rect 18371 15144 18383 15147
rect 18966 15144 18972 15156
rect 18371 15116 18972 15144
rect 18371 15113 18383 15116
rect 18325 15107 18383 15113
rect 18966 15104 18972 15116
rect 19024 15104 19030 15156
rect 20441 15147 20499 15153
rect 20441 15144 20453 15147
rect 19306 15116 20453 15144
rect 16224 15076 16252 15104
rect 12728 15048 16252 15076
rect 12529 15011 12587 15017
rect 12529 15008 12541 15011
rect 11900 14980 12541 15008
rect 11793 14971 11851 14977
rect 12529 14977 12541 14980
rect 12575 15008 12587 15011
rect 12728 15008 12756 15048
rect 16390 15036 16396 15088
rect 16448 15036 16454 15088
rect 18417 15079 18475 15085
rect 18417 15045 18429 15079
rect 18463 15076 18475 15079
rect 19306 15076 19334 15116
rect 20441 15113 20453 15116
rect 20487 15144 20499 15147
rect 20530 15144 20536 15156
rect 20487 15116 20536 15144
rect 20487 15113 20499 15116
rect 20441 15107 20499 15113
rect 20530 15104 20536 15116
rect 20588 15104 20594 15156
rect 20714 15104 20720 15156
rect 20772 15144 20778 15156
rect 20772 15116 21220 15144
rect 20772 15104 20778 15116
rect 21192 15085 21220 15116
rect 21450 15104 21456 15156
rect 21508 15104 21514 15156
rect 21818 15104 21824 15156
rect 21876 15104 21882 15156
rect 22189 15147 22247 15153
rect 22189 15113 22201 15147
rect 22235 15144 22247 15147
rect 22554 15144 22560 15156
rect 22235 15116 22560 15144
rect 22235 15113 22247 15116
rect 22189 15107 22247 15113
rect 22554 15104 22560 15116
rect 22612 15104 22618 15156
rect 23566 15104 23572 15156
rect 23624 15104 23630 15156
rect 23937 15147 23995 15153
rect 23937 15113 23949 15147
rect 23983 15144 23995 15147
rect 24026 15144 24032 15156
rect 23983 15116 24032 15144
rect 23983 15113 23995 15116
rect 23937 15107 23995 15113
rect 24026 15104 24032 15116
rect 24084 15104 24090 15156
rect 24210 15104 24216 15156
rect 24268 15144 24274 15156
rect 24305 15147 24363 15153
rect 24305 15144 24317 15147
rect 24268 15116 24317 15144
rect 24268 15104 24274 15116
rect 24305 15113 24317 15116
rect 24351 15113 24363 15147
rect 24305 15107 24363 15113
rect 26053 15147 26111 15153
rect 26053 15113 26065 15147
rect 26099 15144 26111 15147
rect 26234 15144 26240 15156
rect 26099 15116 26240 15144
rect 26099 15113 26111 15116
rect 26053 15107 26111 15113
rect 26234 15104 26240 15116
rect 26292 15144 26298 15156
rect 27062 15144 27068 15156
rect 26292 15116 27068 15144
rect 26292 15104 26298 15116
rect 27062 15104 27068 15116
rect 27120 15104 27126 15156
rect 29730 15104 29736 15156
rect 29788 15104 29794 15156
rect 30006 15104 30012 15156
rect 30064 15104 30070 15156
rect 30558 15104 30564 15156
rect 30616 15104 30622 15156
rect 30926 15104 30932 15156
rect 30984 15144 30990 15156
rect 30984 15116 32352 15144
rect 30984 15104 30990 15116
rect 18463 15048 19334 15076
rect 20349 15079 20407 15085
rect 18463 15045 18475 15048
rect 18417 15039 18475 15045
rect 20349 15045 20361 15079
rect 20395 15076 20407 15079
rect 21177 15079 21235 15085
rect 20395 15048 20944 15076
rect 20395 15045 20407 15048
rect 20349 15039 20407 15045
rect 12575 14980 12756 15008
rect 14360 15011 14418 15017
rect 12575 14977 12587 14980
rect 12529 14971 12587 14977
rect 14360 14977 14372 15011
rect 14406 15008 14418 15011
rect 14642 15008 14648 15020
rect 14406 14980 14648 15008
rect 14406 14977 14418 14980
rect 14360 14971 14418 14977
rect 14642 14968 14648 14980
rect 14700 14968 14706 15020
rect 16301 15011 16359 15017
rect 16301 14977 16313 15011
rect 16347 15008 16359 15011
rect 16408 15008 16436 15036
rect 20916 15020 20944 15048
rect 21177 15045 21189 15079
rect 21223 15045 21235 15079
rect 21177 15039 21235 15045
rect 22066 15048 28028 15076
rect 16347 14980 19334 15008
rect 16347 14977 16359 14980
rect 16301 14971 16359 14977
rect 10505 14943 10563 14949
rect 10505 14909 10517 14943
rect 10551 14940 10563 14943
rect 10781 14943 10839 14949
rect 10781 14940 10793 14943
rect 10551 14912 10793 14940
rect 10551 14909 10563 14912
rect 10505 14903 10563 14909
rect 10781 14909 10793 14912
rect 10827 14909 10839 14943
rect 10781 14903 10839 14909
rect 11422 14900 11428 14952
rect 11480 14940 11486 14952
rect 11609 14943 11667 14949
rect 11609 14940 11621 14943
rect 11480 14912 11621 14940
rect 11480 14900 11486 14912
rect 11609 14909 11621 14912
rect 11655 14909 11667 14943
rect 11609 14903 11667 14909
rect 12618 14900 12624 14952
rect 12676 14900 12682 14952
rect 12802 14900 12808 14952
rect 12860 14900 12866 14952
rect 14093 14943 14151 14949
rect 14093 14909 14105 14943
rect 14139 14909 14151 14943
rect 14093 14903 14151 14909
rect 1581 14875 1639 14881
rect 1581 14841 1593 14875
rect 1627 14872 1639 14875
rect 1765 14875 1823 14881
rect 1765 14872 1777 14875
rect 1627 14844 1777 14872
rect 1627 14841 1639 14844
rect 1581 14835 1639 14841
rect 1765 14841 1777 14844
rect 1811 14872 1823 14875
rect 11977 14875 12035 14881
rect 1811 14844 7420 14872
rect 1811 14841 1823 14844
rect 1765 14835 1823 14841
rect 3694 14764 3700 14816
rect 3752 14804 3758 14816
rect 4798 14804 4804 14816
rect 3752 14776 4804 14804
rect 3752 14764 3758 14776
rect 4798 14764 4804 14776
rect 4856 14764 4862 14816
rect 5077 14807 5135 14813
rect 5077 14773 5089 14807
rect 5123 14804 5135 14807
rect 5350 14804 5356 14816
rect 5123 14776 5356 14804
rect 5123 14773 5135 14776
rect 5077 14767 5135 14773
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 5442 14764 5448 14816
rect 5500 14804 5506 14816
rect 5997 14807 6055 14813
rect 5997 14804 6009 14807
rect 5500 14776 6009 14804
rect 5500 14764 5506 14776
rect 5997 14773 6009 14776
rect 6043 14804 6055 14807
rect 6362 14804 6368 14816
rect 6043 14776 6368 14804
rect 6043 14773 6055 14776
rect 5997 14767 6055 14773
rect 6362 14764 6368 14776
rect 6420 14764 6426 14816
rect 7392 14804 7420 14844
rect 8312 14844 11652 14872
rect 8312 14804 8340 14844
rect 7392 14776 8340 14804
rect 11238 14764 11244 14816
rect 11296 14764 11302 14816
rect 11514 14764 11520 14816
rect 11572 14764 11578 14816
rect 11624 14804 11652 14844
rect 11977 14841 11989 14875
rect 12023 14872 12035 14875
rect 13722 14872 13728 14884
rect 12023 14844 13728 14872
rect 12023 14841 12035 14844
rect 11977 14835 12035 14841
rect 13722 14832 13728 14844
rect 13780 14832 13786 14884
rect 13998 14804 14004 14816
rect 11624 14776 14004 14804
rect 13998 14764 14004 14776
rect 14056 14764 14062 14816
rect 14108 14804 14136 14903
rect 16114 14900 16120 14952
rect 16172 14940 16178 14952
rect 17129 14943 17187 14949
rect 17129 14940 17141 14943
rect 16172 14912 17141 14940
rect 16172 14900 16178 14912
rect 17129 14909 17141 14912
rect 17175 14909 17187 14943
rect 17129 14903 17187 14909
rect 17313 14943 17371 14949
rect 17313 14909 17325 14943
rect 17359 14940 17371 14943
rect 18601 14943 18659 14949
rect 17359 14912 17632 14940
rect 17359 14909 17371 14912
rect 17313 14903 17371 14909
rect 17604 14816 17632 14912
rect 18601 14909 18613 14943
rect 18647 14909 18659 14943
rect 18601 14903 18659 14909
rect 17770 14832 17776 14884
rect 17828 14872 17834 14884
rect 17865 14875 17923 14881
rect 17865 14872 17877 14875
rect 17828 14844 17877 14872
rect 17828 14832 17834 14844
rect 17865 14841 17877 14844
rect 17911 14872 17923 14875
rect 18616 14872 18644 14903
rect 17911 14844 18644 14872
rect 19306 14872 19334 14980
rect 19518 14968 19524 15020
rect 19576 15008 19582 15020
rect 20809 15011 20867 15017
rect 20809 15008 20821 15011
rect 19576 14980 20821 15008
rect 19576 14968 19582 14980
rect 20809 14977 20821 14980
rect 20855 14977 20867 15011
rect 20809 14971 20867 14977
rect 20898 14968 20904 15020
rect 20956 14968 20962 15020
rect 21082 14968 21088 15020
rect 21140 14968 21146 15020
rect 21315 15011 21373 15017
rect 21315 14977 21327 15011
rect 21361 15008 21373 15011
rect 21726 15008 21732 15020
rect 21361 14980 21732 15008
rect 21361 14977 21373 14980
rect 21315 14971 21373 14977
rect 21726 14968 21732 14980
rect 21784 14968 21790 15020
rect 20530 14900 20536 14952
rect 20588 14900 20594 14952
rect 22066 14940 22094 15048
rect 22281 15011 22339 15017
rect 22281 14977 22293 15011
rect 22327 15008 22339 15011
rect 22646 15008 22652 15020
rect 22327 14980 22652 15008
rect 22327 14977 22339 14980
rect 22281 14971 22339 14977
rect 22646 14968 22652 14980
rect 22704 14968 22710 15020
rect 23385 15011 23443 15017
rect 23385 14977 23397 15011
rect 23431 15008 23443 15011
rect 23474 15008 23480 15020
rect 23431 14980 23480 15008
rect 23431 14977 23443 14980
rect 23385 14971 23443 14977
rect 23474 14968 23480 14980
rect 23532 14968 23538 15020
rect 23753 15011 23811 15017
rect 23753 14977 23765 15011
rect 23799 15008 23811 15011
rect 24118 15008 24124 15020
rect 23799 14980 24124 15008
rect 23799 14977 23811 14980
rect 23753 14971 23811 14977
rect 24118 14968 24124 14980
rect 24176 14968 24182 15020
rect 24210 14968 24216 15020
rect 24268 14968 24274 15020
rect 24670 14968 24676 15020
rect 24728 14968 24734 15020
rect 24940 15011 24998 15017
rect 24940 14977 24952 15011
rect 24986 15008 24998 15011
rect 25222 15008 25228 15020
rect 24986 14980 25228 15008
rect 24986 14977 24998 14980
rect 24940 14971 24998 14977
rect 25222 14968 25228 14980
rect 25280 14968 25286 15020
rect 26145 15011 26203 15017
rect 26145 14977 26157 15011
rect 26191 15008 26203 15011
rect 26789 15011 26847 15017
rect 26789 15008 26801 15011
rect 26191 14980 26801 15008
rect 26191 14977 26203 14980
rect 26145 14971 26203 14977
rect 26789 14977 26801 14980
rect 26835 15008 26847 15011
rect 26878 15008 26884 15020
rect 26835 14980 26884 15008
rect 26835 14977 26847 14980
rect 26789 14971 26847 14977
rect 26878 14968 26884 14980
rect 26936 14968 26942 15020
rect 27062 14968 27068 15020
rect 27120 15008 27126 15020
rect 27229 15011 27287 15017
rect 27229 15008 27241 15011
rect 27120 14980 27241 15008
rect 27120 14968 27126 14980
rect 27229 14977 27241 14980
rect 27275 14977 27287 15011
rect 27229 14971 27287 14977
rect 20640 14912 22094 14940
rect 20640 14872 20668 14912
rect 22462 14900 22468 14952
rect 22520 14900 22526 14952
rect 26970 14900 26976 14952
rect 27028 14900 27034 14952
rect 28000 14940 28028 15048
rect 28902 15036 28908 15088
rect 28960 15076 28966 15088
rect 28960 15048 29132 15076
rect 28960 15036 28966 15048
rect 28445 15011 28503 15017
rect 28445 14977 28457 15011
rect 28491 15008 28503 15011
rect 28534 15008 28540 15020
rect 28491 14980 28540 15008
rect 28491 14977 28503 14980
rect 28445 14971 28503 14977
rect 28534 14968 28540 14980
rect 28592 15008 28598 15020
rect 28718 15008 28724 15020
rect 28592 14980 28724 15008
rect 28592 14968 28598 14980
rect 28718 14968 28724 14980
rect 28776 14968 28782 15020
rect 29104 15017 29132 15048
rect 29914 15036 29920 15088
rect 29972 15036 29978 15088
rect 30466 15036 30472 15088
rect 30524 15036 30530 15088
rect 29089 15011 29147 15017
rect 29089 14977 29101 15011
rect 29135 14977 29147 15011
rect 29089 14971 29147 14977
rect 29178 14968 29184 15020
rect 29236 15008 29242 15020
rect 29236 14980 29281 15008
rect 29236 14968 29242 14980
rect 29362 14968 29368 15020
rect 29420 14968 29426 15020
rect 29454 14968 29460 15020
rect 29512 14968 29518 15020
rect 29546 14968 29552 15020
rect 29604 15017 29610 15020
rect 29604 15011 29653 15017
rect 29604 14977 29607 15011
rect 29641 15008 29653 15011
rect 30190 15008 30196 15020
rect 29641 14980 30196 15008
rect 29641 14977 29653 14980
rect 29604 14971 29653 14977
rect 29604 14968 29610 14971
rect 30190 14968 30196 14980
rect 30248 14968 30254 15020
rect 30576 15008 30604 15104
rect 31018 15036 31024 15088
rect 31076 15076 31082 15088
rect 32324 15085 32352 15116
rect 32674 15104 32680 15156
rect 32732 15104 32738 15156
rect 33134 15104 33140 15156
rect 33192 15144 33198 15156
rect 33192 15116 33548 15144
rect 33192 15104 33198 15116
rect 31665 15079 31723 15085
rect 31665 15076 31677 15079
rect 31076 15048 31677 15076
rect 31076 15036 31082 15048
rect 31665 15045 31677 15048
rect 31711 15045 31723 15079
rect 31665 15039 31723 15045
rect 32309 15079 32367 15085
rect 32309 15045 32321 15079
rect 32355 15045 32367 15079
rect 32309 15039 32367 15045
rect 32401 15079 32459 15085
rect 32401 15045 32413 15079
rect 32447 15076 32459 15079
rect 33410 15076 33416 15088
rect 32447 15048 33416 15076
rect 32447 15045 32459 15048
rect 32401 15039 32459 15045
rect 33410 15036 33416 15048
rect 33468 15036 33474 15088
rect 33520 15076 33548 15116
rect 33520 15048 33994 15076
rect 30929 15011 30987 15017
rect 30929 15008 30941 15011
rect 30576 14980 30941 15008
rect 30929 14977 30941 14980
rect 30975 15008 30987 15011
rect 31205 15011 31263 15017
rect 31205 15008 31217 15011
rect 30975 14980 31217 15008
rect 30975 14977 30987 14980
rect 30929 14971 30987 14977
rect 31205 14977 31217 14980
rect 31251 15008 31263 15011
rect 31389 15011 31447 15017
rect 31389 15008 31401 15011
rect 31251 14980 31401 15008
rect 31251 14977 31263 14980
rect 31205 14971 31263 14977
rect 31389 14977 31401 14980
rect 31435 14977 31447 15011
rect 31389 14971 31447 14977
rect 31846 14968 31852 15020
rect 31904 15008 31910 15020
rect 32125 15011 32183 15017
rect 32125 15008 32137 15011
rect 31904 14980 32137 15008
rect 31904 14968 31910 14980
rect 32125 14977 32137 14980
rect 32171 14977 32183 15011
rect 32125 14971 32183 14977
rect 32493 15011 32551 15017
rect 32493 14977 32505 15011
rect 32539 15008 32551 15011
rect 32582 15008 32588 15020
rect 32539 14980 32588 15008
rect 32539 14977 32551 14980
rect 32493 14971 32551 14977
rect 32582 14968 32588 14980
rect 32640 14968 32646 15020
rect 33229 14943 33287 14949
rect 28000 14912 31754 14940
rect 24026 14872 24032 14884
rect 19306 14844 20668 14872
rect 22066 14844 24032 14872
rect 17911 14841 17923 14844
rect 17865 14835 17923 14841
rect 15102 14804 15108 14816
rect 14108 14776 15108 14804
rect 15102 14764 15108 14776
rect 15160 14764 15166 14816
rect 15746 14764 15752 14816
rect 15804 14804 15810 14816
rect 16482 14804 16488 14816
rect 15804 14776 16488 14804
rect 15804 14764 15810 14776
rect 16482 14764 16488 14776
rect 16540 14764 16546 14816
rect 16669 14807 16727 14813
rect 16669 14773 16681 14807
rect 16715 14804 16727 14807
rect 16758 14804 16764 14816
rect 16715 14776 16764 14804
rect 16715 14773 16727 14776
rect 16669 14767 16727 14773
rect 16758 14764 16764 14776
rect 16816 14764 16822 14816
rect 17586 14764 17592 14816
rect 17644 14764 17650 14816
rect 19978 14764 19984 14816
rect 20036 14764 20042 14816
rect 20530 14764 20536 14816
rect 20588 14804 20594 14816
rect 21545 14807 21603 14813
rect 21545 14804 21557 14807
rect 20588 14776 21557 14804
rect 20588 14764 20594 14776
rect 21545 14773 21557 14776
rect 21591 14804 21603 14807
rect 22066 14804 22094 14844
rect 24026 14832 24032 14844
rect 24084 14832 24090 14884
rect 28166 14832 28172 14884
rect 28224 14872 28230 14884
rect 28626 14872 28632 14884
rect 28224 14844 28632 14872
rect 28224 14832 28230 14844
rect 28626 14832 28632 14844
rect 28684 14832 28690 14884
rect 29362 14832 29368 14884
rect 29420 14872 29426 14884
rect 30745 14875 30803 14881
rect 30745 14872 30757 14875
rect 29420 14844 30757 14872
rect 29420 14832 29426 14844
rect 30745 14841 30757 14844
rect 30791 14841 30803 14875
rect 31726 14872 31754 14912
rect 33229 14909 33241 14943
rect 33275 14909 33287 14943
rect 33229 14903 33287 14909
rect 33505 14943 33563 14949
rect 33505 14909 33517 14943
rect 33551 14940 33563 14943
rect 33962 14940 33968 14952
rect 33551 14912 33968 14940
rect 33551 14909 33563 14912
rect 33505 14903 33563 14909
rect 32030 14872 32036 14884
rect 31726 14844 32036 14872
rect 30745 14835 30803 14841
rect 32030 14832 32036 14844
rect 32088 14832 32094 14884
rect 32122 14832 32128 14884
rect 32180 14872 32186 14884
rect 33042 14872 33048 14884
rect 32180 14844 33048 14872
rect 32180 14832 32186 14844
rect 33042 14832 33048 14844
rect 33100 14872 33106 14884
rect 33244 14872 33272 14903
rect 33962 14900 33968 14912
rect 34020 14900 34026 14952
rect 33100 14844 33272 14872
rect 33100 14832 33106 14844
rect 21591 14776 22094 14804
rect 21591 14773 21603 14776
rect 21545 14767 21603 14773
rect 22462 14764 22468 14816
rect 22520 14804 22526 14816
rect 22741 14807 22799 14813
rect 22741 14804 22753 14807
rect 22520 14776 22753 14804
rect 22520 14764 22526 14776
rect 22741 14773 22753 14776
rect 22787 14804 22799 14807
rect 23198 14804 23204 14816
rect 22787 14776 23204 14804
rect 22787 14773 22799 14776
rect 22741 14767 22799 14773
rect 23198 14764 23204 14776
rect 23256 14764 23262 14816
rect 26326 14764 26332 14816
rect 26384 14804 26390 14816
rect 26510 14804 26516 14816
rect 26384 14776 26516 14804
rect 26384 14764 26390 14776
rect 26510 14764 26516 14776
rect 26568 14764 26574 14816
rect 27982 14764 27988 14816
rect 28040 14804 28046 14816
rect 28353 14807 28411 14813
rect 28353 14804 28365 14807
rect 28040 14776 28365 14804
rect 28040 14764 28046 14776
rect 28353 14773 28365 14776
rect 28399 14773 28411 14807
rect 28353 14767 28411 14773
rect 28442 14764 28448 14816
rect 28500 14804 28506 14816
rect 28718 14804 28724 14816
rect 28500 14776 28724 14804
rect 28500 14764 28506 14776
rect 28718 14764 28724 14776
rect 28776 14804 28782 14816
rect 28813 14807 28871 14813
rect 28813 14804 28825 14807
rect 28776 14776 28825 14804
rect 28776 14764 28782 14776
rect 28813 14773 28825 14776
rect 28859 14773 28871 14807
rect 28813 14767 28871 14773
rect 30006 14764 30012 14816
rect 30064 14804 30070 14816
rect 31021 14807 31079 14813
rect 31021 14804 31033 14807
rect 30064 14776 31033 14804
rect 30064 14764 30070 14776
rect 31021 14773 31033 14776
rect 31067 14773 31079 14807
rect 31021 14767 31079 14773
rect 31478 14764 31484 14816
rect 31536 14804 31542 14816
rect 31757 14807 31815 14813
rect 31757 14804 31769 14807
rect 31536 14776 31769 14804
rect 31536 14764 31542 14776
rect 31757 14773 31769 14776
rect 31803 14804 31815 14807
rect 32769 14807 32827 14813
rect 32769 14804 32781 14807
rect 31803 14776 32781 14804
rect 31803 14773 31815 14776
rect 31757 14767 31815 14773
rect 32769 14773 32781 14776
rect 32815 14773 32827 14807
rect 32769 14767 32827 14773
rect 34790 14764 34796 14816
rect 34848 14804 34854 14816
rect 34977 14807 35035 14813
rect 34977 14804 34989 14807
rect 34848 14776 34989 14804
rect 34848 14764 34854 14776
rect 34977 14773 34989 14776
rect 35023 14773 35035 14807
rect 34977 14767 35035 14773
rect 1104 14714 35328 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 35328 14714
rect 1104 14640 35328 14662
rect 3418 14560 3424 14612
rect 3476 14600 3482 14612
rect 3476 14572 12112 14600
rect 3476 14560 3482 14572
rect 6362 14492 6368 14544
rect 6420 14532 6426 14544
rect 11974 14532 11980 14544
rect 6420 14504 11980 14532
rect 6420 14492 6426 14504
rect 11974 14492 11980 14504
rect 12032 14492 12038 14544
rect 12084 14532 12112 14572
rect 12158 14560 12164 14612
rect 12216 14600 12222 14612
rect 12216 14572 14596 14600
rect 12216 14560 12222 14572
rect 14568 14532 14596 14572
rect 14642 14560 14648 14612
rect 14700 14560 14706 14612
rect 15657 14603 15715 14609
rect 14936 14572 15608 14600
rect 14936 14532 14964 14572
rect 12084 14504 14504 14532
rect 14568 14504 14964 14532
rect 10410 14424 10416 14476
rect 10468 14424 10474 14476
rect 11054 14424 11060 14476
rect 11112 14464 11118 14476
rect 12250 14464 12256 14476
rect 11112 14436 12256 14464
rect 11112 14424 11118 14436
rect 12250 14424 12256 14436
rect 12308 14424 12314 14476
rect 12360 14473 12388 14504
rect 12345 14467 12403 14473
rect 12345 14433 12357 14467
rect 12391 14433 12403 14467
rect 12345 14427 12403 14433
rect 12529 14467 12587 14473
rect 12529 14433 12541 14467
rect 12575 14464 12587 14467
rect 12710 14464 12716 14476
rect 12575 14436 12716 14464
rect 12575 14433 12587 14436
rect 12529 14427 12587 14433
rect 12710 14424 12716 14436
rect 12768 14424 12774 14476
rect 14476 14464 14504 14504
rect 15010 14492 15016 14544
rect 15068 14532 15074 14544
rect 15580 14532 15608 14572
rect 15657 14569 15669 14603
rect 15703 14600 15715 14603
rect 16114 14600 16120 14612
rect 15703 14572 16120 14600
rect 15703 14569 15715 14572
rect 15657 14563 15715 14569
rect 16114 14560 16120 14572
rect 16172 14560 16178 14612
rect 16390 14560 16396 14612
rect 16448 14600 16454 14612
rect 20809 14603 20867 14609
rect 16448 14572 20392 14600
rect 16448 14560 16454 14572
rect 20364 14532 20392 14572
rect 20809 14569 20821 14603
rect 20855 14600 20867 14603
rect 20898 14600 20904 14612
rect 20855 14572 20904 14600
rect 20855 14569 20867 14572
rect 20809 14563 20867 14569
rect 20898 14560 20904 14572
rect 20956 14560 20962 14612
rect 21637 14603 21695 14609
rect 21637 14569 21649 14603
rect 21683 14600 21695 14603
rect 21726 14600 21732 14612
rect 21683 14572 21732 14600
rect 21683 14569 21695 14572
rect 21637 14563 21695 14569
rect 21726 14560 21732 14572
rect 21784 14560 21790 14612
rect 22002 14560 22008 14612
rect 22060 14600 22066 14612
rect 24486 14600 24492 14612
rect 22060 14572 24492 14600
rect 22060 14560 22066 14572
rect 24486 14560 24492 14572
rect 24544 14560 24550 14612
rect 25222 14560 25228 14612
rect 25280 14560 25286 14612
rect 26142 14560 26148 14612
rect 26200 14600 26206 14612
rect 26237 14603 26295 14609
rect 26237 14600 26249 14603
rect 26200 14572 26249 14600
rect 26200 14560 26206 14572
rect 26237 14569 26249 14572
rect 26283 14569 26295 14603
rect 26237 14563 26295 14569
rect 26973 14603 27031 14609
rect 26973 14569 26985 14603
rect 27019 14600 27031 14603
rect 27062 14600 27068 14612
rect 27019 14572 27068 14600
rect 27019 14569 27031 14572
rect 26973 14563 27031 14569
rect 27062 14560 27068 14572
rect 27120 14560 27126 14612
rect 27890 14560 27896 14612
rect 27948 14560 27954 14612
rect 29181 14603 29239 14609
rect 29181 14600 29193 14603
rect 28368 14572 29193 14600
rect 22462 14532 22468 14544
rect 15068 14504 15148 14532
rect 15580 14504 16068 14532
rect 20364 14504 22468 14532
rect 15068 14492 15074 14504
rect 14550 14464 14556 14476
rect 14476 14436 14556 14464
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 15120 14473 15148 14504
rect 15105 14467 15163 14473
rect 15105 14433 15117 14467
rect 15151 14433 15163 14467
rect 15105 14427 15163 14433
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14464 15347 14467
rect 15335 14436 15792 14464
rect 15335 14433 15347 14436
rect 15289 14427 15347 14433
rect 5353 14399 5411 14405
rect 5353 14365 5365 14399
rect 5399 14365 5411 14399
rect 5353 14359 5411 14365
rect 5368 14260 5396 14359
rect 7742 14356 7748 14408
rect 7800 14396 7806 14408
rect 10781 14399 10839 14405
rect 10781 14396 10793 14399
rect 7800 14368 10793 14396
rect 7800 14356 7806 14368
rect 10781 14365 10793 14368
rect 10827 14365 10839 14399
rect 10781 14359 10839 14365
rect 10874 14399 10932 14405
rect 10874 14365 10886 14399
rect 10920 14365 10932 14399
rect 10874 14359 10932 14365
rect 5620 14331 5678 14337
rect 5620 14297 5632 14331
rect 5666 14328 5678 14331
rect 6362 14328 6368 14340
rect 5666 14300 6368 14328
rect 5666 14297 5678 14300
rect 5620 14291 5678 14297
rect 6362 14288 6368 14300
rect 6420 14288 6426 14340
rect 9490 14288 9496 14340
rect 9548 14328 9554 14340
rect 10229 14331 10287 14337
rect 9548 14300 9996 14328
rect 9548 14288 9554 14300
rect 5534 14260 5540 14272
rect 5368 14232 5540 14260
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 6730 14220 6736 14272
rect 6788 14220 6794 14272
rect 9858 14220 9864 14272
rect 9916 14220 9922 14272
rect 9968 14260 9996 14300
rect 10229 14297 10241 14331
rect 10275 14328 10287 14331
rect 10686 14328 10692 14340
rect 10275 14300 10692 14328
rect 10275 14297 10287 14300
rect 10229 14291 10287 14297
rect 10686 14288 10692 14300
rect 10744 14328 10750 14340
rect 10888 14328 10916 14359
rect 11072 14337 11100 14424
rect 11287 14399 11345 14405
rect 11287 14365 11299 14399
rect 11333 14365 11345 14399
rect 11287 14359 11345 14365
rect 10744 14300 10916 14328
rect 11057 14331 11115 14337
rect 10744 14288 10750 14300
rect 11057 14297 11069 14331
rect 11103 14297 11115 14331
rect 11057 14291 11115 14297
rect 10321 14263 10379 14269
rect 10321 14260 10333 14263
rect 9968 14232 10333 14260
rect 10321 14229 10333 14232
rect 10367 14229 10379 14263
rect 10321 14223 10379 14229
rect 10778 14220 10784 14272
rect 10836 14260 10842 14272
rect 11072 14260 11100 14291
rect 11146 14288 11152 14340
rect 11204 14288 11210 14340
rect 11302 14328 11330 14359
rect 11974 14356 11980 14408
rect 12032 14396 12038 14408
rect 12069 14399 12127 14405
rect 12069 14396 12081 14399
rect 12032 14368 12081 14396
rect 12032 14356 12038 14368
rect 12069 14365 12081 14368
rect 12115 14365 12127 14399
rect 15013 14399 15071 14405
rect 12069 14359 12127 14365
rect 12176 14368 12940 14396
rect 12176 14328 12204 14368
rect 12805 14331 12863 14337
rect 12805 14328 12817 14331
rect 11302 14300 12204 14328
rect 12636 14300 12817 14328
rect 10836 14232 11100 14260
rect 11425 14263 11483 14269
rect 10836 14220 10842 14232
rect 11425 14229 11437 14263
rect 11471 14260 11483 14263
rect 12250 14260 12256 14272
rect 11471 14232 12256 14260
rect 11471 14229 11483 14232
rect 11425 14223 11483 14229
rect 12250 14220 12256 14232
rect 12308 14220 12314 14272
rect 12342 14220 12348 14272
rect 12400 14260 12406 14272
rect 12636 14260 12664 14300
rect 12805 14297 12817 14300
rect 12851 14297 12863 14331
rect 12805 14291 12863 14297
rect 12400 14232 12664 14260
rect 12713 14263 12771 14269
rect 12400 14220 12406 14232
rect 12713 14229 12725 14263
rect 12759 14260 12771 14263
rect 12912 14260 12940 14368
rect 15013 14365 15025 14399
rect 15059 14396 15071 14399
rect 15654 14396 15660 14408
rect 15059 14368 15660 14396
rect 15059 14365 15071 14368
rect 15013 14359 15071 14365
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 15565 14331 15623 14337
rect 15565 14297 15577 14331
rect 15611 14328 15623 14331
rect 15764 14328 15792 14436
rect 16040 14396 16068 14504
rect 22462 14492 22468 14504
rect 22520 14492 22526 14544
rect 24213 14535 24271 14541
rect 24213 14501 24225 14535
rect 24259 14501 24271 14535
rect 24213 14495 24271 14501
rect 17037 14467 17095 14473
rect 17037 14433 17049 14467
rect 17083 14464 17095 14467
rect 17494 14464 17500 14476
rect 17083 14436 17500 14464
rect 17083 14433 17095 14436
rect 17037 14427 17095 14433
rect 17494 14424 17500 14436
rect 17552 14424 17558 14476
rect 16040 14368 16712 14396
rect 16684 14328 16712 14368
rect 16758 14356 16764 14408
rect 16816 14405 16822 14408
rect 16816 14396 16828 14405
rect 16816 14368 16861 14396
rect 16816 14359 16828 14368
rect 16816 14356 16822 14359
rect 19426 14356 19432 14408
rect 19484 14356 19490 14408
rect 19696 14399 19754 14405
rect 19696 14365 19708 14399
rect 19742 14396 19754 14399
rect 19978 14396 19984 14408
rect 19742 14368 19984 14396
rect 19742 14365 19754 14368
rect 19696 14359 19754 14365
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 22370 14356 22376 14408
rect 22428 14396 22434 14408
rect 22833 14399 22891 14405
rect 22833 14396 22845 14399
rect 22428 14368 22845 14396
rect 22428 14356 22434 14368
rect 22833 14365 22845 14368
rect 22879 14365 22891 14399
rect 24228 14396 24256 14495
rect 24762 14492 24768 14544
rect 24820 14492 24826 14544
rect 25700 14504 27476 14532
rect 24578 14424 24584 14476
rect 24636 14464 24642 14476
rect 24780 14464 24808 14492
rect 25700 14473 25728 14504
rect 27448 14476 27476 14504
rect 24949 14467 25007 14473
rect 24949 14464 24961 14467
rect 24636 14436 24961 14464
rect 24636 14424 24642 14436
rect 24949 14433 24961 14436
rect 24995 14433 25007 14467
rect 24949 14427 25007 14433
rect 25685 14467 25743 14473
rect 25685 14433 25697 14467
rect 25731 14433 25743 14467
rect 25685 14427 25743 14433
rect 25869 14467 25927 14473
rect 25869 14433 25881 14467
rect 25915 14464 25927 14467
rect 26142 14464 26148 14476
rect 25915 14436 26148 14464
rect 25915 14433 25927 14436
rect 25869 14427 25927 14433
rect 26142 14424 26148 14436
rect 26200 14424 26206 14476
rect 27430 14424 27436 14476
rect 27488 14424 27494 14476
rect 27617 14467 27675 14473
rect 27617 14433 27629 14467
rect 27663 14464 27675 14467
rect 27908 14464 27936 14560
rect 27663 14436 28111 14464
rect 27663 14433 27675 14436
rect 27617 14427 27675 14433
rect 24670 14396 24676 14408
rect 24228 14368 24676 14396
rect 22833 14359 22891 14365
rect 24670 14356 24676 14368
rect 24728 14396 24734 14408
rect 24765 14399 24823 14405
rect 24765 14396 24777 14399
rect 24728 14368 24777 14396
rect 24728 14356 24734 14368
rect 24765 14365 24777 14368
rect 24811 14365 24823 14399
rect 24765 14359 24823 14365
rect 25593 14399 25651 14405
rect 25593 14365 25605 14399
rect 25639 14396 25651 14399
rect 26234 14396 26240 14408
rect 25639 14368 26240 14396
rect 25639 14365 25651 14368
rect 25593 14359 25651 14365
rect 26234 14356 26240 14368
rect 26292 14356 26298 14408
rect 27341 14399 27399 14405
rect 27341 14365 27353 14399
rect 27387 14396 27399 14399
rect 27982 14396 27988 14408
rect 27387 14368 27988 14396
rect 27387 14365 27399 14368
rect 27341 14359 27399 14365
rect 27982 14356 27988 14368
rect 28040 14356 28046 14408
rect 20898 14328 20904 14340
rect 15611 14300 16620 14328
rect 16684 14300 20904 14328
rect 15611 14297 15623 14300
rect 15565 14291 15623 14297
rect 13078 14260 13084 14272
rect 12759 14232 13084 14260
rect 12759 14229 12771 14232
rect 12713 14223 12771 14229
rect 13078 14220 13084 14232
rect 13136 14220 13142 14272
rect 16592 14260 16620 14300
rect 20898 14288 20904 14300
rect 20956 14288 20962 14340
rect 23100 14331 23158 14337
rect 23100 14297 23112 14331
rect 23146 14328 23158 14331
rect 23146 14300 24440 14328
rect 23146 14297 23158 14300
rect 23100 14291 23158 14297
rect 16666 14260 16672 14272
rect 16592 14232 16672 14260
rect 16666 14220 16672 14232
rect 16724 14220 16730 14272
rect 20622 14220 20628 14272
rect 20680 14260 20686 14272
rect 21082 14260 21088 14272
rect 20680 14232 21088 14260
rect 20680 14220 20686 14232
rect 21082 14220 21088 14232
rect 21140 14260 21146 14272
rect 21729 14263 21787 14269
rect 21729 14260 21741 14263
rect 21140 14232 21741 14260
rect 21140 14220 21146 14232
rect 21729 14229 21741 14232
rect 21775 14260 21787 14263
rect 24118 14260 24124 14272
rect 21775 14232 24124 14260
rect 21775 14229 21787 14232
rect 21729 14223 21787 14229
rect 24118 14220 24124 14232
rect 24176 14220 24182 14272
rect 24412 14269 24440 14300
rect 24397 14263 24455 14269
rect 24397 14229 24409 14263
rect 24443 14229 24455 14263
rect 24397 14223 24455 14229
rect 24486 14220 24492 14272
rect 24544 14260 24550 14272
rect 24857 14263 24915 14269
rect 24857 14260 24869 14263
rect 24544 14232 24869 14260
rect 24544 14220 24550 14232
rect 24857 14229 24869 14232
rect 24903 14229 24915 14263
rect 24857 14223 24915 14229
rect 24946 14220 24952 14272
rect 25004 14260 25010 14272
rect 25682 14260 25688 14272
rect 25004 14232 25688 14260
rect 25004 14220 25010 14232
rect 25682 14220 25688 14232
rect 25740 14220 25746 14272
rect 26142 14220 26148 14272
rect 26200 14220 26206 14272
rect 27982 14220 27988 14272
rect 28040 14260 28046 14272
rect 28083 14260 28111 14436
rect 28258 14424 28264 14476
rect 28316 14464 28322 14476
rect 28368 14464 28396 14572
rect 29181 14569 29193 14572
rect 29227 14600 29239 14603
rect 29733 14603 29791 14609
rect 29733 14600 29745 14603
rect 29227 14572 29745 14600
rect 29227 14569 29239 14572
rect 29181 14563 29239 14569
rect 29733 14569 29745 14572
rect 29779 14600 29791 14603
rect 30929 14603 30987 14609
rect 30929 14600 30941 14603
rect 29779 14572 30941 14600
rect 29779 14569 29791 14572
rect 29733 14563 29791 14569
rect 30929 14569 30941 14572
rect 30975 14569 30987 14603
rect 30929 14563 30987 14569
rect 32030 14560 32036 14612
rect 32088 14600 32094 14612
rect 33781 14603 33839 14609
rect 33781 14600 33793 14603
rect 32088 14572 33793 14600
rect 32088 14560 32094 14572
rect 33781 14569 33793 14572
rect 33827 14569 33839 14603
rect 33781 14563 33839 14569
rect 28537 14535 28595 14541
rect 28537 14532 28549 14535
rect 28316 14436 28396 14464
rect 28316 14424 28322 14436
rect 28368 14405 28396 14436
rect 28460 14504 28549 14532
rect 28353 14399 28411 14405
rect 28353 14365 28365 14399
rect 28399 14365 28411 14399
rect 28353 14359 28411 14365
rect 28166 14288 28172 14340
rect 28224 14288 28230 14340
rect 28258 14288 28264 14340
rect 28316 14288 28322 14340
rect 28040 14232 28111 14260
rect 28368 14260 28396 14359
rect 28460 14328 28488 14504
rect 28537 14501 28549 14504
rect 28583 14501 28595 14535
rect 28537 14495 28595 14501
rect 28626 14492 28632 14544
rect 28684 14532 28690 14544
rect 29270 14532 29276 14544
rect 28684 14504 29276 14532
rect 28684 14492 28690 14504
rect 29270 14492 29276 14504
rect 29328 14532 29334 14544
rect 29549 14535 29607 14541
rect 29549 14532 29561 14535
rect 29328 14504 29561 14532
rect 29328 14492 29334 14504
rect 29549 14501 29561 14504
rect 29595 14501 29607 14535
rect 30834 14532 30840 14544
rect 29549 14495 29607 14501
rect 30484 14504 30840 14532
rect 28718 14424 28724 14476
rect 28776 14464 28782 14476
rect 30282 14464 30288 14476
rect 28776 14436 30288 14464
rect 28776 14424 28782 14436
rect 30282 14424 30288 14436
rect 30340 14424 30346 14476
rect 30484 14473 30512 14504
rect 30834 14492 30840 14504
rect 30892 14492 30898 14544
rect 30469 14467 30527 14473
rect 30469 14433 30481 14467
rect 30515 14433 30527 14467
rect 30469 14427 30527 14433
rect 30558 14424 30564 14476
rect 30616 14464 30622 14476
rect 31021 14467 31079 14473
rect 31021 14464 31033 14467
rect 30616 14436 31033 14464
rect 30616 14424 30622 14436
rect 31021 14433 31033 14436
rect 31067 14433 31079 14467
rect 31021 14427 31079 14433
rect 28626 14356 28632 14408
rect 28684 14405 28690 14408
rect 28684 14396 28693 14405
rect 28684 14368 28729 14396
rect 28684 14359 28693 14368
rect 28684 14356 28690 14359
rect 28810 14356 28816 14408
rect 28868 14396 28874 14408
rect 28997 14399 29055 14405
rect 28997 14396 29009 14399
rect 28868 14368 29009 14396
rect 28868 14356 28874 14368
rect 28997 14365 29009 14368
rect 29043 14396 29055 14399
rect 29270 14396 29276 14408
rect 29043 14368 29276 14396
rect 29043 14365 29055 14368
rect 28997 14359 29055 14365
rect 29270 14356 29276 14368
rect 29328 14356 29334 14408
rect 29454 14356 29460 14408
rect 29512 14396 29518 14408
rect 30377 14399 30435 14405
rect 30377 14396 30389 14399
rect 29512 14368 30389 14396
rect 29512 14356 29518 14368
rect 30377 14365 30389 14368
rect 30423 14396 30435 14399
rect 31110 14396 31116 14408
rect 30423 14368 31116 14396
rect 30423 14365 30435 14368
rect 30377 14359 30435 14365
rect 31110 14356 31116 14368
rect 31168 14356 31174 14408
rect 33796 14396 33824 14563
rect 33962 14560 33968 14612
rect 34020 14560 34026 14612
rect 34149 14399 34207 14405
rect 34149 14396 34161 14399
rect 33796 14368 34161 14396
rect 34149 14365 34161 14368
rect 34195 14365 34207 14399
rect 34149 14359 34207 14365
rect 34422 14356 34428 14408
rect 34480 14356 34486 14408
rect 28902 14328 28908 14340
rect 28460 14300 28908 14328
rect 28902 14288 28908 14300
rect 28960 14288 28966 14340
rect 34333 14331 34391 14337
rect 34333 14297 34345 14331
rect 34379 14328 34391 14331
rect 34790 14328 34796 14340
rect 34379 14300 34796 14328
rect 34379 14297 34391 14300
rect 34333 14291 34391 14297
rect 34790 14288 34796 14300
rect 34848 14288 34854 14340
rect 28718 14260 28724 14272
rect 28368 14232 28724 14260
rect 28040 14220 28046 14232
rect 28718 14220 28724 14232
rect 28776 14220 28782 14272
rect 28810 14220 28816 14272
rect 28868 14220 28874 14272
rect 30006 14220 30012 14272
rect 30064 14220 30070 14272
rect 1104 14170 35328 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35328 14170
rect 1104 14096 35328 14118
rect 4893 14059 4951 14065
rect 4893 14025 4905 14059
rect 4939 14056 4951 14059
rect 6270 14056 6276 14068
rect 4939 14028 6276 14056
rect 4939 14025 4951 14028
rect 4893 14019 4951 14025
rect 6270 14016 6276 14028
rect 6328 14016 6334 14068
rect 6362 14016 6368 14068
rect 6420 14016 6426 14068
rect 6730 14016 6736 14068
rect 6788 14016 6794 14068
rect 7742 14016 7748 14068
rect 7800 14016 7806 14068
rect 8113 14059 8171 14065
rect 8113 14025 8125 14059
rect 8159 14056 8171 14059
rect 8386 14056 8392 14068
rect 8159 14028 8392 14056
rect 8159 14025 8171 14028
rect 8113 14019 8171 14025
rect 4525 13991 4583 13997
rect 4525 13957 4537 13991
rect 4571 13988 4583 13991
rect 5077 13991 5135 13997
rect 5077 13988 5089 13991
rect 4571 13960 5089 13988
rect 4571 13957 4583 13960
rect 4525 13951 4583 13957
rect 5077 13957 5089 13960
rect 5123 13988 5135 13991
rect 5442 13988 5448 14000
rect 5123 13960 5448 13988
rect 5123 13957 5135 13960
rect 5077 13951 5135 13957
rect 5442 13948 5448 13960
rect 5500 13948 5506 14000
rect 2866 13880 2872 13932
rect 2924 13920 2930 13932
rect 3418 13920 3424 13932
rect 2924 13892 3424 13920
rect 2924 13880 2930 13892
rect 3418 13880 3424 13892
rect 3476 13880 3482 13932
rect 4154 13880 4160 13932
rect 4212 13920 4218 13932
rect 4341 13923 4399 13929
rect 4341 13920 4353 13923
rect 4212 13892 4353 13920
rect 4212 13880 4218 13892
rect 4341 13889 4353 13892
rect 4387 13889 4399 13923
rect 4341 13883 4399 13889
rect 4614 13880 4620 13932
rect 4672 13880 4678 13932
rect 4709 13923 4767 13929
rect 4709 13889 4721 13923
rect 4755 13920 4767 13923
rect 5258 13920 5264 13932
rect 4755 13892 5264 13920
rect 4755 13889 4767 13892
rect 4709 13883 4767 13889
rect 5258 13880 5264 13892
rect 5316 13880 5322 13932
rect 6748 13920 6776 14016
rect 6914 13948 6920 14000
rect 6972 13988 6978 14000
rect 7469 13991 7527 13997
rect 7469 13988 7481 13991
rect 6972 13960 7481 13988
rect 6972 13948 6978 13960
rect 7469 13957 7481 13960
rect 7515 13957 7527 13991
rect 7469 13951 7527 13957
rect 7650 13948 7656 14000
rect 7708 13988 7714 14000
rect 7837 13991 7895 13997
rect 7837 13988 7849 13991
rect 7708 13960 7849 13988
rect 7708 13948 7714 13960
rect 7837 13957 7849 13960
rect 7883 13957 7895 13991
rect 7837 13951 7895 13957
rect 7193 13923 7251 13929
rect 7193 13920 7205 13923
rect 6748 13892 7205 13920
rect 7193 13889 7205 13892
rect 7239 13889 7251 13923
rect 7193 13883 7251 13889
rect 7377 13923 7435 13929
rect 7377 13889 7389 13923
rect 7423 13889 7435 13923
rect 7377 13883 7435 13889
rect 7561 13923 7619 13929
rect 7561 13889 7573 13923
rect 7607 13920 7619 13923
rect 8128 13920 8156 14019
rect 8386 14016 8392 14028
rect 8444 14056 8450 14068
rect 8754 14056 8760 14068
rect 8444 14028 8760 14056
rect 8444 14016 8450 14028
rect 8754 14016 8760 14028
rect 8812 14016 8818 14068
rect 10686 14016 10692 14068
rect 10744 14016 10750 14068
rect 11146 14016 11152 14068
rect 11204 14056 11210 14068
rect 11882 14056 11888 14068
rect 11204 14028 11888 14056
rect 11204 14016 11210 14028
rect 11882 14016 11888 14028
rect 11940 14056 11946 14068
rect 11977 14059 12035 14065
rect 11977 14056 11989 14059
rect 11940 14028 11989 14056
rect 11940 14016 11946 14028
rect 11977 14025 11989 14028
rect 12023 14025 12035 14059
rect 11977 14019 12035 14025
rect 13262 14016 13268 14068
rect 13320 14056 13326 14068
rect 14461 14059 14519 14065
rect 14461 14056 14473 14059
rect 13320 14028 14473 14056
rect 13320 14016 13326 14028
rect 14461 14025 14473 14028
rect 14507 14025 14519 14059
rect 14461 14019 14519 14025
rect 14550 14016 14556 14068
rect 14608 14056 14614 14068
rect 16574 14056 16580 14068
rect 14608 14028 16580 14056
rect 14608 14016 14614 14028
rect 16574 14016 16580 14028
rect 16632 14016 16638 14068
rect 21269 14059 21327 14065
rect 21269 14056 21281 14059
rect 16684 14028 21281 14056
rect 9576 13991 9634 13997
rect 9576 13957 9588 13991
rect 9622 13988 9634 13991
rect 9858 13988 9864 14000
rect 9622 13960 9864 13988
rect 9622 13957 9634 13960
rect 9576 13951 9634 13957
rect 9858 13948 9864 13960
rect 9916 13948 9922 14000
rect 10410 13948 10416 14000
rect 10468 13988 10474 14000
rect 10781 13991 10839 13997
rect 10781 13988 10793 13991
rect 10468 13960 10793 13988
rect 10468 13948 10474 13960
rect 10781 13957 10793 13960
rect 10827 13957 10839 13991
rect 10781 13951 10839 13957
rect 13998 13948 14004 14000
rect 14056 13988 14062 14000
rect 16684 13988 16712 14028
rect 21269 14025 21281 14028
rect 21315 14025 21327 14059
rect 21269 14019 21327 14025
rect 23845 14059 23903 14065
rect 23845 14025 23857 14059
rect 23891 14025 23903 14059
rect 23845 14019 23903 14025
rect 14056 13960 16712 13988
rect 16776 13960 17540 13988
rect 14056 13948 14062 13960
rect 7607 13892 8156 13920
rect 7607 13889 7619 13892
rect 7561 13883 7619 13889
rect 6825 13855 6883 13861
rect 6825 13821 6837 13855
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 6840 13728 6868 13815
rect 7006 13812 7012 13864
rect 7064 13812 7070 13864
rect 7392 13852 7420 13883
rect 9306 13880 9312 13932
rect 9364 13880 9370 13932
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 11974 13920 11980 13932
rect 11931 13892 11980 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 11974 13880 11980 13892
rect 12032 13880 12038 13932
rect 12345 13923 12403 13929
rect 12345 13889 12357 13923
rect 12391 13920 12403 13923
rect 12434 13920 12440 13932
rect 12391 13892 12440 13920
rect 12391 13889 12403 13892
rect 12345 13883 12403 13889
rect 12434 13880 12440 13892
rect 12492 13880 12498 13932
rect 12618 13929 12624 13932
rect 12612 13883 12624 13929
rect 12618 13880 12624 13883
rect 12676 13880 12682 13932
rect 12986 13880 12992 13932
rect 13044 13920 13050 13932
rect 13817 13923 13875 13929
rect 13817 13920 13829 13923
rect 13044 13892 13829 13920
rect 13044 13880 13050 13892
rect 13817 13889 13829 13892
rect 13863 13889 13875 13923
rect 13817 13883 13875 13889
rect 13910 13923 13968 13929
rect 13910 13889 13922 13923
rect 13956 13889 13968 13923
rect 13910 13883 13968 13889
rect 7650 13852 7656 13864
rect 7392 13824 7656 13852
rect 7650 13812 7656 13824
rect 7708 13812 7714 13864
rect 12161 13855 12219 13861
rect 12161 13821 12173 13855
rect 12207 13821 12219 13855
rect 13924 13852 13952 13883
rect 14090 13880 14096 13932
rect 14148 13880 14154 13932
rect 14182 13880 14188 13932
rect 14240 13880 14246 13932
rect 14274 13880 14280 13932
rect 14332 13929 14338 13932
rect 14332 13923 14381 13929
rect 14332 13889 14335 13923
rect 14369 13920 14381 13923
rect 14369 13892 14872 13920
rect 14369 13889 14381 13892
rect 14332 13883 14381 13889
rect 14332 13880 14338 13883
rect 12161 13815 12219 13821
rect 13740 13824 13952 13852
rect 14108 13852 14136 13880
rect 14642 13852 14648 13864
rect 14108 13824 14648 13852
rect 3605 13719 3663 13725
rect 3605 13685 3617 13719
rect 3651 13716 3663 13719
rect 3694 13716 3700 13728
rect 3651 13688 3700 13716
rect 3651 13685 3663 13688
rect 3605 13679 3663 13685
rect 3694 13676 3700 13688
rect 3752 13676 3758 13728
rect 6822 13676 6828 13728
rect 6880 13716 6886 13728
rect 9490 13716 9496 13728
rect 6880 13688 9496 13716
rect 6880 13676 6886 13688
rect 9490 13676 9496 13688
rect 9548 13676 9554 13728
rect 11514 13676 11520 13728
rect 11572 13676 11578 13728
rect 12176 13716 12204 13815
rect 13740 13728 13768 13824
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 14844 13861 14872 13892
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 16776 13929 16804 13960
rect 17512 13932 17540 13960
rect 16761 13923 16819 13929
rect 16761 13920 16773 13923
rect 15160 13892 16773 13920
rect 15160 13880 15166 13892
rect 16761 13889 16773 13892
rect 16807 13889 16819 13923
rect 16761 13883 16819 13889
rect 17028 13923 17086 13929
rect 17028 13889 17040 13923
rect 17074 13920 17086 13923
rect 17310 13920 17316 13932
rect 17074 13892 17316 13920
rect 17074 13889 17086 13892
rect 17028 13883 17086 13889
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 17494 13880 17500 13932
rect 17552 13920 17558 13932
rect 18325 13923 18383 13929
rect 18325 13920 18337 13923
rect 17552 13892 18337 13920
rect 17552 13880 17558 13892
rect 18325 13889 18337 13892
rect 18371 13889 18383 13923
rect 18325 13883 18383 13889
rect 18592 13923 18650 13929
rect 18592 13889 18604 13923
rect 18638 13920 18650 13923
rect 19150 13920 19156 13932
rect 18638 13892 19156 13920
rect 18638 13889 18650 13892
rect 18592 13883 18650 13889
rect 19150 13880 19156 13892
rect 19208 13880 19214 13932
rect 21284 13920 21312 14019
rect 22640 13991 22698 13997
rect 22640 13957 22652 13991
rect 22686 13988 22698 13991
rect 23860 13988 23888 14019
rect 24118 14016 24124 14068
rect 24176 14056 24182 14068
rect 24854 14056 24860 14068
rect 24176 14028 24860 14056
rect 24176 14016 24182 14028
rect 24854 14016 24860 14028
rect 24912 14016 24918 14068
rect 25225 14059 25283 14065
rect 25225 14025 25237 14059
rect 25271 14056 25283 14059
rect 26418 14056 26424 14068
rect 25271 14028 26424 14056
rect 25271 14025 25283 14028
rect 25225 14019 25283 14025
rect 26418 14016 26424 14028
rect 26476 14016 26482 14068
rect 27062 14016 27068 14068
rect 27120 14016 27126 14068
rect 27890 14016 27896 14068
rect 27948 14056 27954 14068
rect 27985 14059 28043 14065
rect 27985 14056 27997 14059
rect 27948 14028 27997 14056
rect 27948 14016 27954 14028
rect 27985 14025 27997 14028
rect 28031 14025 28043 14059
rect 27985 14019 28043 14025
rect 28258 14016 28264 14068
rect 28316 14056 28322 14068
rect 28810 14056 28816 14068
rect 28316 14028 28816 14056
rect 28316 14016 28322 14028
rect 28810 14016 28816 14028
rect 28868 14056 28874 14068
rect 29549 14059 29607 14065
rect 29549 14056 29561 14059
rect 28868 14028 29561 14056
rect 28868 14016 28874 14028
rect 29549 14025 29561 14028
rect 29595 14025 29607 14059
rect 29549 14019 29607 14025
rect 31110 14016 31116 14068
rect 31168 14016 31174 14068
rect 22686 13960 23888 13988
rect 24213 13991 24271 13997
rect 22686 13957 22698 13960
rect 22640 13951 22698 13957
rect 24213 13957 24225 13991
rect 24259 13988 24271 13991
rect 24949 13991 25007 13997
rect 24949 13988 24961 13991
rect 24259 13960 24961 13988
rect 24259 13957 24271 13960
rect 24213 13951 24271 13957
rect 24949 13957 24961 13960
rect 24995 13957 25007 13991
rect 24949 13951 25007 13957
rect 21453 13923 21511 13929
rect 21453 13920 21465 13923
rect 21284 13892 21465 13920
rect 21453 13889 21465 13892
rect 21499 13889 21511 13923
rect 21453 13883 21511 13889
rect 22097 13923 22155 13929
rect 22097 13889 22109 13923
rect 22143 13920 22155 13923
rect 22278 13920 22284 13932
rect 22143 13892 22284 13920
rect 22143 13889 22155 13892
rect 22097 13883 22155 13889
rect 22278 13880 22284 13892
rect 22336 13880 22342 13932
rect 14829 13855 14887 13861
rect 14829 13821 14841 13855
rect 14875 13852 14887 13855
rect 15010 13852 15016 13864
rect 14875 13824 15016 13852
rect 14875 13821 14887 13824
rect 14829 13815 14887 13821
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 22370 13812 22376 13864
rect 22428 13812 22434 13864
rect 24228 13852 24256 13951
rect 25406 13948 25412 14000
rect 25464 13988 25470 14000
rect 25961 13991 26019 13997
rect 25961 13988 25973 13991
rect 25464 13960 25973 13988
rect 25464 13948 25470 13960
rect 25961 13957 25973 13960
rect 26007 13957 26019 13991
rect 25961 13951 26019 13957
rect 26142 13948 26148 14000
rect 26200 13988 26206 14000
rect 26329 13991 26387 13997
rect 26329 13988 26341 13991
rect 26200 13960 26341 13988
rect 26200 13948 26206 13960
rect 26329 13957 26341 13960
rect 26375 13988 26387 13991
rect 27080 13988 27108 14016
rect 28442 13997 28448 14000
rect 26375 13960 27108 13988
rect 26375 13957 26387 13960
rect 26329 13951 26387 13957
rect 28436 13951 28448 13997
rect 28442 13948 28448 13951
rect 28500 13948 28506 14000
rect 32122 13988 32128 14000
rect 29748 13960 32128 13988
rect 24670 13880 24676 13932
rect 24728 13880 24734 13932
rect 24854 13880 24860 13932
rect 24912 13880 24918 13932
rect 25041 13923 25099 13929
rect 25041 13889 25053 13923
rect 25087 13889 25099 13923
rect 25041 13883 25099 13889
rect 25593 13923 25651 13929
rect 25593 13889 25605 13923
rect 25639 13920 25651 13923
rect 26050 13920 26056 13932
rect 25639 13892 26056 13920
rect 25639 13889 25651 13892
rect 25593 13883 25651 13889
rect 23768 13824 24256 13852
rect 24305 13855 24363 13861
rect 21637 13787 21695 13793
rect 17696 13756 18276 13784
rect 12710 13716 12716 13728
rect 12176 13688 12716 13716
rect 12710 13676 12716 13688
rect 12768 13716 12774 13728
rect 13538 13716 13544 13728
rect 12768 13688 13544 13716
rect 12768 13676 12774 13688
rect 13538 13676 13544 13688
rect 13596 13676 13602 13728
rect 13722 13676 13728 13728
rect 13780 13676 13786 13728
rect 16482 13676 16488 13728
rect 16540 13716 16546 13728
rect 17696 13716 17724 13756
rect 16540 13688 17724 13716
rect 16540 13676 16546 13688
rect 17954 13676 17960 13728
rect 18012 13716 18018 13728
rect 18141 13719 18199 13725
rect 18141 13716 18153 13719
rect 18012 13688 18153 13716
rect 18012 13676 18018 13688
rect 18141 13685 18153 13688
rect 18187 13685 18199 13719
rect 18248 13716 18276 13756
rect 21637 13753 21649 13787
rect 21683 13784 21695 13787
rect 21726 13784 21732 13796
rect 21683 13756 21732 13784
rect 21683 13753 21695 13756
rect 21637 13747 21695 13753
rect 21726 13744 21732 13756
rect 21784 13784 21790 13796
rect 23768 13793 23796 13824
rect 24305 13821 24317 13855
rect 24351 13821 24363 13855
rect 24305 13815 24363 13821
rect 23753 13787 23811 13793
rect 21784 13756 22416 13784
rect 21784 13744 21790 13756
rect 18690 13716 18696 13728
rect 18248 13688 18696 13716
rect 18141 13679 18199 13685
rect 18690 13676 18696 13688
rect 18748 13676 18754 13728
rect 19702 13676 19708 13728
rect 19760 13676 19766 13728
rect 21913 13719 21971 13725
rect 21913 13685 21925 13719
rect 21959 13716 21971 13719
rect 22094 13716 22100 13728
rect 21959 13688 22100 13716
rect 21959 13685 21971 13688
rect 21913 13679 21971 13685
rect 22094 13676 22100 13688
rect 22152 13716 22158 13728
rect 22189 13719 22247 13725
rect 22189 13716 22201 13719
rect 22152 13688 22201 13716
rect 22152 13676 22158 13688
rect 22189 13685 22201 13688
rect 22235 13685 22247 13719
rect 22388 13716 22416 13756
rect 23753 13753 23765 13787
rect 23799 13753 23811 13787
rect 24320 13784 24348 13815
rect 24394 13812 24400 13864
rect 24452 13812 24458 13864
rect 24762 13812 24768 13864
rect 24820 13852 24826 13864
rect 25056 13852 25084 13883
rect 26050 13880 26056 13892
rect 26108 13880 26114 13932
rect 26970 13880 26976 13932
rect 27028 13920 27034 13932
rect 27798 13920 27804 13932
rect 27028 13892 27804 13920
rect 27028 13880 27034 13892
rect 27798 13880 27804 13892
rect 27856 13920 27862 13932
rect 28169 13923 28227 13929
rect 28169 13920 28181 13923
rect 27856 13892 28181 13920
rect 27856 13880 27862 13892
rect 28169 13889 28181 13892
rect 28215 13889 28227 13923
rect 29546 13920 29552 13932
rect 28169 13883 28227 13889
rect 28276 13892 29552 13920
rect 26421 13855 26479 13861
rect 26421 13852 26433 13855
rect 24820 13824 26433 13852
rect 24820 13812 24826 13824
rect 25424 13793 25452 13824
rect 26421 13821 26433 13824
rect 26467 13852 26479 13855
rect 26605 13855 26663 13861
rect 26605 13852 26617 13855
rect 26467 13824 26617 13852
rect 26467 13821 26479 13824
rect 26421 13815 26479 13821
rect 26605 13821 26617 13824
rect 26651 13821 26663 13855
rect 26605 13815 26663 13821
rect 27246 13812 27252 13864
rect 27304 13852 27310 13864
rect 28276 13852 28304 13892
rect 29546 13880 29552 13892
rect 29604 13880 29610 13932
rect 29748 13864 29776 13960
rect 32122 13948 32128 13960
rect 32180 13948 32186 14000
rect 30006 13929 30012 13932
rect 30000 13920 30012 13929
rect 29967 13892 30012 13920
rect 30000 13883 30012 13892
rect 30006 13880 30012 13883
rect 30064 13880 30070 13932
rect 27304 13824 28304 13852
rect 27304 13812 27310 13824
rect 29730 13812 29736 13864
rect 29788 13812 29794 13864
rect 23753 13747 23811 13753
rect 24228 13756 24348 13784
rect 25409 13787 25467 13793
rect 24228 13716 24256 13756
rect 25409 13753 25421 13787
rect 25455 13753 25467 13787
rect 26510 13784 26516 13796
rect 25409 13747 25467 13753
rect 25608 13756 26516 13784
rect 25608 13716 25636 13756
rect 26510 13744 26516 13756
rect 26568 13744 26574 13796
rect 22388 13688 25636 13716
rect 22189 13679 22247 13685
rect 25682 13676 25688 13728
rect 25740 13676 25746 13728
rect 1104 13626 35328 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 35328 13626
rect 1104 13552 35328 13574
rect 3605 13515 3663 13521
rect 3605 13481 3617 13515
rect 3651 13512 3663 13515
rect 4062 13512 4068 13524
rect 3651 13484 4068 13512
rect 3651 13481 3663 13484
rect 3605 13475 3663 13481
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 6914 13472 6920 13524
rect 6972 13472 6978 13524
rect 7006 13472 7012 13524
rect 7064 13512 7070 13524
rect 7285 13515 7343 13521
rect 7285 13512 7297 13515
rect 7064 13484 7297 13512
rect 7064 13472 7070 13484
rect 7285 13481 7297 13484
rect 7331 13512 7343 13515
rect 7331 13484 11468 13512
rect 7331 13481 7343 13484
rect 7285 13475 7343 13481
rect 11440 13444 11468 13484
rect 11882 13472 11888 13524
rect 11940 13472 11946 13524
rect 12250 13472 12256 13524
rect 12308 13472 12314 13524
rect 12618 13472 12624 13524
rect 12676 13512 12682 13524
rect 12805 13515 12863 13521
rect 12805 13512 12817 13515
rect 12676 13484 12817 13512
rect 12676 13472 12682 13484
rect 12805 13481 12817 13484
rect 12851 13481 12863 13515
rect 12805 13475 12863 13481
rect 14918 13472 14924 13524
rect 14976 13472 14982 13524
rect 17310 13472 17316 13524
rect 17368 13472 17374 13524
rect 19150 13472 19156 13524
rect 19208 13512 19214 13524
rect 19245 13515 19303 13521
rect 19245 13512 19257 13515
rect 19208 13484 19257 13512
rect 19208 13472 19214 13484
rect 19245 13481 19257 13484
rect 19291 13481 19303 13515
rect 23753 13515 23811 13521
rect 19245 13475 19303 13481
rect 19812 13484 22784 13512
rect 12710 13444 12716 13456
rect 11440 13416 12716 13444
rect 12710 13404 12716 13416
rect 12768 13404 12774 13456
rect 13170 13404 13176 13456
rect 13228 13444 13234 13456
rect 13630 13444 13636 13456
rect 13228 13416 13636 13444
rect 13228 13404 13234 13416
rect 5534 13336 5540 13388
rect 5592 13336 5598 13388
rect 9122 13336 9128 13388
rect 9180 13376 9186 13388
rect 9493 13379 9551 13385
rect 9493 13376 9505 13379
rect 9180 13348 9505 13376
rect 9180 13336 9186 13348
rect 9493 13345 9505 13348
rect 9539 13376 9551 13379
rect 9582 13376 9588 13388
rect 9539 13348 9588 13376
rect 9539 13345 9551 13348
rect 9493 13339 9551 13345
rect 9582 13336 9588 13348
rect 9640 13376 9646 13388
rect 9769 13379 9827 13385
rect 9769 13376 9781 13379
rect 9640 13348 9781 13376
rect 9640 13336 9646 13348
rect 9769 13345 9781 13348
rect 9815 13345 9827 13379
rect 9769 13339 9827 13345
rect 12345 13379 12403 13385
rect 12345 13345 12357 13379
rect 12391 13376 12403 13379
rect 13262 13376 13268 13388
rect 12391 13348 13268 13376
rect 12391 13345 12403 13348
rect 12345 13339 12403 13345
rect 13262 13336 13268 13348
rect 13320 13336 13326 13388
rect 13372 13385 13400 13416
rect 13630 13404 13636 13416
rect 13688 13404 13694 13456
rect 13357 13379 13415 13385
rect 13357 13345 13369 13379
rect 13403 13345 13415 13379
rect 13357 13339 13415 13345
rect 14182 13336 14188 13388
rect 14240 13376 14246 13388
rect 14553 13379 14611 13385
rect 14553 13376 14565 13379
rect 14240 13348 14565 13376
rect 14240 13336 14246 13348
rect 14553 13345 14565 13348
rect 14599 13345 14611 13379
rect 14553 13339 14611 13345
rect 14737 13379 14795 13385
rect 14737 13345 14749 13379
rect 14783 13376 14795 13379
rect 14826 13376 14832 13388
rect 14783 13348 14832 13376
rect 14783 13345 14795 13348
rect 14737 13339 14795 13345
rect 14826 13336 14832 13348
rect 14884 13376 14890 13388
rect 14936 13376 14964 13472
rect 17586 13404 17592 13456
rect 17644 13444 17650 13456
rect 17644 13416 18276 13444
rect 17644 13404 17650 13416
rect 14884 13348 14964 13376
rect 14884 13336 14890 13348
rect 15102 13336 15108 13388
rect 15160 13336 15166 13388
rect 17865 13379 17923 13385
rect 17865 13345 17877 13379
rect 17911 13376 17923 13379
rect 18141 13379 18199 13385
rect 18141 13376 18153 13379
rect 17911 13348 18153 13376
rect 17911 13345 17923 13348
rect 17865 13339 17923 13345
rect 18141 13345 18153 13348
rect 18187 13345 18199 13379
rect 18248 13376 18276 13416
rect 18506 13404 18512 13456
rect 18564 13444 18570 13456
rect 18877 13447 18935 13453
rect 18877 13444 18889 13447
rect 18564 13416 18889 13444
rect 18564 13404 18570 13416
rect 18877 13413 18889 13416
rect 18923 13444 18935 13447
rect 19812 13444 19840 13484
rect 18923 13416 19840 13444
rect 21821 13447 21879 13453
rect 18923 13413 18935 13416
rect 18877 13407 18935 13413
rect 21821 13413 21833 13447
rect 21867 13444 21879 13447
rect 22186 13444 22192 13456
rect 21867 13416 22192 13444
rect 21867 13413 21879 13416
rect 21821 13407 21879 13413
rect 22186 13404 22192 13416
rect 22244 13404 22250 13456
rect 22756 13444 22784 13484
rect 23753 13481 23765 13515
rect 23799 13512 23811 13515
rect 24394 13512 24400 13524
rect 23799 13484 24400 13512
rect 23799 13481 23811 13484
rect 23753 13475 23811 13481
rect 24394 13472 24400 13484
rect 24452 13472 24458 13524
rect 24489 13515 24547 13521
rect 24489 13481 24501 13515
rect 24535 13512 24547 13515
rect 24578 13512 24584 13524
rect 24535 13484 24584 13512
rect 24535 13481 24547 13484
rect 24489 13475 24547 13481
rect 24578 13472 24584 13484
rect 24636 13472 24642 13524
rect 26326 13512 26332 13524
rect 24964 13484 26332 13512
rect 24964 13444 24992 13484
rect 26326 13472 26332 13484
rect 26384 13512 26390 13524
rect 26384 13484 26740 13512
rect 26384 13472 26390 13484
rect 22756 13416 24992 13444
rect 26712 13444 26740 13484
rect 27246 13472 27252 13524
rect 27304 13472 27310 13524
rect 27522 13472 27528 13524
rect 27580 13512 27586 13524
rect 28261 13515 28319 13521
rect 28261 13512 28273 13515
rect 27580 13484 28273 13512
rect 27580 13472 27586 13484
rect 28261 13481 28273 13484
rect 28307 13481 28319 13515
rect 28261 13475 28319 13481
rect 26878 13444 26884 13456
rect 26712 13416 26884 13444
rect 19610 13376 19616 13388
rect 18248 13348 19616 13376
rect 18141 13339 18199 13345
rect 2225 13311 2283 13317
rect 2225 13277 2237 13311
rect 2271 13308 2283 13311
rect 2774 13308 2780 13320
rect 2271 13280 2780 13308
rect 2271 13277 2283 13280
rect 2225 13271 2283 13277
rect 2774 13268 2780 13280
rect 2832 13308 2838 13320
rect 3789 13311 3847 13317
rect 3789 13308 3801 13311
rect 2832 13280 3801 13308
rect 2832 13268 2838 13280
rect 3789 13277 3801 13280
rect 3835 13277 3847 13311
rect 5552 13308 5580 13336
rect 7377 13311 7435 13317
rect 7377 13308 7389 13311
rect 5552 13280 7389 13308
rect 3789 13271 3847 13277
rect 7377 13277 7389 13280
rect 7423 13277 7435 13311
rect 7377 13271 7435 13277
rect 9306 13268 9312 13320
rect 9364 13308 9370 13320
rect 10505 13311 10563 13317
rect 10505 13308 10517 13311
rect 9364 13280 10517 13308
rect 9364 13268 9370 13280
rect 10505 13277 10517 13280
rect 10551 13277 10563 13311
rect 10505 13271 10563 13277
rect 10772 13311 10830 13317
rect 10772 13277 10784 13311
rect 10818 13308 10830 13311
rect 11514 13308 11520 13320
rect 10818 13280 11520 13308
rect 10818 13277 10830 13280
rect 10772 13271 10830 13277
rect 11514 13268 11520 13280
rect 11572 13268 11578 13320
rect 12250 13268 12256 13320
rect 12308 13268 12314 13320
rect 13173 13311 13231 13317
rect 13173 13277 13185 13311
rect 13219 13308 13231 13311
rect 13722 13308 13728 13320
rect 13219 13280 13728 13308
rect 13219 13277 13231 13280
rect 13173 13271 13231 13277
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 13832 13280 14504 13308
rect 2492 13243 2550 13249
rect 2492 13209 2504 13243
rect 2538 13240 2550 13243
rect 2958 13240 2964 13252
rect 2538 13212 2964 13240
rect 2538 13209 2550 13212
rect 2492 13203 2550 13209
rect 2958 13200 2964 13212
rect 3016 13200 3022 13252
rect 4062 13249 4068 13252
rect 4056 13203 4068 13249
rect 4062 13200 4068 13203
rect 4120 13200 4126 13252
rect 5804 13243 5862 13249
rect 5804 13209 5816 13243
rect 5850 13240 5862 13243
rect 6362 13240 6368 13252
rect 5850 13212 6368 13240
rect 5850 13209 5862 13212
rect 5804 13203 5862 13209
rect 6362 13200 6368 13212
rect 6420 13200 6426 13252
rect 7644 13243 7702 13249
rect 7644 13209 7656 13243
rect 7690 13240 7702 13243
rect 9401 13243 9459 13249
rect 7690 13212 8984 13240
rect 7690 13209 7702 13212
rect 7644 13203 7702 13209
rect 4338 13132 4344 13184
rect 4396 13172 4402 13184
rect 4614 13172 4620 13184
rect 4396 13144 4620 13172
rect 4396 13132 4402 13144
rect 4614 13132 4620 13144
rect 4672 13172 4678 13184
rect 5169 13175 5227 13181
rect 5169 13172 5181 13175
rect 4672 13144 5181 13172
rect 4672 13132 4678 13144
rect 5169 13141 5181 13144
rect 5215 13141 5227 13175
rect 5169 13135 5227 13141
rect 8757 13175 8815 13181
rect 8757 13141 8769 13175
rect 8803 13172 8815 13175
rect 8846 13172 8852 13184
rect 8803 13144 8852 13172
rect 8803 13141 8815 13144
rect 8757 13135 8815 13141
rect 8846 13132 8852 13144
rect 8904 13132 8910 13184
rect 8956 13181 8984 13212
rect 9401 13209 9413 13243
rect 9447 13240 9459 13243
rect 9490 13240 9496 13252
rect 9447 13212 9496 13240
rect 9447 13209 9459 13212
rect 9401 13203 9459 13209
rect 9490 13200 9496 13212
rect 9548 13200 9554 13252
rect 11974 13200 11980 13252
rect 12032 13240 12038 13252
rect 12434 13240 12440 13252
rect 12032 13212 12440 13240
rect 12032 13200 12038 13212
rect 12434 13200 12440 13212
rect 12492 13240 12498 13252
rect 13265 13243 13323 13249
rect 13265 13240 13277 13243
rect 12492 13212 13277 13240
rect 12492 13200 12498 13212
rect 13265 13209 13277 13212
rect 13311 13240 13323 13243
rect 13832 13240 13860 13280
rect 13311 13212 13860 13240
rect 13311 13209 13323 13212
rect 13265 13203 13323 13209
rect 8941 13175 8999 13181
rect 8941 13141 8953 13175
rect 8987 13141 8999 13175
rect 8941 13135 8999 13141
rect 9030 13132 9036 13184
rect 9088 13172 9094 13184
rect 9309 13175 9367 13181
rect 9309 13172 9321 13175
rect 9088 13144 9321 13172
rect 9088 13132 9094 13144
rect 9309 13141 9321 13144
rect 9355 13141 9367 13175
rect 9309 13135 9367 13141
rect 12618 13132 12624 13184
rect 12676 13132 12682 13184
rect 12894 13132 12900 13184
rect 12952 13172 12958 13184
rect 13170 13172 13176 13184
rect 12952 13144 13176 13172
rect 12952 13132 12958 13144
rect 13170 13132 13176 13144
rect 13228 13132 13234 13184
rect 14090 13132 14096 13184
rect 14148 13132 14154 13184
rect 14476 13181 14504 13280
rect 16574 13268 16580 13320
rect 16632 13268 16638 13320
rect 17681 13311 17739 13317
rect 17681 13277 17693 13311
rect 17727 13308 17739 13311
rect 17954 13308 17960 13320
rect 17727 13280 17960 13308
rect 17727 13277 17739 13280
rect 17681 13271 17739 13277
rect 17954 13268 17960 13280
rect 18012 13268 18018 13320
rect 18156 13308 18184 13339
rect 19610 13336 19616 13348
rect 19668 13376 19674 13388
rect 19797 13379 19855 13385
rect 19797 13376 19809 13379
rect 19668 13348 19809 13376
rect 19668 13336 19674 13348
rect 19797 13345 19809 13348
rect 19843 13376 19855 13379
rect 20073 13379 20131 13385
rect 20073 13376 20085 13379
rect 19843 13348 20085 13376
rect 19843 13345 19855 13348
rect 19797 13339 19855 13345
rect 20073 13345 20085 13348
rect 20119 13345 20131 13379
rect 20073 13339 20131 13345
rect 22370 13336 22376 13388
rect 22428 13376 22434 13388
rect 22741 13379 22799 13385
rect 22741 13376 22753 13379
rect 22428 13348 22753 13376
rect 22428 13336 22434 13348
rect 22741 13345 22753 13348
rect 22787 13376 22799 13379
rect 24949 13379 25007 13385
rect 24949 13376 24961 13379
rect 22787 13348 24961 13376
rect 22787 13345 22799 13348
rect 22741 13339 22799 13345
rect 24949 13345 24961 13348
rect 24995 13345 25007 13379
rect 24949 13339 25007 13345
rect 18156 13280 19380 13308
rect 15372 13243 15430 13249
rect 15372 13209 15384 13243
rect 15418 13240 15430 13243
rect 15654 13240 15660 13252
rect 15418 13212 15660 13240
rect 15418 13209 15430 13212
rect 15372 13203 15430 13209
rect 15654 13200 15660 13212
rect 15712 13200 15718 13252
rect 19352 13240 19380 13280
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 20441 13311 20499 13317
rect 20441 13308 20453 13311
rect 19484 13280 20453 13308
rect 19484 13268 19490 13280
rect 20441 13277 20453 13280
rect 20487 13277 20499 13311
rect 20441 13271 20499 13277
rect 20990 13268 20996 13320
rect 21048 13308 21054 13320
rect 23842 13308 23848 13320
rect 21048 13280 23848 13308
rect 21048 13268 21054 13280
rect 23842 13268 23848 13280
rect 23900 13268 23906 13320
rect 26418 13268 26424 13320
rect 26476 13268 26482 13320
rect 26712 13317 26740 13416
rect 26878 13404 26884 13416
rect 26936 13404 26942 13456
rect 28276 13444 28304 13475
rect 28442 13472 28448 13524
rect 28500 13472 28506 13524
rect 29270 13472 29276 13524
rect 29328 13472 29334 13524
rect 30558 13444 30564 13456
rect 28276 13416 30564 13444
rect 30558 13404 30564 13416
rect 30616 13404 30622 13456
rect 27985 13379 28043 13385
rect 27985 13376 27997 13379
rect 27356 13348 27997 13376
rect 27356 13320 27384 13348
rect 27985 13345 27997 13348
rect 28031 13345 28043 13379
rect 27985 13339 28043 13345
rect 28074 13336 28080 13388
rect 28132 13376 28138 13388
rect 28905 13379 28963 13385
rect 28905 13376 28917 13379
rect 28132 13348 28917 13376
rect 28132 13336 28138 13348
rect 28905 13345 28917 13348
rect 28951 13345 28963 13379
rect 28905 13339 28963 13345
rect 28997 13379 29055 13385
rect 28997 13345 29009 13379
rect 29043 13345 29055 13379
rect 28997 13339 29055 13345
rect 26514 13311 26572 13317
rect 26514 13277 26526 13311
rect 26560 13277 26572 13311
rect 26514 13271 26572 13277
rect 26697 13311 26755 13317
rect 26697 13277 26709 13311
rect 26743 13277 26755 13311
rect 26697 13271 26755 13277
rect 26927 13311 26985 13317
rect 26927 13277 26939 13311
rect 26973 13308 26985 13311
rect 27246 13308 27252 13320
rect 26973 13280 27252 13308
rect 26973 13277 26985 13280
rect 26927 13271 26985 13277
rect 20530 13240 20536 13252
rect 15764 13212 17899 13240
rect 19352 13212 20536 13240
rect 14461 13175 14519 13181
rect 14461 13141 14473 13175
rect 14507 13172 14519 13175
rect 15764 13172 15792 13212
rect 14507 13144 15792 13172
rect 14507 13141 14519 13144
rect 14461 13135 14519 13141
rect 16022 13132 16028 13184
rect 16080 13172 16086 13184
rect 16485 13175 16543 13181
rect 16485 13172 16497 13175
rect 16080 13144 16497 13172
rect 16080 13132 16086 13144
rect 16485 13141 16497 13144
rect 16531 13141 16543 13175
rect 16485 13135 16543 13141
rect 16758 13132 16764 13184
rect 16816 13172 16822 13184
rect 17494 13172 17500 13184
rect 16816 13144 17500 13172
rect 16816 13132 16822 13144
rect 17494 13132 17500 13144
rect 17552 13172 17558 13184
rect 17773 13175 17831 13181
rect 17773 13172 17785 13175
rect 17552 13144 17785 13172
rect 17552 13132 17558 13144
rect 17773 13141 17785 13144
rect 17819 13141 17831 13175
rect 17871 13172 17899 13212
rect 20530 13200 20536 13212
rect 20588 13200 20594 13252
rect 20708 13243 20766 13249
rect 20708 13209 20720 13243
rect 20754 13240 20766 13243
rect 21818 13240 21824 13252
rect 20754 13212 21824 13240
rect 20754 13209 20766 13212
rect 20708 13203 20766 13209
rect 21818 13200 21824 13212
rect 21876 13200 21882 13252
rect 21913 13243 21971 13249
rect 21913 13209 21925 13243
rect 21959 13209 21971 13243
rect 21913 13203 21971 13209
rect 25216 13243 25274 13249
rect 25216 13209 25228 13243
rect 25262 13240 25274 13243
rect 25498 13240 25504 13252
rect 25262 13212 25504 13240
rect 25262 13209 25274 13212
rect 25216 13203 25274 13209
rect 19613 13175 19671 13181
rect 19613 13172 19625 13175
rect 17871 13144 19625 13172
rect 17773 13135 17831 13141
rect 19613 13141 19625 13144
rect 19659 13141 19671 13175
rect 19613 13135 19671 13141
rect 19702 13132 19708 13184
rect 19760 13132 19766 13184
rect 21928 13172 21956 13203
rect 25498 13200 25504 13212
rect 25556 13200 25562 13252
rect 26528 13240 26556 13271
rect 27246 13268 27252 13280
rect 27304 13268 27310 13320
rect 27338 13268 27344 13320
rect 27396 13268 27402 13320
rect 27709 13311 27767 13317
rect 27709 13277 27721 13311
rect 27755 13308 27767 13311
rect 27890 13308 27896 13320
rect 27755 13280 27896 13308
rect 27755 13277 27767 13280
rect 27709 13271 27767 13277
rect 27890 13268 27896 13280
rect 27948 13268 27954 13320
rect 28810 13268 28816 13320
rect 28868 13268 28874 13320
rect 29012 13308 29040 13339
rect 28920 13280 29040 13308
rect 26344 13212 26556 13240
rect 26789 13243 26847 13249
rect 26344 13184 26372 13212
rect 26789 13209 26801 13243
rect 26835 13240 26847 13243
rect 27798 13240 27804 13252
rect 26835 13212 27804 13240
rect 26835 13209 26847 13212
rect 26789 13203 26847 13209
rect 27798 13200 27804 13212
rect 27856 13200 27862 13252
rect 28626 13200 28632 13252
rect 28684 13240 28690 13252
rect 28920 13240 28948 13280
rect 28684 13212 28948 13240
rect 28684 13200 28690 13212
rect 22830 13172 22836 13184
rect 21928 13144 22836 13172
rect 22830 13132 22836 13144
rect 22888 13172 22894 13184
rect 22925 13175 22983 13181
rect 22925 13172 22937 13175
rect 22888 13144 22937 13172
rect 22888 13132 22894 13144
rect 22925 13141 22937 13144
rect 22971 13141 22983 13175
rect 22925 13135 22983 13141
rect 23382 13132 23388 13184
rect 23440 13172 23446 13184
rect 23937 13175 23995 13181
rect 23937 13172 23949 13175
rect 23440 13144 23949 13172
rect 23440 13132 23446 13144
rect 23937 13141 23949 13144
rect 23983 13172 23995 13175
rect 24118 13172 24124 13184
rect 23983 13144 24124 13172
rect 23983 13141 23995 13144
rect 23937 13135 23995 13141
rect 24118 13132 24124 13144
rect 24176 13132 24182 13184
rect 26326 13132 26332 13184
rect 26384 13132 26390 13184
rect 26602 13132 26608 13184
rect 26660 13172 26666 13184
rect 27065 13175 27123 13181
rect 27065 13172 27077 13175
rect 26660 13144 27077 13172
rect 26660 13132 26666 13144
rect 27065 13141 27077 13144
rect 27111 13141 27123 13175
rect 27065 13135 27123 13141
rect 1104 13082 35328 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35328 13082
rect 1104 13008 35328 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 2866 12968 2872 12980
rect 1627 12940 2872 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 2866 12928 2872 12940
rect 2924 12928 2930 12980
rect 2958 12928 2964 12980
rect 3016 12928 3022 12980
rect 3973 12971 4031 12977
rect 3973 12937 3985 12971
rect 4019 12968 4031 12971
rect 4062 12968 4068 12980
rect 4019 12940 4068 12968
rect 4019 12937 4031 12940
rect 3973 12931 4031 12937
rect 4062 12928 4068 12940
rect 4120 12928 4126 12980
rect 4338 12928 4344 12980
rect 4396 12928 4402 12980
rect 6362 12928 6368 12980
rect 6420 12928 6426 12980
rect 6733 12971 6791 12977
rect 6733 12937 6745 12971
rect 6779 12968 6791 12971
rect 6914 12968 6920 12980
rect 6779 12940 6920 12968
rect 6779 12937 6791 12940
rect 6733 12931 6791 12937
rect 6914 12928 6920 12940
rect 6972 12928 6978 12980
rect 9217 12971 9275 12977
rect 9217 12937 9229 12971
rect 9263 12968 9275 12971
rect 12250 12968 12256 12980
rect 9263 12940 12256 12968
rect 9263 12937 9275 12940
rect 9217 12931 9275 12937
rect 12250 12928 12256 12940
rect 12308 12928 12314 12980
rect 14182 12928 14188 12980
rect 14240 12968 14246 12980
rect 15105 12971 15163 12977
rect 15105 12968 15117 12971
rect 14240 12940 15117 12968
rect 14240 12928 14246 12940
rect 15105 12937 15117 12940
rect 15151 12937 15163 12971
rect 15105 12931 15163 12937
rect 15654 12928 15660 12980
rect 15712 12928 15718 12980
rect 16022 12928 16028 12980
rect 16080 12928 16086 12980
rect 16117 12971 16175 12977
rect 16117 12937 16129 12971
rect 16163 12968 16175 12971
rect 16758 12968 16764 12980
rect 16163 12940 16764 12968
rect 16163 12937 16175 12940
rect 16117 12931 16175 12937
rect 16758 12928 16764 12940
rect 16816 12928 16822 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 17052 12940 17785 12968
rect 3421 12903 3479 12909
rect 3421 12869 3433 12903
rect 3467 12900 3479 12903
rect 4154 12900 4160 12912
rect 3467 12872 4160 12900
rect 3467 12869 3479 12872
rect 3421 12863 3479 12869
rect 4154 12860 4160 12872
rect 4212 12860 4218 12912
rect 6270 12860 6276 12912
rect 6328 12900 6334 12912
rect 9398 12900 9404 12912
rect 6328 12872 8800 12900
rect 6328 12860 6334 12872
rect 1302 12792 1308 12844
rect 1360 12832 1366 12844
rect 1397 12835 1455 12841
rect 1397 12832 1409 12835
rect 1360 12804 1409 12832
rect 1360 12792 1366 12804
rect 1397 12801 1409 12804
rect 1443 12832 1455 12835
rect 1673 12835 1731 12841
rect 1673 12832 1685 12835
rect 1443 12804 1685 12832
rect 1443 12801 1455 12804
rect 1397 12795 1455 12801
rect 1673 12801 1685 12804
rect 1719 12801 1731 12835
rect 1673 12795 1731 12801
rect 3329 12835 3387 12841
rect 3329 12801 3341 12835
rect 3375 12832 3387 12835
rect 3694 12832 3700 12844
rect 3375 12804 3700 12832
rect 3375 12801 3387 12804
rect 3329 12795 3387 12801
rect 3694 12792 3700 12804
rect 3752 12832 3758 12844
rect 4433 12835 4491 12841
rect 4433 12832 4445 12835
rect 3752 12804 4445 12832
rect 3752 12792 3758 12804
rect 4433 12801 4445 12804
rect 4479 12832 4491 12835
rect 6822 12832 6828 12844
rect 4479 12804 6828 12832
rect 4479 12801 4491 12804
rect 4433 12795 4491 12801
rect 6822 12792 6828 12804
rect 6880 12792 6886 12844
rect 8772 12841 8800 12872
rect 9048 12872 9404 12900
rect 8665 12835 8723 12841
rect 8665 12801 8677 12835
rect 8711 12801 8723 12835
rect 8665 12795 8723 12801
rect 8757 12835 8815 12841
rect 8757 12801 8769 12835
rect 8803 12801 8815 12835
rect 8757 12795 8815 12801
rect 3605 12767 3663 12773
rect 3605 12733 3617 12767
rect 3651 12764 3663 12767
rect 4617 12767 4675 12773
rect 3651 12736 3924 12764
rect 3651 12733 3663 12736
rect 3605 12727 3663 12733
rect 3896 12637 3924 12736
rect 4617 12733 4629 12767
rect 4663 12764 4675 12767
rect 4706 12764 4712 12776
rect 4663 12736 4712 12764
rect 4663 12733 4675 12736
rect 4617 12727 4675 12733
rect 4706 12724 4712 12736
rect 4764 12764 4770 12776
rect 5258 12764 5264 12776
rect 4764 12736 5264 12764
rect 4764 12724 4770 12736
rect 5258 12724 5264 12736
rect 5316 12724 5322 12776
rect 7009 12767 7067 12773
rect 7009 12733 7021 12767
rect 7055 12764 7067 12767
rect 7190 12764 7196 12776
rect 7055 12736 7196 12764
rect 7055 12733 7067 12736
rect 7009 12727 7067 12733
rect 7190 12724 7196 12736
rect 7248 12764 7254 12776
rect 8202 12764 8208 12776
rect 7248 12736 8208 12764
rect 7248 12724 7254 12736
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 8680 12764 8708 12795
rect 8846 12792 8852 12844
rect 8904 12832 8910 12844
rect 9048 12841 9076 12872
rect 9398 12860 9404 12872
rect 9456 12860 9462 12912
rect 9585 12903 9643 12909
rect 9585 12869 9597 12903
rect 9631 12900 9643 12903
rect 11146 12900 11152 12912
rect 9631 12872 11152 12900
rect 9631 12869 9643 12872
rect 9585 12863 9643 12869
rect 8941 12835 8999 12841
rect 8941 12832 8953 12835
rect 8904 12804 8953 12832
rect 8904 12792 8910 12804
rect 8941 12801 8953 12804
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12801 9091 12835
rect 9033 12795 9091 12801
rect 9600 12764 9628 12863
rect 11146 12860 11152 12872
rect 11204 12860 11210 12912
rect 13992 12903 14050 12909
rect 13992 12869 14004 12903
rect 14038 12900 14050 12903
rect 14090 12900 14096 12912
rect 14038 12872 14096 12900
rect 14038 12869 14050 12872
rect 13992 12863 14050 12869
rect 14090 12860 14096 12872
rect 14148 12860 14154 12912
rect 9674 12792 9680 12844
rect 9732 12832 9738 12844
rect 10042 12832 10048 12844
rect 9732 12804 10048 12832
rect 9732 12792 9738 12804
rect 10042 12792 10048 12804
rect 10100 12832 10106 12844
rect 16040 12832 16068 12928
rect 16942 12860 16948 12912
rect 17000 12900 17006 12912
rect 17052 12909 17080 12940
rect 17773 12937 17785 12940
rect 17819 12968 17831 12971
rect 24762 12968 24768 12980
rect 17819 12940 24768 12968
rect 17819 12937 17831 12940
rect 17773 12931 17831 12937
rect 24762 12928 24768 12940
rect 24820 12928 24826 12980
rect 25498 12928 25504 12980
rect 25556 12928 25562 12980
rect 25869 12971 25927 12977
rect 25869 12937 25881 12971
rect 25915 12968 25927 12971
rect 26326 12968 26332 12980
rect 25915 12940 26332 12968
rect 25915 12937 25927 12940
rect 25869 12931 25927 12937
rect 26326 12928 26332 12940
rect 26384 12928 26390 12980
rect 26605 12971 26663 12977
rect 26605 12937 26617 12971
rect 26651 12968 26663 12971
rect 26878 12968 26884 12980
rect 26651 12940 26884 12968
rect 26651 12937 26663 12940
rect 26605 12931 26663 12937
rect 26878 12928 26884 12940
rect 26936 12928 26942 12980
rect 27798 12928 27804 12980
rect 27856 12968 27862 12980
rect 28353 12971 28411 12977
rect 28353 12968 28365 12971
rect 27856 12940 28365 12968
rect 27856 12928 27862 12940
rect 28353 12937 28365 12940
rect 28399 12937 28411 12971
rect 28353 12931 28411 12937
rect 17037 12903 17095 12909
rect 17037 12900 17049 12903
rect 17000 12872 17049 12900
rect 17000 12860 17006 12872
rect 17037 12869 17049 12872
rect 17083 12869 17095 12903
rect 17037 12863 17095 12869
rect 17954 12860 17960 12912
rect 18012 12900 18018 12912
rect 20990 12900 20996 12912
rect 18012 12872 18184 12900
rect 18012 12860 18018 12872
rect 16853 12835 16911 12841
rect 16853 12832 16865 12835
rect 10100 12804 15976 12832
rect 16040 12804 16865 12832
rect 10100 12792 10106 12804
rect 8680 12736 9628 12764
rect 12526 12724 12532 12776
rect 12584 12764 12590 12776
rect 13725 12767 13783 12773
rect 13725 12764 13737 12767
rect 12584 12736 13737 12764
rect 12584 12724 12590 12736
rect 13725 12733 13737 12736
rect 13771 12733 13783 12767
rect 15948 12764 15976 12804
rect 16853 12801 16865 12804
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 17126 12792 17132 12844
rect 17184 12792 17190 12844
rect 17221 12835 17279 12841
rect 17221 12801 17233 12835
rect 17267 12832 17279 12835
rect 17497 12835 17555 12841
rect 17497 12832 17509 12835
rect 17267 12804 17509 12832
rect 17267 12801 17279 12804
rect 17221 12795 17279 12801
rect 17497 12801 17509 12804
rect 17543 12832 17555 12835
rect 17586 12832 17592 12844
rect 17543 12804 17592 12832
rect 17543 12801 17555 12804
rect 17497 12795 17555 12801
rect 16301 12767 16359 12773
rect 16301 12764 16313 12767
rect 15948 12736 16313 12764
rect 13725 12727 13783 12733
rect 16301 12733 16313 12736
rect 16347 12733 16359 12767
rect 16301 12727 16359 12733
rect 6454 12656 6460 12708
rect 6512 12696 6518 12708
rect 7377 12699 7435 12705
rect 7377 12696 7389 12699
rect 6512 12668 7389 12696
rect 6512 12656 6518 12668
rect 7377 12665 7389 12668
rect 7423 12665 7435 12699
rect 16316 12696 16344 12727
rect 16574 12724 16580 12776
rect 16632 12764 16638 12776
rect 17236 12764 17264 12795
rect 17586 12792 17592 12804
rect 17644 12792 17650 12844
rect 18156 12841 18184 12872
rect 18248 12872 20996 12900
rect 18049 12835 18107 12841
rect 18049 12801 18061 12835
rect 18095 12801 18107 12835
rect 18049 12795 18107 12801
rect 18142 12835 18200 12841
rect 18142 12801 18154 12835
rect 18188 12801 18200 12835
rect 18142 12795 18200 12801
rect 16632 12736 17264 12764
rect 16632 12724 16638 12736
rect 16761 12699 16819 12705
rect 16761 12696 16773 12699
rect 16316 12668 16773 12696
rect 7377 12659 7435 12665
rect 16761 12665 16773 12668
rect 16807 12696 16819 12699
rect 17405 12699 17463 12705
rect 16807 12668 16988 12696
rect 16807 12665 16819 12668
rect 16761 12659 16819 12665
rect 3881 12631 3939 12637
rect 3881 12597 3893 12631
rect 3927 12628 3939 12631
rect 5350 12628 5356 12640
rect 3927 12600 5356 12628
rect 3927 12597 3939 12600
rect 3881 12591 3939 12597
rect 5350 12588 5356 12600
rect 5408 12588 5414 12640
rect 12710 12588 12716 12640
rect 12768 12628 12774 12640
rect 15930 12628 15936 12640
rect 12768 12600 15936 12628
rect 12768 12588 12774 12600
rect 15930 12588 15936 12600
rect 15988 12628 15994 12640
rect 16850 12628 16856 12640
rect 15988 12600 16856 12628
rect 15988 12588 15994 12600
rect 16850 12588 16856 12600
rect 16908 12588 16914 12640
rect 16960 12628 16988 12668
rect 17405 12665 17417 12699
rect 17451 12696 17463 12699
rect 18064 12696 18092 12795
rect 17451 12668 18092 12696
rect 17451 12665 17463 12668
rect 17405 12659 17463 12665
rect 18248 12628 18276 12872
rect 20990 12860 20996 12872
rect 21048 12860 21054 12912
rect 21269 12903 21327 12909
rect 21269 12900 21281 12903
rect 21192 12872 21281 12900
rect 18325 12835 18383 12841
rect 18325 12801 18337 12835
rect 18371 12801 18383 12835
rect 18325 12795 18383 12801
rect 16960 12600 18276 12628
rect 18340 12628 18368 12795
rect 18414 12792 18420 12844
rect 18472 12792 18478 12844
rect 18506 12792 18512 12844
rect 18564 12841 18570 12844
rect 18564 12832 18572 12841
rect 18564 12804 18609 12832
rect 18564 12795 18572 12804
rect 18564 12792 18570 12795
rect 18782 12792 18788 12844
rect 18840 12792 18846 12844
rect 18969 12835 19027 12841
rect 18969 12801 18981 12835
rect 19015 12801 19027 12835
rect 18969 12795 19027 12801
rect 18984 12764 19012 12795
rect 19058 12792 19064 12844
rect 19116 12792 19122 12844
rect 19150 12792 19156 12844
rect 19208 12792 19214 12844
rect 19337 12835 19395 12841
rect 19337 12801 19349 12835
rect 19383 12832 19395 12835
rect 19702 12832 19708 12844
rect 19383 12804 19708 12832
rect 19383 12801 19395 12804
rect 19337 12795 19395 12801
rect 19702 12792 19708 12804
rect 19760 12792 19766 12844
rect 20898 12792 20904 12844
rect 20956 12792 20962 12844
rect 21082 12792 21088 12844
rect 21140 12792 21146 12844
rect 18708 12736 19012 12764
rect 18708 12705 18736 12736
rect 19242 12724 19248 12776
rect 19300 12764 19306 12776
rect 19613 12767 19671 12773
rect 19613 12764 19625 12767
rect 19300 12736 19625 12764
rect 19300 12724 19306 12736
rect 19613 12733 19625 12736
rect 19659 12733 19671 12767
rect 20916 12764 20944 12792
rect 21192 12764 21220 12872
rect 21269 12869 21281 12872
rect 21315 12869 21327 12903
rect 21269 12863 21327 12869
rect 21361 12903 21419 12909
rect 21361 12869 21373 12903
rect 21407 12900 21419 12903
rect 22186 12900 22192 12912
rect 21407 12872 22192 12900
rect 21407 12869 21419 12872
rect 21361 12863 21419 12869
rect 22186 12860 22192 12872
rect 22244 12860 22250 12912
rect 24670 12900 24676 12912
rect 24504 12872 24676 12900
rect 21453 12835 21511 12841
rect 21453 12801 21465 12835
rect 21499 12832 21511 12835
rect 21499 12804 21588 12832
rect 21499 12801 21511 12804
rect 21453 12795 21511 12801
rect 20916 12736 21220 12764
rect 19613 12727 19671 12733
rect 18693 12699 18751 12705
rect 18693 12665 18705 12699
rect 18739 12665 18751 12699
rect 18693 12659 18751 12665
rect 18782 12656 18788 12708
rect 18840 12696 18846 12708
rect 19260 12696 19288 12724
rect 19797 12699 19855 12705
rect 19797 12696 19809 12699
rect 18840 12668 19288 12696
rect 19444 12668 19809 12696
rect 18840 12656 18846 12668
rect 19444 12628 19472 12668
rect 19797 12665 19809 12668
rect 19843 12696 19855 12699
rect 20622 12696 20628 12708
rect 19843 12668 20628 12696
rect 19843 12665 19855 12668
rect 19797 12659 19855 12665
rect 20622 12656 20628 12668
rect 20680 12656 20686 12708
rect 20806 12656 20812 12708
rect 20864 12696 20870 12708
rect 21560 12696 21588 12804
rect 21726 12792 21732 12844
rect 21784 12832 21790 12844
rect 21913 12835 21971 12841
rect 21913 12832 21925 12835
rect 21784 12804 21925 12832
rect 21784 12792 21790 12804
rect 21913 12801 21925 12804
rect 21959 12801 21971 12835
rect 23201 12835 23259 12841
rect 23201 12832 23213 12835
rect 21913 12795 21971 12801
rect 22066 12804 23213 12832
rect 20864 12668 21588 12696
rect 20864 12656 20870 12668
rect 18340 12600 19472 12628
rect 19518 12588 19524 12640
rect 19576 12588 19582 12640
rect 19702 12588 19708 12640
rect 19760 12628 19766 12640
rect 19981 12631 20039 12637
rect 19981 12628 19993 12631
rect 19760 12600 19993 12628
rect 19760 12588 19766 12600
rect 19981 12597 19993 12600
rect 20027 12597 20039 12631
rect 21560 12628 21588 12668
rect 21637 12699 21695 12705
rect 21637 12665 21649 12699
rect 21683 12696 21695 12699
rect 22066 12696 22094 12804
rect 23201 12801 23213 12804
rect 23247 12801 23259 12835
rect 23201 12795 23259 12801
rect 23290 12792 23296 12844
rect 23348 12792 23354 12844
rect 23382 12792 23388 12844
rect 23440 12832 23446 12844
rect 23477 12835 23535 12841
rect 23477 12832 23489 12835
rect 23440 12804 23489 12832
rect 23440 12792 23446 12804
rect 23477 12801 23489 12804
rect 23523 12801 23535 12835
rect 23477 12795 23535 12801
rect 23566 12792 23572 12844
rect 23624 12792 23630 12844
rect 23658 12792 23664 12844
rect 23716 12841 23722 12844
rect 24504 12841 24532 12872
rect 24670 12860 24676 12872
rect 24728 12900 24734 12912
rect 25133 12903 25191 12909
rect 25133 12900 25145 12903
rect 24728 12872 25145 12900
rect 24728 12860 24734 12872
rect 25133 12869 25145 12872
rect 25179 12900 25191 12903
rect 26694 12900 26700 12912
rect 25179 12872 26700 12900
rect 25179 12869 25191 12872
rect 25133 12863 25191 12869
rect 26694 12860 26700 12872
rect 26752 12860 26758 12912
rect 27338 12860 27344 12912
rect 27396 12900 27402 12912
rect 28445 12903 28503 12909
rect 28445 12900 28457 12903
rect 27396 12872 28457 12900
rect 27396 12860 27402 12872
rect 28445 12869 28457 12872
rect 28491 12900 28503 12903
rect 28813 12903 28871 12909
rect 28813 12900 28825 12903
rect 28491 12872 28825 12900
rect 28491 12869 28503 12872
rect 28445 12863 28503 12869
rect 28813 12869 28825 12872
rect 28859 12869 28871 12903
rect 28813 12863 28871 12869
rect 33134 12860 33140 12912
rect 33192 12860 33198 12912
rect 23716 12832 23724 12841
rect 24489 12835 24547 12841
rect 23716 12804 23761 12832
rect 23716 12795 23724 12804
rect 24489 12801 24501 12835
rect 24535 12801 24547 12835
rect 24489 12795 24547 12801
rect 23716 12792 23722 12795
rect 26510 12792 26516 12844
rect 26568 12792 26574 12844
rect 26970 12792 26976 12844
rect 27028 12792 27034 12844
rect 27246 12841 27252 12844
rect 27240 12795 27252 12841
rect 27246 12792 27252 12795
rect 27304 12792 27310 12844
rect 32122 12792 32128 12844
rect 32180 12792 32186 12844
rect 33870 12792 33876 12844
rect 33928 12832 33934 12844
rect 34517 12835 34575 12841
rect 34517 12832 34529 12835
rect 33928 12804 34529 12832
rect 33928 12792 33934 12804
rect 34517 12801 34529 12804
rect 34563 12801 34575 12835
rect 34517 12795 34575 12801
rect 22189 12767 22247 12773
rect 22189 12733 22201 12767
rect 22235 12764 22247 12767
rect 22554 12764 22560 12776
rect 22235 12736 22560 12764
rect 22235 12733 22247 12736
rect 22189 12727 22247 12733
rect 22554 12724 22560 12736
rect 22612 12724 22618 12776
rect 24765 12767 24823 12773
rect 24765 12733 24777 12767
rect 24811 12764 24823 12767
rect 25222 12764 25228 12776
rect 24811 12736 25228 12764
rect 24811 12733 24823 12736
rect 24765 12727 24823 12733
rect 25222 12724 25228 12736
rect 25280 12724 25286 12776
rect 25961 12767 26019 12773
rect 25961 12733 25973 12767
rect 26007 12733 26019 12767
rect 25961 12727 26019 12733
rect 21683 12668 22094 12696
rect 21683 12665 21695 12668
rect 21637 12659 21695 12665
rect 22738 12656 22744 12708
rect 22796 12696 22802 12708
rect 23017 12699 23075 12705
rect 23017 12696 23029 12699
rect 22796 12668 23029 12696
rect 22796 12656 22802 12668
rect 23017 12665 23029 12668
rect 23063 12665 23075 12699
rect 23017 12659 23075 12665
rect 23845 12699 23903 12705
rect 23845 12665 23857 12699
rect 23891 12696 23903 12699
rect 24946 12696 24952 12708
rect 23891 12668 24952 12696
rect 23891 12665 23903 12668
rect 23845 12659 23903 12665
rect 24946 12656 24952 12668
rect 25004 12656 25010 12708
rect 25976 12696 26004 12727
rect 26142 12724 26148 12776
rect 26200 12724 26206 12776
rect 32398 12724 32404 12776
rect 32456 12724 32462 12776
rect 34793 12767 34851 12773
rect 34793 12733 34805 12767
rect 34839 12764 34851 12767
rect 35342 12764 35348 12776
rect 34839 12736 35348 12764
rect 34839 12733 34851 12736
rect 34793 12727 34851 12733
rect 35342 12724 35348 12736
rect 35400 12724 35406 12776
rect 26329 12699 26387 12705
rect 26329 12696 26341 12699
rect 25976 12668 26341 12696
rect 26329 12665 26341 12668
rect 26375 12696 26387 12699
rect 26418 12696 26424 12708
rect 26375 12668 26424 12696
rect 26375 12665 26387 12668
rect 26329 12659 26387 12665
rect 26418 12656 26424 12668
rect 26476 12656 26482 12708
rect 22833 12631 22891 12637
rect 22833 12628 22845 12631
rect 21560 12600 22845 12628
rect 19981 12591 20039 12597
rect 22833 12597 22845 12600
rect 22879 12597 22891 12631
rect 22833 12591 22891 12597
rect 24854 12588 24860 12640
rect 24912 12588 24918 12640
rect 25590 12588 25596 12640
rect 25648 12628 25654 12640
rect 28626 12628 28632 12640
rect 25648 12600 28632 12628
rect 25648 12588 25654 12600
rect 28626 12588 28632 12600
rect 28684 12588 28690 12640
rect 33870 12588 33876 12640
rect 33928 12588 33934 12640
rect 1104 12538 35328 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 35328 12538
rect 1104 12464 35328 12486
rect 12986 12384 12992 12436
rect 13044 12384 13050 12436
rect 13357 12427 13415 12433
rect 13357 12393 13369 12427
rect 13403 12424 13415 12427
rect 13906 12424 13912 12436
rect 13403 12396 13912 12424
rect 13403 12393 13415 12396
rect 13357 12387 13415 12393
rect 13906 12384 13912 12396
rect 13964 12384 13970 12436
rect 16298 12384 16304 12436
rect 16356 12424 16362 12436
rect 20990 12424 20996 12436
rect 16356 12396 20996 12424
rect 16356 12384 16362 12396
rect 20990 12384 20996 12396
rect 21048 12384 21054 12436
rect 21082 12384 21088 12436
rect 21140 12424 21146 12436
rect 21177 12427 21235 12433
rect 21177 12424 21189 12427
rect 21140 12396 21189 12424
rect 21140 12384 21146 12396
rect 21177 12393 21189 12396
rect 21223 12393 21235 12427
rect 21177 12387 21235 12393
rect 21818 12384 21824 12436
rect 21876 12384 21882 12436
rect 22094 12384 22100 12436
rect 22152 12424 22158 12436
rect 22738 12424 22744 12436
rect 22152 12396 22744 12424
rect 22152 12384 22158 12396
rect 22738 12384 22744 12396
rect 22796 12384 22802 12436
rect 23566 12384 23572 12436
rect 23624 12424 23630 12436
rect 24213 12427 24271 12433
rect 24213 12424 24225 12427
rect 23624 12396 24225 12424
rect 23624 12384 23630 12396
rect 23860 12368 23888 12396
rect 24213 12393 24225 12396
rect 24259 12393 24271 12427
rect 25133 12427 25191 12433
rect 25133 12424 25145 12427
rect 24213 12387 24271 12393
rect 24504 12396 25145 12424
rect 24504 12368 24532 12396
rect 25133 12393 25145 12396
rect 25179 12393 25191 12427
rect 25133 12387 25191 12393
rect 25774 12384 25780 12436
rect 25832 12384 25838 12436
rect 26602 12384 26608 12436
rect 26660 12384 26666 12436
rect 26789 12427 26847 12433
rect 26789 12393 26801 12427
rect 26835 12424 26847 12427
rect 27062 12424 27068 12436
rect 26835 12396 27068 12424
rect 26835 12393 26847 12396
rect 26789 12387 26847 12393
rect 27062 12384 27068 12396
rect 27120 12384 27126 12436
rect 27246 12384 27252 12436
rect 27304 12384 27310 12436
rect 29454 12384 29460 12436
rect 29512 12424 29518 12436
rect 29822 12424 29828 12436
rect 29512 12396 29828 12424
rect 29512 12384 29518 12396
rect 29822 12384 29828 12396
rect 29880 12424 29886 12436
rect 32217 12427 32275 12433
rect 29880 12396 31754 12424
rect 29880 12384 29886 12396
rect 8478 12316 8484 12368
rect 8536 12356 8542 12368
rect 10134 12356 10140 12368
rect 8536 12328 10140 12356
rect 8536 12316 8542 12328
rect 10134 12316 10140 12328
rect 10192 12316 10198 12368
rect 10318 12316 10324 12368
rect 10376 12356 10382 12368
rect 18693 12359 18751 12365
rect 18693 12356 18705 12359
rect 10376 12328 18705 12356
rect 10376 12316 10382 12328
rect 18693 12325 18705 12328
rect 18739 12356 18751 12359
rect 19521 12359 19579 12365
rect 19521 12356 19533 12359
rect 18739 12328 19533 12356
rect 18739 12325 18751 12328
rect 18693 12319 18751 12325
rect 19521 12325 19533 12328
rect 19567 12356 19579 12359
rect 19610 12356 19616 12368
rect 19567 12328 19616 12356
rect 19567 12325 19579 12328
rect 19521 12319 19579 12325
rect 19610 12316 19616 12328
rect 19668 12316 19674 12368
rect 20898 12316 20904 12368
rect 20956 12356 20962 12368
rect 21266 12356 21272 12368
rect 20956 12328 21272 12356
rect 20956 12316 20962 12328
rect 21266 12316 21272 12328
rect 21324 12356 21330 12368
rect 21453 12359 21511 12365
rect 21453 12356 21465 12359
rect 21324 12328 21465 12356
rect 21324 12316 21330 12328
rect 21453 12325 21465 12328
rect 21499 12356 21511 12359
rect 22649 12359 22707 12365
rect 22649 12356 22661 12359
rect 21499 12328 22661 12356
rect 21499 12325 21511 12328
rect 21453 12319 21511 12325
rect 22649 12325 22661 12328
rect 22695 12325 22707 12359
rect 22649 12319 22707 12325
rect 23842 12316 23848 12368
rect 23900 12316 23906 12368
rect 24118 12316 24124 12368
rect 24176 12356 24182 12368
rect 24486 12356 24492 12368
rect 24176 12328 24492 12356
rect 24176 12316 24182 12328
rect 24486 12316 24492 12328
rect 24544 12316 24550 12368
rect 26234 12316 26240 12368
rect 26292 12356 26298 12368
rect 26881 12359 26939 12365
rect 26881 12356 26893 12359
rect 26292 12328 26893 12356
rect 26292 12316 26298 12328
rect 26881 12325 26893 12328
rect 26927 12325 26939 12359
rect 29638 12356 29644 12368
rect 26881 12319 26939 12325
rect 26988 12328 29644 12356
rect 7653 12291 7711 12297
rect 7653 12257 7665 12291
rect 7699 12288 7711 12291
rect 7926 12288 7932 12300
rect 7699 12260 7932 12288
rect 7699 12257 7711 12260
rect 7653 12251 7711 12257
rect 7926 12248 7932 12260
rect 7984 12248 7990 12300
rect 8665 12291 8723 12297
rect 8665 12288 8677 12291
rect 8220 12260 8677 12288
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 8021 12223 8079 12229
rect 8021 12220 8033 12223
rect 5592 12192 6776 12220
rect 5592 12180 5598 12192
rect 6748 12164 6776 12192
rect 7392 12192 8033 12220
rect 5994 12112 6000 12164
rect 6052 12152 6058 12164
rect 6454 12152 6460 12164
rect 6052 12124 6460 12152
rect 6052 12112 6058 12124
rect 6454 12112 6460 12124
rect 6512 12112 6518 12164
rect 6730 12112 6736 12164
rect 6788 12112 6794 12164
rect 7392 12096 7420 12192
rect 8021 12189 8033 12192
rect 8067 12189 8079 12223
rect 8021 12183 8079 12189
rect 8110 12180 8116 12232
rect 8168 12220 8174 12232
rect 8220 12229 8248 12260
rect 8665 12257 8677 12260
rect 8711 12257 8723 12291
rect 13170 12288 13176 12300
rect 8665 12251 8723 12257
rect 12636 12260 13176 12288
rect 8205 12223 8263 12229
rect 8205 12220 8217 12223
rect 8168 12192 8217 12220
rect 8168 12180 8174 12192
rect 8205 12189 8217 12192
rect 8251 12189 8263 12223
rect 8205 12183 8263 12189
rect 8389 12223 8447 12229
rect 8389 12189 8401 12223
rect 8435 12220 8447 12223
rect 8754 12220 8760 12232
rect 8435 12192 8760 12220
rect 8435 12189 8447 12192
rect 8389 12183 8447 12189
rect 8754 12180 8760 12192
rect 8812 12220 8818 12232
rect 8941 12223 8999 12229
rect 8941 12220 8953 12223
rect 8812 12192 8953 12220
rect 8812 12180 8818 12192
rect 8941 12189 8953 12192
rect 8987 12189 8999 12223
rect 8941 12183 8999 12189
rect 11330 12180 11336 12232
rect 11388 12220 11394 12232
rect 12636 12229 12664 12260
rect 13170 12248 13176 12260
rect 13228 12288 13234 12300
rect 13722 12288 13728 12300
rect 13228 12260 13728 12288
rect 13228 12248 13234 12260
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 18598 12248 18604 12300
rect 18656 12288 18662 12300
rect 19334 12288 19340 12300
rect 18656 12260 19340 12288
rect 18656 12248 18662 12260
rect 12437 12223 12495 12229
rect 12437 12220 12449 12223
rect 11388 12192 12449 12220
rect 11388 12180 11394 12192
rect 12437 12189 12449 12192
rect 12483 12189 12495 12223
rect 12437 12183 12495 12189
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12189 12679 12223
rect 12621 12183 12679 12189
rect 12805 12223 12863 12229
rect 12805 12189 12817 12223
rect 12851 12220 12863 12223
rect 13998 12220 14004 12232
rect 12851 12192 14004 12220
rect 12851 12189 12863 12192
rect 12805 12183 12863 12189
rect 13998 12180 14004 12192
rect 14056 12180 14062 12232
rect 14274 12180 14280 12232
rect 14332 12220 14338 12232
rect 14826 12220 14832 12232
rect 14332 12192 14832 12220
rect 14332 12180 14338 12192
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 17034 12180 17040 12232
rect 17092 12220 17098 12232
rect 17678 12220 17684 12232
rect 17092 12192 17684 12220
rect 17092 12180 17098 12192
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 18892 12229 18920 12260
rect 19334 12248 19340 12260
rect 19392 12248 19398 12300
rect 19426 12248 19432 12300
rect 19484 12288 19490 12300
rect 19797 12291 19855 12297
rect 19797 12288 19809 12291
rect 19484 12260 19809 12288
rect 19484 12248 19490 12260
rect 19797 12257 19809 12260
rect 19843 12257 19855 12291
rect 19797 12251 19855 12257
rect 20806 12248 20812 12300
rect 20864 12288 20870 12300
rect 22094 12288 22100 12300
rect 20864 12260 22100 12288
rect 20864 12248 20870 12260
rect 22094 12248 22100 12260
rect 22152 12288 22158 12300
rect 22373 12291 22431 12297
rect 22373 12288 22385 12291
rect 22152 12260 22385 12288
rect 22152 12248 22158 12260
rect 22373 12257 22385 12260
rect 22419 12257 22431 12291
rect 22373 12251 22431 12257
rect 24946 12248 24952 12300
rect 25004 12288 25010 12300
rect 26513 12291 26571 12297
rect 26513 12288 26525 12291
rect 25004 12260 26525 12288
rect 25004 12248 25010 12260
rect 26513 12257 26525 12260
rect 26559 12257 26571 12291
rect 26513 12251 26571 12257
rect 18877 12223 18935 12229
rect 18877 12189 18889 12223
rect 18923 12189 18935 12223
rect 21637 12223 21695 12229
rect 18877 12183 18935 12189
rect 18984 12192 21588 12220
rect 8297 12155 8355 12161
rect 8297 12121 8309 12155
rect 8343 12152 8355 12155
rect 8343 12124 8432 12152
rect 8343 12121 8355 12124
rect 8297 12115 8355 12121
rect 8404 12096 8432 12124
rect 9398 12112 9404 12164
rect 9456 12152 9462 12164
rect 12713 12155 12771 12161
rect 9456 12124 12434 12152
rect 9456 12112 9462 12124
rect 7006 12044 7012 12096
rect 7064 12044 7070 12096
rect 7374 12044 7380 12096
rect 7432 12044 7438 12096
rect 7466 12044 7472 12096
rect 7524 12044 7530 12096
rect 7926 12044 7932 12096
rect 7984 12044 7990 12096
rect 8386 12044 8392 12096
rect 8444 12044 8450 12096
rect 8573 12087 8631 12093
rect 8573 12053 8585 12087
rect 8619 12084 8631 12087
rect 10686 12084 10692 12096
rect 8619 12056 10692 12084
rect 8619 12053 8631 12056
rect 8573 12047 8631 12053
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 12406 12084 12434 12124
rect 12713 12121 12725 12155
rect 12759 12152 12771 12155
rect 13170 12152 13176 12164
rect 12759 12124 13176 12152
rect 12759 12121 12771 12124
rect 12713 12115 12771 12121
rect 13170 12112 13176 12124
rect 13228 12112 13234 12164
rect 16574 12152 16580 12164
rect 13280 12124 16580 12152
rect 13280 12084 13308 12124
rect 16574 12112 16580 12124
rect 16632 12152 16638 12164
rect 17310 12152 17316 12164
rect 16632 12124 17316 12152
rect 16632 12112 16638 12124
rect 17310 12112 17316 12124
rect 17368 12152 17374 12164
rect 18984 12152 19012 12192
rect 17368 12124 19012 12152
rect 20064 12155 20122 12161
rect 17368 12112 17374 12124
rect 20064 12121 20076 12155
rect 20110 12152 20122 12155
rect 20346 12152 20352 12164
rect 20110 12124 20352 12152
rect 20110 12121 20122 12124
rect 20064 12115 20122 12121
rect 20346 12112 20352 12124
rect 20404 12112 20410 12164
rect 21560 12152 21588 12192
rect 21637 12189 21649 12223
rect 21683 12220 21695 12223
rect 22002 12220 22008 12232
rect 21683 12192 22008 12220
rect 21683 12189 21695 12192
rect 21637 12183 21695 12189
rect 22002 12180 22008 12192
rect 22060 12180 22066 12232
rect 22186 12180 22192 12232
rect 22244 12180 22250 12232
rect 22462 12180 22468 12232
rect 22520 12220 22526 12232
rect 22833 12223 22891 12229
rect 22833 12220 22845 12223
rect 22520 12192 22845 12220
rect 22520 12180 22526 12192
rect 22833 12189 22845 12192
rect 22879 12220 22891 12223
rect 22922 12220 22928 12232
rect 22879 12192 22928 12220
rect 22879 12189 22891 12192
rect 22833 12183 22891 12189
rect 22922 12180 22928 12192
rect 22980 12180 22986 12232
rect 23658 12220 23664 12232
rect 23032 12192 23664 12220
rect 23032 12152 23060 12192
rect 23658 12180 23664 12192
rect 23716 12180 23722 12232
rect 24673 12223 24731 12229
rect 24673 12189 24685 12223
rect 24719 12189 24731 12223
rect 24673 12183 24731 12189
rect 25041 12223 25099 12229
rect 25041 12189 25053 12223
rect 25087 12220 25099 12223
rect 25774 12220 25780 12232
rect 25087 12192 25780 12220
rect 25087 12189 25099 12192
rect 25041 12183 25099 12189
rect 21560 12124 23060 12152
rect 23100 12155 23158 12161
rect 23100 12121 23112 12155
rect 23146 12152 23158 12155
rect 23474 12152 23480 12164
rect 23146 12124 23480 12152
rect 23146 12121 23158 12124
rect 23100 12115 23158 12121
rect 23474 12112 23480 12124
rect 23532 12112 23538 12164
rect 12406 12056 13308 12084
rect 19610 12044 19616 12096
rect 19668 12084 19674 12096
rect 20162 12084 20168 12096
rect 19668 12056 20168 12084
rect 19668 12044 19674 12056
rect 20162 12044 20168 12056
rect 20220 12044 20226 12096
rect 22281 12087 22339 12093
rect 22281 12053 22293 12087
rect 22327 12084 22339 12087
rect 22646 12084 22652 12096
rect 22327 12056 22652 12084
rect 22327 12053 22339 12056
rect 22281 12047 22339 12053
rect 22646 12044 22652 12056
rect 22704 12044 22710 12096
rect 23676 12084 23704 12180
rect 24688 12152 24716 12183
rect 25774 12180 25780 12192
rect 25832 12180 25838 12232
rect 26326 12180 26332 12232
rect 26384 12220 26390 12232
rect 26421 12223 26479 12229
rect 26421 12220 26433 12223
rect 26384 12192 26433 12220
rect 26384 12180 26390 12192
rect 26421 12189 26433 12192
rect 26467 12189 26479 12223
rect 26421 12183 26479 12189
rect 25409 12155 25467 12161
rect 25409 12152 25421 12155
rect 24688 12124 25421 12152
rect 25409 12121 25421 12124
rect 25455 12152 25467 12155
rect 26988 12152 27016 12328
rect 29638 12316 29644 12328
rect 29696 12316 29702 12368
rect 31726 12356 31754 12396
rect 32217 12393 32229 12427
rect 32263 12424 32275 12427
rect 32398 12424 32404 12436
rect 32263 12396 32404 12424
rect 32263 12393 32275 12396
rect 32217 12387 32275 12393
rect 32398 12384 32404 12396
rect 32456 12384 32462 12436
rect 33134 12384 33140 12436
rect 33192 12424 33198 12436
rect 33229 12427 33287 12433
rect 33229 12424 33241 12427
rect 33192 12396 33241 12424
rect 33192 12384 33198 12396
rect 33229 12393 33241 12396
rect 33275 12393 33287 12427
rect 33229 12387 33287 12393
rect 32858 12356 32864 12368
rect 31726 12328 32864 12356
rect 32858 12316 32864 12328
rect 32916 12316 32922 12368
rect 27522 12248 27528 12300
rect 27580 12288 27586 12300
rect 27801 12291 27859 12297
rect 27801 12288 27813 12291
rect 27580 12260 27813 12288
rect 27580 12248 27586 12260
rect 27801 12257 27813 12260
rect 27847 12288 27859 12291
rect 28077 12291 28135 12297
rect 28077 12288 28089 12291
rect 27847 12260 28089 12288
rect 27847 12257 27859 12260
rect 27801 12251 27859 12257
rect 28077 12257 28089 12260
rect 28123 12257 28135 12291
rect 28077 12251 28135 12257
rect 29730 12248 29736 12300
rect 29788 12288 29794 12300
rect 29825 12291 29883 12297
rect 29825 12288 29837 12291
rect 29788 12260 29837 12288
rect 29788 12248 29794 12260
rect 29825 12257 29837 12260
rect 29871 12257 29883 12291
rect 33870 12288 33876 12300
rect 29825 12251 29883 12257
rect 31956 12260 33876 12288
rect 27617 12223 27675 12229
rect 27617 12189 27629 12223
rect 27663 12220 27675 12223
rect 27890 12220 27896 12232
rect 27663 12192 27896 12220
rect 27663 12189 27675 12192
rect 27617 12183 27675 12189
rect 27890 12180 27896 12192
rect 27948 12180 27954 12232
rect 30024 12192 30236 12220
rect 25455 12124 27016 12152
rect 25455 12121 25467 12124
rect 25409 12115 25467 12121
rect 27062 12112 27068 12164
rect 27120 12152 27126 12164
rect 30024 12152 30052 12192
rect 30098 12161 30104 12164
rect 27120 12124 30052 12152
rect 27120 12112 27126 12124
rect 30092 12115 30104 12161
rect 30098 12112 30104 12115
rect 30156 12112 30162 12164
rect 30208 12152 30236 12192
rect 31386 12180 31392 12232
rect 31444 12220 31450 12232
rect 31956 12229 31984 12260
rect 33870 12248 33876 12260
rect 33928 12248 33934 12300
rect 31665 12223 31723 12229
rect 31665 12220 31677 12223
rect 31444 12192 31677 12220
rect 31444 12180 31450 12192
rect 31665 12189 31677 12192
rect 31711 12189 31723 12223
rect 31665 12183 31723 12189
rect 31941 12223 31999 12229
rect 31941 12189 31953 12223
rect 31987 12189 31999 12223
rect 31941 12183 31999 12189
rect 32033 12223 32091 12229
rect 32033 12189 32045 12223
rect 32079 12220 32091 12223
rect 34422 12220 34428 12232
rect 32079 12192 34428 12220
rect 32079 12189 32091 12192
rect 32033 12183 32091 12189
rect 34422 12180 34428 12192
rect 34480 12180 34486 12232
rect 31849 12155 31907 12161
rect 31849 12152 31861 12155
rect 30208 12124 31861 12152
rect 31849 12121 31861 12124
rect 31895 12121 31907 12155
rect 31849 12115 31907 12121
rect 32858 12112 32864 12164
rect 32916 12152 32922 12164
rect 33137 12155 33195 12161
rect 33137 12152 33149 12155
rect 32916 12124 33149 12152
rect 32916 12112 32922 12124
rect 33137 12121 33149 12124
rect 33183 12121 33195 12155
rect 33137 12115 33195 12121
rect 24854 12084 24860 12096
rect 23676 12056 24860 12084
rect 24854 12044 24860 12056
rect 24912 12084 24918 12096
rect 25501 12087 25559 12093
rect 25501 12084 25513 12087
rect 24912 12056 25513 12084
rect 24912 12044 24918 12056
rect 25501 12053 25513 12056
rect 25547 12053 25559 12087
rect 25501 12047 25559 12053
rect 25866 12044 25872 12096
rect 25924 12044 25930 12096
rect 26418 12044 26424 12096
rect 26476 12084 26482 12096
rect 27522 12084 27528 12096
rect 26476 12056 27528 12084
rect 26476 12044 26482 12056
rect 27522 12044 27528 12056
rect 27580 12084 27586 12096
rect 27709 12087 27767 12093
rect 27709 12084 27721 12087
rect 27580 12056 27721 12084
rect 27580 12044 27586 12056
rect 27709 12053 27721 12056
rect 27755 12053 27767 12087
rect 27709 12047 27767 12053
rect 28258 12044 28264 12096
rect 28316 12044 28322 12096
rect 30926 12044 30932 12096
rect 30984 12084 30990 12096
rect 31205 12087 31263 12093
rect 31205 12084 31217 12087
rect 30984 12056 31217 12084
rect 30984 12044 30990 12056
rect 31205 12053 31217 12056
rect 31251 12053 31263 12087
rect 31205 12047 31263 12053
rect 1104 11994 35328 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35328 11994
rect 1104 11920 35328 11942
rect 7926 11840 7932 11892
rect 7984 11880 7990 11892
rect 11238 11880 11244 11892
rect 7984 11852 11244 11880
rect 7984 11840 7990 11852
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 11330 11840 11336 11892
rect 11388 11840 11394 11892
rect 13170 11840 13176 11892
rect 13228 11840 13234 11892
rect 13538 11840 13544 11892
rect 13596 11880 13602 11892
rect 14093 11883 14151 11889
rect 14093 11880 14105 11883
rect 13596 11852 14105 11880
rect 13596 11840 13602 11852
rect 14093 11849 14105 11852
rect 14139 11880 14151 11883
rect 16942 11880 16948 11892
rect 14139 11852 16948 11880
rect 14139 11849 14151 11852
rect 14093 11843 14151 11849
rect 16942 11840 16948 11852
rect 17000 11840 17006 11892
rect 17037 11883 17095 11889
rect 17037 11849 17049 11883
rect 17083 11880 17095 11883
rect 17126 11880 17132 11892
rect 17083 11852 17132 11880
rect 17083 11849 17095 11852
rect 17037 11843 17095 11849
rect 17126 11840 17132 11852
rect 17184 11840 17190 11892
rect 18414 11840 18420 11892
rect 18472 11880 18478 11892
rect 18969 11883 19027 11889
rect 18969 11880 18981 11883
rect 18472 11852 18981 11880
rect 18472 11840 18478 11852
rect 18969 11849 18981 11852
rect 19015 11849 19027 11883
rect 18969 11843 19027 11849
rect 20346 11840 20352 11892
rect 20404 11840 20410 11892
rect 20714 11840 20720 11892
rect 20772 11840 20778 11892
rect 20809 11883 20867 11889
rect 20809 11849 20821 11883
rect 20855 11880 20867 11883
rect 21082 11880 21088 11892
rect 20855 11852 21088 11880
rect 20855 11849 20867 11852
rect 20809 11843 20867 11849
rect 21082 11840 21088 11852
rect 21140 11840 21146 11892
rect 21192 11852 23428 11880
rect 3234 11812 3240 11824
rect 2884 11784 3240 11812
rect 2884 11753 2912 11784
rect 3234 11772 3240 11784
rect 3292 11812 3298 11824
rect 5534 11812 5540 11824
rect 3292 11784 5540 11812
rect 3292 11772 3298 11784
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11713 2927 11747
rect 2869 11707 2927 11713
rect 3136 11747 3194 11753
rect 3136 11713 3148 11747
rect 3182 11744 3194 11747
rect 3694 11744 3700 11756
rect 3182 11716 3700 11744
rect 3182 11713 3194 11716
rect 3136 11707 3194 11713
rect 3694 11704 3700 11716
rect 3752 11704 3758 11756
rect 4356 11753 4384 11784
rect 5534 11772 5540 11784
rect 5592 11772 5598 11824
rect 7024 11784 9996 11812
rect 4341 11747 4399 11753
rect 4341 11713 4353 11747
rect 4387 11713 4399 11747
rect 4341 11707 4399 11713
rect 4608 11747 4666 11753
rect 4608 11713 4620 11747
rect 4654 11744 4666 11747
rect 4890 11744 4896 11756
rect 4654 11716 4896 11744
rect 4654 11713 4666 11716
rect 4608 11707 4666 11713
rect 4890 11704 4896 11716
rect 4948 11704 4954 11756
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11744 6607 11747
rect 6730 11744 6736 11756
rect 6595 11716 6736 11744
rect 6595 11713 6607 11716
rect 6549 11707 6607 11713
rect 6730 11704 6736 11716
rect 6788 11744 6794 11756
rect 7024 11753 7052 11784
rect 7009 11747 7067 11753
rect 7009 11744 7021 11747
rect 6788 11716 7021 11744
rect 6788 11704 6794 11716
rect 7009 11713 7021 11716
rect 7055 11713 7067 11747
rect 7009 11707 7067 11713
rect 7276 11747 7334 11753
rect 7276 11713 7288 11747
rect 7322 11744 7334 11747
rect 7650 11744 7656 11756
rect 7322 11716 7656 11744
rect 7322 11713 7334 11716
rect 7276 11707 7334 11713
rect 7650 11704 7656 11716
rect 7708 11704 7714 11756
rect 8496 11753 8524 11784
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 8748 11747 8806 11753
rect 8748 11713 8760 11747
rect 8794 11744 8806 11747
rect 9306 11744 9312 11756
rect 8794 11716 9312 11744
rect 8794 11713 8806 11716
rect 8748 11707 8806 11713
rect 9306 11704 9312 11716
rect 9364 11704 9370 11756
rect 9968 11753 9996 11784
rect 11146 11772 11152 11824
rect 11204 11812 11210 11824
rect 11204 11784 12480 11812
rect 11204 11772 11210 11784
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11713 10011 11747
rect 9953 11707 10011 11713
rect 10220 11747 10278 11753
rect 10220 11713 10232 11747
rect 10266 11744 10278 11747
rect 10962 11744 10968 11756
rect 10266 11716 10968 11744
rect 10266 11713 10278 11716
rect 10220 11707 10278 11713
rect 10962 11704 10968 11716
rect 11020 11704 11026 11756
rect 12060 11747 12118 11753
rect 12060 11713 12072 11747
rect 12106 11744 12118 11747
rect 12342 11744 12348 11756
rect 12106 11716 12348 11744
rect 12106 11713 12118 11716
rect 12060 11707 12118 11713
rect 12342 11704 12348 11716
rect 12400 11704 12406 11756
rect 12452 11744 12480 11784
rect 12526 11772 12532 11824
rect 12584 11812 12590 11824
rect 15289 11815 15347 11821
rect 15289 11812 15301 11815
rect 12584 11784 15301 11812
rect 12584 11772 12590 11784
rect 15289 11781 15301 11784
rect 15335 11812 15347 11815
rect 15470 11812 15476 11824
rect 15335 11784 15476 11812
rect 15335 11781 15347 11784
rect 15289 11775 15347 11781
rect 15470 11772 15476 11784
rect 15528 11812 15534 11824
rect 15528 11784 17632 11812
rect 15528 11772 15534 11784
rect 14642 11744 14648 11756
rect 12452 11716 14648 11744
rect 14642 11704 14648 11716
rect 14700 11704 14706 11756
rect 14737 11747 14795 11753
rect 14737 11713 14749 11747
rect 14783 11713 14795 11747
rect 14737 11707 14795 11713
rect 11793 11679 11851 11685
rect 11793 11645 11805 11679
rect 11839 11645 11851 11679
rect 11793 11639 11851 11645
rect 7944 11580 8524 11608
rect 4249 11543 4307 11549
rect 4249 11509 4261 11543
rect 4295 11540 4307 11543
rect 4614 11540 4620 11552
rect 4295 11512 4620 11540
rect 4295 11509 4307 11512
rect 4249 11503 4307 11509
rect 4614 11500 4620 11512
rect 4672 11500 4678 11552
rect 5258 11500 5264 11552
rect 5316 11540 5322 11552
rect 5721 11543 5779 11549
rect 5721 11540 5733 11543
rect 5316 11512 5733 11540
rect 5316 11500 5322 11512
rect 5721 11509 5733 11512
rect 5767 11509 5779 11543
rect 5721 11503 5779 11509
rect 6086 11500 6092 11552
rect 6144 11540 6150 11552
rect 7944 11540 7972 11580
rect 6144 11512 7972 11540
rect 6144 11500 6150 11512
rect 8386 11500 8392 11552
rect 8444 11500 8450 11552
rect 8496 11540 8524 11580
rect 9416 11580 9996 11608
rect 9416 11540 9444 11580
rect 8496 11512 9444 11540
rect 9766 11500 9772 11552
rect 9824 11540 9830 11552
rect 9861 11543 9919 11549
rect 9861 11540 9873 11543
rect 9824 11512 9873 11540
rect 9824 11500 9830 11512
rect 9861 11509 9873 11512
rect 9907 11509 9919 11543
rect 9968 11540 9996 11580
rect 10318 11540 10324 11552
rect 9968 11512 10324 11540
rect 9861 11503 9919 11509
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 11808 11540 11836 11639
rect 13906 11636 13912 11688
rect 13964 11676 13970 11688
rect 14752 11676 14780 11707
rect 14918 11704 14924 11756
rect 14976 11704 14982 11756
rect 15013 11747 15071 11753
rect 15013 11713 15025 11747
rect 15059 11744 15071 11747
rect 16117 11747 16175 11753
rect 16117 11744 16129 11747
rect 15059 11716 16129 11744
rect 15059 11713 15071 11716
rect 15013 11707 15071 11713
rect 16117 11713 16129 11716
rect 16163 11744 16175 11747
rect 16574 11744 16580 11756
rect 16163 11716 16580 11744
rect 16163 11713 16175 11716
rect 16117 11707 16175 11713
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 17129 11747 17187 11753
rect 17129 11713 17141 11747
rect 17175 11744 17187 11747
rect 17310 11744 17316 11756
rect 17175 11716 17316 11744
rect 17175 11713 17187 11716
rect 17129 11707 17187 11713
rect 17310 11704 17316 11716
rect 17368 11744 17374 11756
rect 17494 11744 17500 11756
rect 17368 11716 17500 11744
rect 17368 11704 17374 11716
rect 17494 11704 17500 11716
rect 17552 11704 17558 11756
rect 17604 11753 17632 11784
rect 17678 11772 17684 11824
rect 17736 11812 17742 11824
rect 21192 11812 21220 11852
rect 22462 11812 22468 11824
rect 17736 11784 21220 11812
rect 21836 11784 22468 11812
rect 17736 11772 17742 11784
rect 17862 11753 17868 11756
rect 17589 11747 17647 11753
rect 17589 11713 17601 11747
rect 17635 11713 17647 11747
rect 17589 11707 17647 11713
rect 17856 11707 17868 11753
rect 17862 11704 17868 11707
rect 17920 11704 17926 11756
rect 13964 11648 14780 11676
rect 13964 11636 13970 11648
rect 16666 11636 16672 11688
rect 16724 11676 16730 11688
rect 17221 11679 17279 11685
rect 17221 11676 17233 11679
rect 16724 11648 17233 11676
rect 16724 11636 16730 11648
rect 17221 11645 17233 11648
rect 17267 11676 17279 11679
rect 17267 11648 17632 11676
rect 17267 11645 17279 11648
rect 17221 11639 17279 11645
rect 17604 11620 17632 11648
rect 20070 11636 20076 11688
rect 20128 11676 20134 11688
rect 20257 11679 20315 11685
rect 20257 11676 20269 11679
rect 20128 11648 20269 11676
rect 20128 11636 20134 11648
rect 20257 11645 20269 11648
rect 20303 11676 20315 11679
rect 20993 11679 21051 11685
rect 20993 11676 21005 11679
rect 20303 11648 21005 11676
rect 20303 11645 20315 11648
rect 20257 11639 20315 11645
rect 20993 11645 21005 11648
rect 21039 11676 21051 11679
rect 21358 11676 21364 11688
rect 21039 11648 21364 11676
rect 21039 11645 21051 11648
rect 20993 11639 21051 11645
rect 21358 11636 21364 11648
rect 21416 11636 21422 11688
rect 21836 11685 21864 11784
rect 22462 11772 22468 11784
rect 22520 11772 22526 11824
rect 22094 11753 22100 11756
rect 22088 11707 22100 11753
rect 22094 11704 22100 11707
rect 22152 11704 22158 11756
rect 23400 11744 23428 11852
rect 23474 11840 23480 11892
rect 23532 11840 23538 11892
rect 23842 11840 23848 11892
rect 23900 11840 23906 11892
rect 25038 11840 25044 11892
rect 25096 11880 25102 11892
rect 25593 11883 25651 11889
rect 25593 11880 25605 11883
rect 25096 11852 25605 11880
rect 25096 11840 25102 11852
rect 25593 11849 25605 11852
rect 25639 11880 25651 11883
rect 25866 11880 25872 11892
rect 25639 11852 25872 11880
rect 25639 11849 25651 11852
rect 25593 11843 25651 11849
rect 25866 11840 25872 11852
rect 25924 11880 25930 11892
rect 26605 11883 26663 11889
rect 26605 11880 26617 11883
rect 25924 11852 26617 11880
rect 25924 11840 25930 11852
rect 26605 11849 26617 11852
rect 26651 11849 26663 11883
rect 26605 11843 26663 11849
rect 27246 11840 27252 11892
rect 27304 11880 27310 11892
rect 27304 11852 29684 11880
rect 27304 11840 27310 11852
rect 23658 11772 23664 11824
rect 23716 11812 23722 11824
rect 23716 11784 25176 11812
rect 23716 11772 23722 11784
rect 24305 11747 24363 11753
rect 23400 11716 24072 11744
rect 21821 11679 21879 11685
rect 21821 11645 21833 11679
rect 21867 11645 21879 11679
rect 21821 11639 21879 11645
rect 15933 11611 15991 11617
rect 15933 11608 15945 11611
rect 14752 11580 15945 11608
rect 12526 11540 12532 11552
rect 11808 11512 12532 11540
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 12710 11500 12716 11552
rect 12768 11540 12774 11552
rect 13538 11540 13544 11552
rect 12768 11512 13544 11540
rect 12768 11500 12774 11512
rect 13538 11500 13544 11512
rect 13596 11500 13602 11552
rect 14642 11500 14648 11552
rect 14700 11540 14706 11552
rect 14752 11540 14780 11580
rect 15933 11577 15945 11580
rect 15979 11608 15991 11611
rect 16942 11608 16948 11620
rect 15979 11580 16948 11608
rect 15979 11577 15991 11580
rect 15933 11571 15991 11577
rect 16942 11568 16948 11580
rect 17000 11568 17006 11620
rect 17586 11568 17592 11620
rect 17644 11568 17650 11620
rect 20346 11568 20352 11620
rect 20404 11608 20410 11620
rect 21836 11608 21864 11639
rect 23934 11636 23940 11688
rect 23992 11636 23998 11688
rect 24044 11685 24072 11716
rect 24305 11713 24317 11747
rect 24351 11744 24363 11747
rect 24670 11744 24676 11756
rect 24351 11716 24676 11744
rect 24351 11713 24363 11716
rect 24305 11707 24363 11713
rect 24670 11704 24676 11716
rect 24728 11744 24734 11756
rect 24728 11716 24992 11744
rect 24728 11704 24734 11716
rect 24029 11679 24087 11685
rect 24029 11645 24041 11679
rect 24075 11676 24087 11679
rect 24964 11676 24992 11716
rect 25038 11704 25044 11756
rect 25096 11704 25102 11756
rect 25148 11744 25176 11784
rect 26142 11772 26148 11824
rect 26200 11812 26206 11824
rect 27617 11815 27675 11821
rect 27617 11812 27629 11815
rect 26200 11784 27629 11812
rect 26200 11772 26206 11784
rect 27617 11781 27629 11784
rect 27663 11812 27675 11815
rect 27663 11784 27844 11812
rect 27663 11781 27675 11784
rect 27617 11775 27675 11781
rect 25409 11747 25467 11753
rect 25409 11744 25421 11747
rect 25148 11716 25421 11744
rect 25409 11713 25421 11716
rect 25455 11713 25467 11747
rect 25409 11707 25467 11713
rect 25961 11747 26019 11753
rect 25961 11713 25973 11747
rect 26007 11713 26019 11747
rect 25961 11707 26019 11713
rect 26237 11747 26295 11753
rect 26237 11713 26249 11747
rect 26283 11713 26295 11747
rect 26237 11707 26295 11713
rect 26329 11747 26387 11753
rect 26329 11713 26341 11747
rect 26375 11744 26387 11747
rect 26375 11716 26464 11744
rect 26375 11713 26387 11716
rect 26329 11707 26387 11713
rect 25777 11679 25835 11685
rect 25777 11676 25789 11679
rect 24075 11648 24532 11676
rect 24964 11648 25789 11676
rect 24075 11645 24087 11648
rect 24029 11639 24087 11645
rect 20404 11580 21864 11608
rect 23201 11611 23259 11617
rect 20404 11568 20410 11580
rect 23201 11577 23213 11611
rect 23247 11608 23259 11611
rect 23290 11608 23296 11620
rect 23247 11580 23296 11608
rect 23247 11577 23259 11580
rect 23201 11571 23259 11577
rect 23290 11568 23296 11580
rect 23348 11568 23354 11620
rect 23952 11608 23980 11636
rect 24394 11608 24400 11620
rect 23952 11580 24400 11608
rect 24394 11568 24400 11580
rect 24452 11568 24458 11620
rect 24504 11617 24532 11648
rect 25777 11645 25789 11648
rect 25823 11645 25835 11679
rect 25777 11639 25835 11645
rect 24489 11611 24547 11617
rect 24489 11577 24501 11611
rect 24535 11608 24547 11611
rect 24673 11611 24731 11617
rect 24673 11608 24685 11611
rect 24535 11580 24685 11608
rect 24535 11577 24547 11580
rect 24489 11571 24547 11577
rect 24673 11577 24685 11580
rect 24719 11608 24731 11611
rect 24857 11611 24915 11617
rect 24857 11608 24869 11611
rect 24719 11580 24869 11608
rect 24719 11577 24731 11580
rect 24673 11571 24731 11577
rect 24857 11577 24869 11580
rect 24903 11577 24915 11611
rect 25976 11608 26004 11707
rect 26050 11636 26056 11688
rect 26108 11676 26114 11688
rect 26252 11676 26280 11707
rect 26108 11648 26280 11676
rect 26436 11676 26464 11716
rect 26510 11704 26516 11756
rect 26568 11744 26574 11756
rect 27065 11747 27123 11753
rect 27065 11744 27077 11747
rect 26568 11716 27077 11744
rect 26568 11704 26574 11716
rect 27065 11713 27077 11716
rect 27111 11713 27123 11747
rect 27065 11707 27123 11713
rect 27706 11704 27712 11756
rect 27764 11704 27770 11756
rect 27816 11744 27844 11784
rect 28166 11772 28172 11824
rect 28224 11812 28230 11824
rect 29549 11815 29607 11821
rect 29549 11812 29561 11815
rect 28224 11784 29561 11812
rect 28224 11772 28230 11784
rect 29549 11781 29561 11784
rect 29595 11781 29607 11815
rect 29656 11812 29684 11852
rect 30098 11840 30104 11892
rect 30156 11840 30162 11892
rect 31386 11840 31392 11892
rect 31444 11840 31450 11892
rect 31478 11840 31484 11892
rect 31536 11840 31542 11892
rect 31496 11812 31524 11840
rect 29656 11784 30328 11812
rect 29549 11775 29607 11781
rect 30300 11756 30328 11784
rect 31036 11784 31524 11812
rect 28718 11744 28724 11756
rect 27816 11716 28724 11744
rect 28718 11704 28724 11716
rect 28776 11704 28782 11756
rect 29086 11704 29092 11756
rect 29144 11753 29150 11756
rect 29144 11707 29156 11753
rect 29144 11704 29150 11707
rect 30282 11704 30288 11756
rect 30340 11744 30346 11756
rect 30469 11747 30527 11753
rect 30469 11744 30481 11747
rect 30340 11716 30481 11744
rect 30340 11704 30346 11716
rect 30469 11713 30481 11716
rect 30515 11713 30527 11747
rect 30469 11707 30527 11713
rect 30561 11747 30619 11753
rect 30561 11713 30573 11747
rect 30607 11744 30619 11747
rect 30926 11744 30932 11756
rect 30607 11716 30932 11744
rect 30607 11713 30619 11716
rect 30561 11707 30619 11713
rect 30926 11704 30932 11716
rect 30984 11704 30990 11756
rect 31036 11753 31064 11784
rect 31021 11747 31079 11753
rect 31021 11713 31033 11747
rect 31067 11713 31079 11747
rect 31021 11707 31079 11713
rect 31205 11747 31263 11753
rect 31205 11713 31217 11747
rect 31251 11744 31263 11747
rect 31294 11744 31300 11756
rect 31251 11716 31300 11744
rect 31251 11713 31263 11716
rect 31205 11707 31263 11713
rect 31294 11704 31300 11716
rect 31352 11704 31358 11756
rect 34514 11704 34520 11756
rect 34572 11704 34578 11756
rect 26786 11676 26792 11688
rect 26436 11648 26792 11676
rect 26108 11636 26114 11648
rect 26786 11636 26792 11648
rect 26844 11676 26850 11688
rect 27341 11679 27399 11685
rect 27341 11676 27353 11679
rect 26844 11648 27353 11676
rect 26844 11636 26850 11648
rect 27341 11645 27353 11648
rect 27387 11645 27399 11679
rect 27341 11639 27399 11645
rect 27614 11636 27620 11688
rect 27672 11676 27678 11688
rect 28350 11676 28356 11688
rect 27672 11648 28356 11676
rect 27672 11636 27678 11648
rect 28350 11636 28356 11648
rect 28408 11636 28414 11688
rect 29365 11679 29423 11685
rect 29365 11645 29377 11679
rect 29411 11676 29423 11679
rect 29822 11676 29828 11688
rect 29411 11648 29828 11676
rect 29411 11645 29423 11648
rect 29365 11639 29423 11645
rect 29822 11636 29828 11648
rect 29880 11636 29886 11688
rect 30650 11636 30656 11688
rect 30708 11636 30714 11688
rect 34790 11636 34796 11688
rect 34848 11636 34854 11688
rect 27982 11608 27988 11620
rect 25976 11580 27988 11608
rect 24857 11571 24915 11577
rect 27982 11568 27988 11580
rect 28040 11568 28046 11620
rect 30668 11608 30696 11636
rect 29380 11580 30696 11608
rect 14700 11512 14780 11540
rect 14700 11500 14706 11512
rect 15194 11500 15200 11552
rect 15252 11500 15258 11552
rect 16666 11500 16672 11552
rect 16724 11500 16730 11552
rect 20714 11500 20720 11552
rect 20772 11540 20778 11552
rect 22554 11540 22560 11552
rect 20772 11512 22560 11540
rect 20772 11500 20778 11512
rect 22554 11500 22560 11512
rect 22612 11500 22618 11552
rect 25225 11543 25283 11549
rect 25225 11509 25237 11543
rect 25271 11540 25283 11543
rect 25498 11540 25504 11552
rect 25271 11512 25504 11540
rect 25271 11509 25283 11512
rect 25225 11503 25283 11509
rect 25498 11500 25504 11512
rect 25556 11500 25562 11552
rect 26510 11500 26516 11552
rect 26568 11500 26574 11552
rect 26694 11500 26700 11552
rect 26752 11540 26758 11552
rect 29380 11540 29408 11580
rect 26752 11512 29408 11540
rect 26752 11500 26758 11512
rect 29546 11500 29552 11552
rect 29604 11540 29610 11552
rect 29641 11543 29699 11549
rect 29641 11540 29653 11543
rect 29604 11512 29653 11540
rect 29604 11500 29610 11512
rect 29641 11509 29653 11512
rect 29687 11540 29699 11543
rect 29825 11543 29883 11549
rect 29825 11540 29837 11543
rect 29687 11512 29837 11540
rect 29687 11509 29699 11512
rect 29641 11503 29699 11509
rect 29825 11509 29837 11512
rect 29871 11509 29883 11543
rect 29825 11503 29883 11509
rect 1104 11450 35328 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 35328 11450
rect 1104 11376 35328 11398
rect 3694 11296 3700 11348
rect 3752 11336 3758 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 3752 11308 3801 11336
rect 3752 11296 3758 11308
rect 3789 11305 3801 11308
rect 3835 11305 3847 11339
rect 3789 11299 3847 11305
rect 4890 11296 4896 11348
rect 4948 11296 4954 11348
rect 5736 11308 7328 11336
rect 5074 11268 5080 11280
rect 4264 11240 5080 11268
rect 4264 11212 4292 11240
rect 5074 11228 5080 11240
rect 5132 11228 5138 11280
rect 2961 11203 3019 11209
rect 2961 11169 2973 11203
rect 3007 11200 3019 11203
rect 3329 11203 3387 11209
rect 3329 11200 3341 11203
rect 3007 11172 3341 11200
rect 3007 11169 3019 11172
rect 2961 11163 3019 11169
rect 3329 11169 3341 11172
rect 3375 11200 3387 11203
rect 3605 11203 3663 11209
rect 3605 11200 3617 11203
rect 3375 11172 3617 11200
rect 3375 11169 3387 11172
rect 3329 11163 3387 11169
rect 3605 11169 3617 11172
rect 3651 11200 3663 11203
rect 4246 11200 4252 11212
rect 3651 11172 4252 11200
rect 3651 11169 3663 11172
rect 3605 11163 3663 11169
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 5736 11209 5764 11308
rect 5997 11271 6055 11277
rect 5997 11237 6009 11271
rect 6043 11268 6055 11271
rect 6086 11268 6092 11280
rect 6043 11240 6092 11268
rect 6043 11237 6055 11240
rect 5997 11231 6055 11237
rect 4433 11203 4491 11209
rect 4433 11169 4445 11203
rect 4479 11200 4491 11203
rect 5537 11203 5595 11209
rect 4479 11172 5488 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 1302 11092 1308 11144
rect 1360 11132 1366 11144
rect 1397 11135 1455 11141
rect 1397 11132 1409 11135
rect 1360 11104 1409 11132
rect 1360 11092 1366 11104
rect 1397 11101 1409 11104
rect 1443 11132 1455 11135
rect 1673 11135 1731 11141
rect 1673 11132 1685 11135
rect 1443 11104 1685 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 1673 11101 1685 11104
rect 1719 11101 1731 11135
rect 1673 11095 1731 11101
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4614 11132 4620 11144
rect 4203 11104 4620 11132
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 4801 11135 4859 11141
rect 4801 11101 4813 11135
rect 4847 11132 4859 11135
rect 4847 11104 5120 11132
rect 4847 11101 4859 11104
rect 4801 11095 4859 11101
rect 5092 11076 5120 11104
rect 5258 11092 5264 11144
rect 5316 11092 5322 11144
rect 5460 11132 5488 11172
rect 5537 11169 5549 11203
rect 5583 11200 5595 11203
rect 5721 11203 5779 11209
rect 5721 11200 5733 11203
rect 5583 11172 5733 11200
rect 5583 11169 5595 11172
rect 5537 11163 5595 11169
rect 5721 11169 5733 11172
rect 5767 11169 5779 11203
rect 5721 11163 5779 11169
rect 6012 11132 6040 11231
rect 6086 11228 6092 11240
rect 6144 11228 6150 11280
rect 5460 11104 6040 11132
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11132 6147 11135
rect 6730 11132 6736 11144
rect 6135 11104 6736 11132
rect 6135 11101 6147 11104
rect 6089 11095 6147 11101
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 3142 11064 3148 11076
rect 1596 11036 3148 11064
rect 1596 11005 1624 11036
rect 3142 11024 3148 11036
rect 3200 11024 3206 11076
rect 5074 11024 5080 11076
rect 5132 11064 5138 11076
rect 5353 11067 5411 11073
rect 5353 11064 5365 11067
rect 5132 11036 5365 11064
rect 5132 11024 5138 11036
rect 5353 11033 5365 11036
rect 5399 11033 5411 11067
rect 5353 11027 5411 11033
rect 6356 11067 6414 11073
rect 6356 11033 6368 11067
rect 6402 11064 6414 11067
rect 7006 11064 7012 11076
rect 6402 11036 7012 11064
rect 6402 11033 6414 11036
rect 6356 11027 6414 11033
rect 7006 11024 7012 11036
rect 7064 11024 7070 11076
rect 7300 11064 7328 11308
rect 7374 11296 7380 11348
rect 7432 11336 7438 11348
rect 7469 11339 7527 11345
rect 7469 11336 7481 11339
rect 7432 11308 7481 11336
rect 7432 11296 7438 11308
rect 7469 11305 7481 11308
rect 7515 11305 7527 11339
rect 7469 11299 7527 11305
rect 7650 11296 7656 11348
rect 7708 11296 7714 11348
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 9401 11339 9459 11345
rect 9401 11336 9413 11339
rect 9364 11308 9413 11336
rect 9364 11296 9370 11308
rect 9401 11305 9413 11308
rect 9447 11305 9459 11339
rect 10410 11336 10416 11348
rect 9401 11299 9459 11305
rect 9508 11308 10416 11336
rect 7466 11160 7472 11212
rect 7524 11200 7530 11212
rect 8113 11203 8171 11209
rect 8113 11200 8125 11203
rect 7524 11172 8125 11200
rect 7524 11160 7530 11172
rect 8113 11169 8125 11172
rect 8159 11169 8171 11203
rect 8113 11163 8171 11169
rect 8202 11160 8208 11212
rect 8260 11200 8266 11212
rect 8481 11203 8539 11209
rect 8481 11200 8493 11203
rect 8260 11172 8493 11200
rect 8260 11160 8266 11172
rect 8481 11169 8493 11172
rect 8527 11169 8539 11203
rect 8481 11163 8539 11169
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11132 8079 11135
rect 8386 11132 8392 11144
rect 8067 11104 8392 11132
rect 8067 11101 8079 11104
rect 8021 11095 8079 11101
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 9508 11064 9536 11308
rect 10410 11296 10416 11308
rect 10468 11336 10474 11348
rect 10870 11336 10876 11348
rect 10468 11308 10876 11336
rect 10468 11296 10474 11308
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 10962 11296 10968 11348
rect 11020 11296 11026 11348
rect 12342 11296 12348 11348
rect 12400 11296 12406 11348
rect 13906 11296 13912 11348
rect 13964 11296 13970 11348
rect 14461 11339 14519 11345
rect 14461 11305 14473 11339
rect 14507 11336 14519 11339
rect 14918 11336 14924 11348
rect 14507 11308 14924 11336
rect 14507 11305 14519 11308
rect 14461 11299 14519 11305
rect 14918 11296 14924 11308
rect 14976 11336 14982 11348
rect 16114 11336 16120 11348
rect 14976 11308 16120 11336
rect 14976 11296 14982 11308
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 17126 11296 17132 11348
rect 17184 11336 17190 11348
rect 17313 11339 17371 11345
rect 17313 11336 17325 11339
rect 17184 11308 17325 11336
rect 17184 11296 17190 11308
rect 17313 11305 17325 11308
rect 17359 11305 17371 11339
rect 17313 11299 17371 11305
rect 17586 11296 17592 11348
rect 17644 11296 17650 11348
rect 17862 11296 17868 11348
rect 17920 11336 17926 11348
rect 18049 11339 18107 11345
rect 18049 11336 18061 11339
rect 17920 11308 18061 11336
rect 17920 11296 17926 11308
rect 18049 11305 18061 11308
rect 18095 11305 18107 11339
rect 18049 11299 18107 11305
rect 18969 11339 19027 11345
rect 18969 11305 18981 11339
rect 19015 11336 19027 11339
rect 19610 11336 19616 11348
rect 19015 11308 19616 11336
rect 19015 11305 19027 11308
rect 18969 11299 19027 11305
rect 19610 11296 19616 11308
rect 19668 11296 19674 11348
rect 20990 11296 20996 11348
rect 21048 11336 21054 11348
rect 21177 11339 21235 11345
rect 21177 11336 21189 11339
rect 21048 11308 21189 11336
rect 21048 11296 21054 11308
rect 21177 11305 21189 11308
rect 21223 11336 21235 11339
rect 21453 11339 21511 11345
rect 21453 11336 21465 11339
rect 21223 11308 21465 11336
rect 21223 11305 21235 11308
rect 21177 11299 21235 11305
rect 21453 11305 21465 11308
rect 21499 11336 21511 11339
rect 21726 11336 21732 11348
rect 21499 11308 21732 11336
rect 21499 11305 21511 11308
rect 21453 11299 21511 11305
rect 21726 11296 21732 11308
rect 21784 11296 21790 11348
rect 22094 11296 22100 11348
rect 22152 11336 22158 11348
rect 22189 11339 22247 11345
rect 22189 11336 22201 11339
rect 22152 11308 22201 11336
rect 22152 11296 22158 11308
rect 22189 11305 22201 11308
rect 22235 11305 22247 11339
rect 25777 11339 25835 11345
rect 22189 11299 22247 11305
rect 24412 11308 25728 11336
rect 12710 11268 12716 11280
rect 10428 11240 12716 11268
rect 9674 11160 9680 11212
rect 9732 11200 9738 11212
rect 9861 11203 9919 11209
rect 9861 11200 9873 11203
rect 9732 11172 9873 11200
rect 9732 11160 9738 11172
rect 9861 11169 9873 11172
rect 9907 11169 9919 11203
rect 9861 11163 9919 11169
rect 10042 11160 10048 11212
rect 10100 11160 10106 11212
rect 10134 11160 10140 11212
rect 10192 11200 10198 11212
rect 10428 11200 10456 11240
rect 12710 11228 12716 11240
rect 12768 11228 12774 11280
rect 16942 11228 16948 11280
rect 17000 11268 17006 11280
rect 24412 11268 24440 11308
rect 17000 11240 24440 11268
rect 25700 11268 25728 11308
rect 25777 11305 25789 11339
rect 25823 11336 25835 11339
rect 26050 11336 26056 11348
rect 25823 11308 26056 11336
rect 25823 11305 25835 11308
rect 25777 11299 25835 11305
rect 26050 11296 26056 11308
rect 26108 11296 26114 11348
rect 26326 11296 26332 11348
rect 26384 11296 26390 11348
rect 26510 11296 26516 11348
rect 26568 11336 26574 11348
rect 26697 11339 26755 11345
rect 26697 11336 26709 11339
rect 26568 11308 26709 11336
rect 26568 11296 26574 11308
rect 26697 11305 26709 11308
rect 26743 11305 26755 11339
rect 26697 11299 26755 11305
rect 26789 11339 26847 11345
rect 26789 11305 26801 11339
rect 26835 11336 26847 11339
rect 28534 11336 28540 11348
rect 26835 11308 28540 11336
rect 26835 11305 26847 11308
rect 26789 11299 26847 11305
rect 28534 11296 28540 11308
rect 28592 11296 28598 11348
rect 29086 11296 29092 11348
rect 29144 11296 29150 11348
rect 30561 11339 30619 11345
rect 30561 11305 30573 11339
rect 30607 11336 30619 11339
rect 30650 11336 30656 11348
rect 30607 11308 30656 11336
rect 30607 11305 30619 11308
rect 30561 11299 30619 11305
rect 30650 11296 30656 11308
rect 30708 11296 30714 11348
rect 26605 11271 26663 11277
rect 26605 11268 26617 11271
rect 25700 11240 26617 11268
rect 17000 11228 17006 11240
rect 26605 11237 26617 11240
rect 26651 11268 26663 11271
rect 27433 11271 27491 11277
rect 27433 11268 27445 11271
rect 26651 11240 27445 11268
rect 26651 11237 26663 11240
rect 26605 11231 26663 11237
rect 27433 11237 27445 11240
rect 27479 11268 27491 11271
rect 27706 11268 27712 11280
rect 27479 11240 27712 11268
rect 27479 11237 27491 11240
rect 27433 11231 27491 11237
rect 27706 11228 27712 11240
rect 27764 11268 27770 11280
rect 29181 11271 29239 11277
rect 29181 11268 29193 11271
rect 27764 11240 29193 11268
rect 27764 11228 27770 11240
rect 29181 11237 29193 11240
rect 29227 11237 29239 11271
rect 29181 11231 29239 11237
rect 10192 11172 10456 11200
rect 10192 11160 10198 11172
rect 10428 11144 10456 11172
rect 11238 11160 11244 11212
rect 11296 11200 11302 11212
rect 11609 11203 11667 11209
rect 11609 11200 11621 11203
rect 11296 11172 11621 11200
rect 11296 11160 11302 11172
rect 11609 11169 11621 11172
rect 11655 11200 11667 11203
rect 11885 11203 11943 11209
rect 11885 11200 11897 11203
rect 11655 11172 11897 11200
rect 11655 11169 11667 11172
rect 11609 11163 11667 11169
rect 11885 11169 11897 11172
rect 11931 11200 11943 11203
rect 12802 11200 12808 11212
rect 11931 11172 12808 11200
rect 11931 11169 11943 11172
rect 11885 11163 11943 11169
rect 12802 11160 12808 11172
rect 12860 11160 12866 11212
rect 12989 11203 13047 11209
rect 12989 11169 13001 11203
rect 13035 11200 13047 11203
rect 13265 11203 13323 11209
rect 13265 11200 13277 11203
rect 13035 11172 13277 11200
rect 13035 11169 13047 11172
rect 12989 11163 13047 11169
rect 13265 11169 13277 11172
rect 13311 11200 13323 11203
rect 13311 11172 14320 11200
rect 13311 11169 13323 11172
rect 13265 11163 13323 11169
rect 9766 11092 9772 11144
rect 9824 11092 9830 11144
rect 10226 11092 10232 11144
rect 10284 11092 10290 11144
rect 10410 11092 10416 11144
rect 10468 11092 10474 11144
rect 10505 11135 10563 11141
rect 10505 11101 10517 11135
rect 10551 11101 10563 11135
rect 10505 11095 10563 11101
rect 7300 11036 9536 11064
rect 9784 11064 9812 11092
rect 10520 11064 10548 11095
rect 10686 11092 10692 11144
rect 10744 11092 10750 11144
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11132 10839 11135
rect 11146 11132 11152 11144
rect 10827 11104 11152 11132
rect 10827 11101 10839 11104
rect 10781 11095 10839 11101
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 11330 11092 11336 11144
rect 11388 11092 11394 11144
rect 12713 11135 12771 11141
rect 12713 11101 12725 11135
rect 12759 11132 12771 11135
rect 13170 11132 13176 11144
rect 12759 11104 13176 11132
rect 12759 11101 12771 11104
rect 12713 11095 12771 11101
rect 13170 11092 13176 11104
rect 13228 11092 13234 11144
rect 13354 11092 13360 11144
rect 13412 11092 13418 11144
rect 13538 11092 13544 11144
rect 13596 11092 13602 11144
rect 13722 11092 13728 11144
rect 13780 11132 13786 11144
rect 14185 11135 14243 11141
rect 14185 11132 14197 11135
rect 13780 11104 14197 11132
rect 13780 11092 13786 11104
rect 14185 11101 14197 11104
rect 14231 11101 14243 11135
rect 14292 11132 14320 11172
rect 17310 11160 17316 11212
rect 17368 11200 17374 11212
rect 18509 11203 18567 11209
rect 18509 11200 18521 11203
rect 17368 11172 18521 11200
rect 17368 11160 17374 11172
rect 18509 11169 18521 11172
rect 18555 11169 18567 11203
rect 18509 11163 18567 11169
rect 18693 11203 18751 11209
rect 18693 11169 18705 11203
rect 18739 11200 18751 11203
rect 19610 11200 19616 11212
rect 18739 11172 19616 11200
rect 18739 11169 18751 11172
rect 18693 11163 18751 11169
rect 19610 11160 19616 11172
rect 19668 11160 19674 11212
rect 22094 11160 22100 11212
rect 22152 11200 22158 11212
rect 22741 11203 22799 11209
rect 22741 11200 22753 11203
rect 22152 11172 22753 11200
rect 22152 11160 22158 11172
rect 22741 11169 22753 11172
rect 22787 11169 22799 11203
rect 22741 11163 22799 11169
rect 22922 11160 22928 11212
rect 22980 11200 22986 11212
rect 24397 11203 24455 11209
rect 24397 11200 24409 11203
rect 22980 11172 24409 11200
rect 22980 11160 22986 11172
rect 24397 11169 24409 11172
rect 24443 11169 24455 11203
rect 24397 11163 24455 11169
rect 26237 11203 26295 11209
rect 26237 11169 26249 11203
rect 26283 11200 26295 11203
rect 27614 11200 27620 11212
rect 26283 11172 27620 11200
rect 26283 11169 26295 11172
rect 26237 11163 26295 11169
rect 15102 11132 15108 11144
rect 14292 11104 15108 11132
rect 14185 11095 14243 11101
rect 15102 11092 15108 11104
rect 15160 11092 15166 11144
rect 15841 11135 15899 11141
rect 15841 11132 15853 11135
rect 15488 11104 15853 11132
rect 15488 11076 15516 11104
rect 15841 11101 15853 11104
rect 15887 11132 15899 11135
rect 15933 11135 15991 11141
rect 15933 11132 15945 11135
rect 15887 11104 15945 11132
rect 15887 11101 15899 11104
rect 15841 11095 15899 11101
rect 15933 11101 15945 11104
rect 15979 11101 15991 11135
rect 15933 11095 15991 11101
rect 16200 11135 16258 11141
rect 16200 11101 16212 11135
rect 16246 11132 16258 11135
rect 16666 11132 16672 11144
rect 16246 11104 16672 11132
rect 16246 11101 16258 11104
rect 16200 11095 16258 11101
rect 16666 11092 16672 11104
rect 16724 11092 16730 11144
rect 18414 11092 18420 11144
rect 18472 11092 18478 11144
rect 19797 11135 19855 11141
rect 19797 11101 19809 11135
rect 19843 11101 19855 11135
rect 19797 11095 19855 11101
rect 21361 11135 21419 11141
rect 21361 11101 21373 11135
rect 21407 11132 21419 11135
rect 22462 11132 22468 11144
rect 21407 11104 22468 11132
rect 21407 11101 21419 11104
rect 21361 11095 21419 11101
rect 9784 11036 10548 11064
rect 11425 11067 11483 11073
rect 11425 11033 11437 11067
rect 11471 11064 11483 11067
rect 12434 11064 12440 11076
rect 11471 11036 12440 11064
rect 11471 11033 11483 11036
rect 11425 11027 11483 11033
rect 12434 11024 12440 11036
rect 12492 11064 12498 11076
rect 12805 11067 12863 11073
rect 12805 11064 12817 11067
rect 12492 11036 12817 11064
rect 12492 11024 12498 11036
rect 12805 11033 12817 11036
rect 12851 11033 12863 11067
rect 12805 11027 12863 11033
rect 13633 11067 13691 11073
rect 13633 11033 13645 11067
rect 13679 11064 13691 11067
rect 13906 11064 13912 11076
rect 13679 11036 13912 11064
rect 13679 11033 13691 11036
rect 13633 11027 13691 11033
rect 13906 11024 13912 11036
rect 13964 11024 13970 11076
rect 15470 11024 15476 11076
rect 15528 11024 15534 11076
rect 15596 11067 15654 11073
rect 15596 11033 15608 11067
rect 15642 11064 15654 11067
rect 15746 11064 15752 11076
rect 15642 11036 15752 11064
rect 15642 11033 15654 11036
rect 15596 11027 15654 11033
rect 15746 11024 15752 11036
rect 15804 11024 15810 11076
rect 19610 11024 19616 11076
rect 19668 11064 19674 11076
rect 19812 11064 19840 11095
rect 22462 11092 22468 11104
rect 22520 11092 22526 11144
rect 22557 11135 22615 11141
rect 22557 11101 22569 11135
rect 22603 11132 22615 11135
rect 23290 11132 23296 11144
rect 22603 11104 23296 11132
rect 22603 11101 22615 11104
rect 22557 11095 22615 11101
rect 23290 11092 23296 11104
rect 23348 11092 23354 11144
rect 23382 11092 23388 11144
rect 23440 11132 23446 11144
rect 26142 11132 26148 11144
rect 23440 11104 26148 11132
rect 23440 11092 23446 11104
rect 26142 11092 26148 11104
rect 26200 11092 26206 11144
rect 27080 11141 27108 11172
rect 27614 11160 27620 11172
rect 27672 11160 27678 11212
rect 27798 11160 27804 11212
rect 27856 11200 27862 11212
rect 28074 11200 28080 11212
rect 27856 11172 28080 11200
rect 27856 11160 27862 11172
rect 27065 11135 27123 11141
rect 27065 11101 27077 11135
rect 27111 11101 27123 11135
rect 27065 11095 27123 11101
rect 27249 11135 27307 11141
rect 27249 11101 27261 11135
rect 27295 11132 27307 11135
rect 27430 11132 27436 11144
rect 27295 11104 27436 11132
rect 27295 11101 27307 11104
rect 27249 11095 27307 11101
rect 27430 11092 27436 11104
rect 27488 11132 27494 11144
rect 27706 11132 27712 11144
rect 27488 11104 27712 11132
rect 27488 11092 27494 11104
rect 27706 11092 27712 11104
rect 27764 11092 27770 11144
rect 27908 11141 27936 11172
rect 28074 11160 28080 11172
rect 28132 11160 28138 11212
rect 28537 11203 28595 11209
rect 28537 11169 28549 11203
rect 28583 11200 28595 11203
rect 28626 11200 28632 11212
rect 28583 11172 28632 11200
rect 28583 11169 28595 11172
rect 28537 11163 28595 11169
rect 28626 11160 28632 11172
rect 28684 11160 28690 11212
rect 30653 11203 30711 11209
rect 30653 11200 30665 11203
rect 29564 11172 30665 11200
rect 29564 11144 29592 11172
rect 30653 11169 30665 11172
rect 30699 11200 30711 11203
rect 30742 11200 30748 11212
rect 30699 11172 30748 11200
rect 30699 11169 30711 11172
rect 30653 11163 30711 11169
rect 30742 11160 30748 11172
rect 30800 11160 30806 11212
rect 27893 11135 27951 11141
rect 27893 11101 27905 11135
rect 27939 11101 27951 11135
rect 27893 11095 27951 11101
rect 27982 11092 27988 11144
rect 28040 11132 28046 11144
rect 28721 11135 28779 11141
rect 28721 11132 28733 11135
rect 28040 11104 28733 11132
rect 28040 11092 28046 11104
rect 28721 11101 28733 11104
rect 28767 11101 28779 11135
rect 28721 11095 28779 11101
rect 29546 11092 29552 11144
rect 29604 11092 29610 11144
rect 29638 11092 29644 11144
rect 29696 11132 29702 11144
rect 29825 11135 29883 11141
rect 29825 11132 29837 11135
rect 29696 11104 29837 11132
rect 29696 11092 29702 11104
rect 29825 11101 29837 11104
rect 29871 11132 29883 11135
rect 30190 11132 30196 11144
rect 29871 11104 30196 11132
rect 29871 11101 29883 11104
rect 29825 11095 29883 11101
rect 30190 11092 30196 11104
rect 30248 11092 30254 11144
rect 34146 11092 34152 11144
rect 34204 11092 34210 11144
rect 34422 11092 34428 11144
rect 34480 11092 34486 11144
rect 19668 11036 19840 11064
rect 19668 11024 19674 11036
rect 22094 11024 22100 11076
rect 22152 11024 22158 11076
rect 22646 11024 22652 11076
rect 22704 11064 22710 11076
rect 23934 11064 23940 11076
rect 22704 11036 23940 11064
rect 22704 11024 22710 11036
rect 23934 11024 23940 11036
rect 23992 11024 23998 11076
rect 24664 11067 24722 11073
rect 24664 11033 24676 11067
rect 24710 11064 24722 11067
rect 24946 11064 24952 11076
rect 24710 11036 24952 11064
rect 24710 11033 24722 11036
rect 24664 11027 24722 11033
rect 24946 11024 24952 11036
rect 25004 11024 25010 11076
rect 27154 11064 27160 11076
rect 25424 11036 26004 11064
rect 1581 10999 1639 11005
rect 1581 10965 1593 10999
rect 1627 10965 1639 10999
rect 1581 10959 1639 10965
rect 4338 10956 4344 11008
rect 4396 10996 4402 11008
rect 5166 10996 5172 11008
rect 4396 10968 5172 10996
rect 4396 10956 4402 10968
rect 5166 10956 5172 10968
rect 5224 10996 5230 11008
rect 5442 10996 5448 11008
rect 5224 10968 5448 10996
rect 5224 10956 5230 10968
rect 5442 10956 5448 10968
rect 5500 10956 5506 11008
rect 8662 10956 8668 11008
rect 8720 10996 8726 11008
rect 13998 10996 14004 11008
rect 8720 10968 14004 10996
rect 8720 10956 8726 10968
rect 13998 10956 14004 10968
rect 14056 10956 14062 11008
rect 14826 10956 14832 11008
rect 14884 10996 14890 11008
rect 17770 10996 17776 11008
rect 14884 10968 17776 10996
rect 14884 10956 14890 10968
rect 17770 10956 17776 10968
rect 17828 10956 17834 11008
rect 19981 10999 20039 11005
rect 19981 10965 19993 10999
rect 20027 10996 20039 10999
rect 20622 10996 20628 11008
rect 20027 10968 20628 10996
rect 20027 10965 20039 10968
rect 19981 10959 20039 10965
rect 20622 10956 20628 10968
rect 20680 10956 20686 11008
rect 22370 10956 22376 11008
rect 22428 10996 22434 11008
rect 25424 10996 25452 11036
rect 22428 10968 25452 10996
rect 22428 10956 22434 10968
rect 25498 10956 25504 11008
rect 25556 10996 25562 11008
rect 25869 10999 25927 11005
rect 25869 10996 25881 10999
rect 25556 10968 25881 10996
rect 25556 10956 25562 10968
rect 25869 10965 25881 10968
rect 25915 10965 25927 10999
rect 25976 10996 26004 11036
rect 26896 11036 27160 11064
rect 26896 10996 26924 11036
rect 27154 11024 27160 11036
rect 27212 11024 27218 11076
rect 27522 11024 27528 11076
rect 27580 11024 27586 11076
rect 27614 11024 27620 11076
rect 27672 11024 27678 11076
rect 28629 11067 28687 11073
rect 28629 11064 28641 11067
rect 27724 11036 28641 11064
rect 25976 10968 26924 10996
rect 25869 10959 25927 10965
rect 26970 10956 26976 11008
rect 27028 10956 27034 11008
rect 27540 10996 27568 11024
rect 27724 10996 27752 11036
rect 28629 11033 28641 11036
rect 28675 11033 28687 11067
rect 28629 11027 28687 11033
rect 34333 11067 34391 11073
rect 34333 11033 34345 11067
rect 34379 11064 34391 11067
rect 34514 11064 34520 11076
rect 34379 11036 34520 11064
rect 34379 11033 34391 11036
rect 34333 11027 34391 11033
rect 34514 11024 34520 11036
rect 34572 11064 34578 11076
rect 34974 11064 34980 11076
rect 34572 11036 34980 11064
rect 34572 11024 34578 11036
rect 34974 11024 34980 11036
rect 35032 11024 35038 11076
rect 27540 10968 27752 10996
rect 28074 10956 28080 11008
rect 28132 10996 28138 11008
rect 28258 10996 28264 11008
rect 28132 10968 28264 10996
rect 28132 10956 28138 10968
rect 28258 10956 28264 10968
rect 28316 10956 28322 11008
rect 33502 10956 33508 11008
rect 33560 10996 33566 11008
rect 33965 10999 34023 11005
rect 33965 10996 33977 10999
rect 33560 10968 33977 10996
rect 33560 10956 33566 10968
rect 33965 10965 33977 10968
rect 34011 10965 34023 10999
rect 33965 10959 34023 10965
rect 1104 10906 35328 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35328 10906
rect 1104 10832 35328 10854
rect 3329 10795 3387 10801
rect 3329 10761 3341 10795
rect 3375 10761 3387 10795
rect 3329 10755 3387 10761
rect 2992 10727 3050 10733
rect 2992 10693 3004 10727
rect 3038 10724 3050 10727
rect 3344 10724 3372 10755
rect 3602 10752 3608 10804
rect 3660 10792 3666 10804
rect 3789 10795 3847 10801
rect 3789 10792 3801 10795
rect 3660 10764 3801 10792
rect 3660 10752 3666 10764
rect 3789 10761 3801 10764
rect 3835 10792 3847 10795
rect 4246 10792 4252 10804
rect 3835 10764 4252 10792
rect 3835 10761 3847 10764
rect 3789 10755 3847 10761
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 4709 10795 4767 10801
rect 4709 10761 4721 10795
rect 4755 10761 4767 10795
rect 4709 10755 4767 10761
rect 4433 10727 4491 10733
rect 4433 10724 4445 10727
rect 3038 10696 3372 10724
rect 3712 10696 4445 10724
rect 3038 10693 3050 10696
rect 2992 10687 3050 10693
rect 3234 10616 3240 10668
rect 3292 10616 3298 10668
rect 3712 10665 3740 10696
rect 4433 10693 4445 10696
rect 4479 10693 4491 10727
rect 4433 10687 4491 10693
rect 3697 10659 3755 10665
rect 3697 10625 3709 10659
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 1857 10455 1915 10461
rect 1857 10421 1869 10455
rect 1903 10452 1915 10455
rect 3712 10452 3740 10619
rect 4154 10616 4160 10668
rect 4212 10616 4218 10668
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 4525 10659 4583 10665
rect 4387 10628 4476 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 3973 10591 4031 10597
rect 3973 10557 3985 10591
rect 4019 10588 4031 10591
rect 4246 10588 4252 10600
rect 4019 10560 4252 10588
rect 4019 10557 4031 10560
rect 3973 10551 4031 10557
rect 4246 10548 4252 10560
rect 4304 10548 4310 10600
rect 1903 10424 3740 10452
rect 4448 10452 4476 10628
rect 4525 10625 4537 10659
rect 4571 10625 4583 10659
rect 4724 10656 4752 10755
rect 5074 10752 5080 10804
rect 5132 10792 5138 10804
rect 5132 10764 5396 10792
rect 5132 10752 5138 10764
rect 5258 10684 5264 10736
rect 5316 10684 5322 10736
rect 5368 10724 5396 10764
rect 5718 10752 5724 10804
rect 5776 10792 5782 10804
rect 8754 10792 8760 10804
rect 5776 10764 8760 10792
rect 5776 10752 5782 10764
rect 8754 10752 8760 10764
rect 8812 10752 8818 10804
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 10229 10795 10287 10801
rect 10229 10792 10241 10795
rect 10100 10764 10241 10792
rect 10100 10752 10106 10764
rect 10229 10761 10241 10764
rect 10275 10761 10287 10795
rect 10229 10755 10287 10761
rect 10410 10752 10416 10804
rect 10468 10792 10474 10804
rect 10873 10795 10931 10801
rect 10873 10792 10885 10795
rect 10468 10764 10885 10792
rect 10468 10752 10474 10764
rect 10873 10761 10885 10764
rect 10919 10761 10931 10795
rect 10873 10755 10931 10761
rect 11146 10752 11152 10804
rect 11204 10752 11210 10804
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 13817 10795 13875 10801
rect 13817 10792 13829 10795
rect 12860 10764 13829 10792
rect 12860 10752 12866 10764
rect 13817 10761 13829 10764
rect 13863 10792 13875 10795
rect 14001 10795 14059 10801
rect 14001 10792 14013 10795
rect 13863 10764 14013 10792
rect 13863 10761 13875 10764
rect 13817 10755 13875 10761
rect 14001 10761 14013 10764
rect 14047 10792 14059 10795
rect 14826 10792 14832 10804
rect 14047 10764 14832 10792
rect 14047 10761 14059 10764
rect 14001 10755 14059 10761
rect 14826 10752 14832 10764
rect 14884 10752 14890 10804
rect 15746 10752 15752 10804
rect 15804 10752 15810 10804
rect 16114 10752 16120 10804
rect 16172 10752 16178 10804
rect 18785 10795 18843 10801
rect 18785 10761 18797 10795
rect 18831 10792 18843 10795
rect 20625 10795 20683 10801
rect 20625 10792 20637 10795
rect 18831 10764 20637 10792
rect 18831 10761 18843 10764
rect 18785 10755 18843 10761
rect 20625 10761 20637 10764
rect 20671 10761 20683 10795
rect 22465 10795 22523 10801
rect 22465 10792 22477 10795
rect 20625 10755 20683 10761
rect 21330 10764 22477 10792
rect 12434 10724 12440 10736
rect 5368 10696 12440 10724
rect 12434 10684 12440 10696
rect 12492 10684 12498 10736
rect 14645 10727 14703 10733
rect 14645 10693 14657 10727
rect 14691 10724 14703 10727
rect 14734 10724 14740 10736
rect 14691 10696 14740 10724
rect 14691 10693 14703 10696
rect 14645 10687 14703 10693
rect 14734 10684 14740 10696
rect 14792 10684 14798 10736
rect 15470 10684 15476 10736
rect 15528 10684 15534 10736
rect 17126 10684 17132 10736
rect 17184 10684 17190 10736
rect 19426 10684 19432 10736
rect 19484 10724 19490 10736
rect 19484 10696 20208 10724
rect 19484 10684 19490 10696
rect 4893 10659 4951 10665
rect 4893 10656 4905 10659
rect 4724 10628 4905 10656
rect 4525 10619 4583 10625
rect 4893 10625 4905 10628
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 4986 10659 5044 10665
rect 4986 10625 4998 10659
rect 5032 10625 5044 10659
rect 4986 10619 5044 10625
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10625 5227 10659
rect 5169 10619 5227 10625
rect 5399 10659 5457 10665
rect 5399 10625 5411 10659
rect 5445 10656 5457 10659
rect 5445 10628 5856 10656
rect 5445 10625 5457 10628
rect 5399 10619 5457 10625
rect 4540 10520 4568 10619
rect 4614 10548 4620 10600
rect 4672 10588 4678 10600
rect 5000 10588 5028 10619
rect 4672 10560 5028 10588
rect 5184 10588 5212 10619
rect 5718 10588 5724 10600
rect 5184 10560 5724 10588
rect 4672 10548 4678 10560
rect 5718 10548 5724 10560
rect 5776 10548 5782 10600
rect 5828 10588 5856 10628
rect 5902 10616 5908 10668
rect 5960 10656 5966 10668
rect 12621 10659 12679 10665
rect 12621 10656 12633 10659
rect 5960 10628 12633 10656
rect 5960 10616 5966 10628
rect 12621 10625 12633 10628
rect 12667 10625 12679 10659
rect 12621 10619 12679 10625
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10656 14243 10659
rect 16758 10656 16764 10668
rect 14231 10628 14504 10656
rect 14231 10625 14243 10628
rect 14185 10619 14243 10625
rect 5828 10560 5948 10588
rect 4798 10520 4804 10532
rect 4540 10492 4804 10520
rect 4798 10480 4804 10492
rect 4856 10480 4862 10532
rect 4890 10452 4896 10464
rect 4448 10424 4896 10452
rect 1903 10421 1915 10424
rect 1857 10415 1915 10421
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 5534 10412 5540 10464
rect 5592 10412 5598 10464
rect 5920 10461 5948 10560
rect 10042 10548 10048 10600
rect 10100 10588 10106 10600
rect 12250 10588 12256 10600
rect 10100 10560 12256 10588
rect 10100 10548 10106 10560
rect 12250 10548 12256 10560
rect 12308 10588 12314 10600
rect 12897 10591 12955 10597
rect 12897 10588 12909 10591
rect 12308 10560 12909 10588
rect 12308 10548 12314 10560
rect 12897 10557 12909 10560
rect 12943 10557 12955 10591
rect 12897 10551 12955 10557
rect 14476 10529 14504 10628
rect 16408 10628 16764 10656
rect 14550 10548 14556 10600
rect 14608 10588 14614 10600
rect 16408 10597 16436 10628
rect 16758 10616 16764 10628
rect 16816 10656 16822 10668
rect 16942 10656 16948 10668
rect 16816 10628 16948 10656
rect 16816 10616 16822 10628
rect 16942 10616 16948 10628
rect 17000 10616 17006 10668
rect 17034 10616 17040 10668
rect 17092 10616 17098 10668
rect 17773 10659 17831 10665
rect 17773 10625 17785 10659
rect 17819 10656 17831 10659
rect 18141 10659 18199 10665
rect 18141 10656 18153 10659
rect 17819 10628 18153 10656
rect 17819 10625 17831 10628
rect 17773 10619 17831 10625
rect 18141 10625 18153 10628
rect 18187 10656 18199 10659
rect 18322 10656 18328 10668
rect 18187 10628 18328 10656
rect 18187 10625 18199 10628
rect 18141 10619 18199 10625
rect 18322 10616 18328 10628
rect 18380 10616 18386 10668
rect 20180 10665 20208 10696
rect 19909 10659 19967 10665
rect 19909 10625 19921 10659
rect 19955 10656 19967 10659
rect 20165 10659 20223 10665
rect 19955 10628 20116 10656
rect 19955 10625 19967 10628
rect 19909 10619 19967 10625
rect 16209 10591 16267 10597
rect 16209 10588 16221 10591
rect 14608 10560 16221 10588
rect 14608 10548 14614 10560
rect 16209 10557 16221 10560
rect 16255 10557 16267 10591
rect 16209 10551 16267 10557
rect 16393 10591 16451 10597
rect 16393 10557 16405 10591
rect 16439 10557 16451 10591
rect 16393 10551 16451 10557
rect 16850 10548 16856 10600
rect 16908 10588 16914 10600
rect 17221 10591 17279 10597
rect 17221 10588 17233 10591
rect 16908 10560 17233 10588
rect 16908 10548 16914 10560
rect 17221 10557 17233 10560
rect 17267 10588 17279 10591
rect 17865 10591 17923 10597
rect 17865 10588 17877 10591
rect 17267 10560 17877 10588
rect 17267 10557 17279 10560
rect 17221 10551 17279 10557
rect 17604 10529 17632 10560
rect 17865 10557 17877 10560
rect 17911 10588 17923 10591
rect 18233 10591 18291 10597
rect 18233 10588 18245 10591
rect 17911 10560 18245 10588
rect 17911 10557 17923 10560
rect 17865 10551 17923 10557
rect 18233 10557 18245 10560
rect 18279 10557 18291 10591
rect 20088 10588 20116 10628
rect 20165 10625 20177 10659
rect 20211 10656 20223 10659
rect 20346 10656 20352 10668
rect 20211 10628 20352 10656
rect 20211 10625 20223 10628
rect 20165 10619 20223 10625
rect 20346 10616 20352 10628
rect 20404 10616 20410 10668
rect 20640 10656 20668 10755
rect 21330 10724 21358 10764
rect 22465 10761 22477 10764
rect 22511 10792 22523 10795
rect 23382 10792 23388 10804
rect 22511 10764 23388 10792
rect 22511 10761 22523 10764
rect 22465 10755 22523 10761
rect 23382 10752 23388 10764
rect 23440 10752 23446 10804
rect 24946 10752 24952 10804
rect 25004 10752 25010 10804
rect 25409 10795 25467 10801
rect 25409 10761 25421 10795
rect 25455 10792 25467 10795
rect 26050 10792 26056 10804
rect 25455 10764 26056 10792
rect 25455 10761 25467 10764
rect 25409 10755 25467 10761
rect 26050 10752 26056 10764
rect 26108 10752 26114 10804
rect 26970 10752 26976 10804
rect 27028 10752 27034 10804
rect 28994 10792 29000 10804
rect 27356 10764 29000 10792
rect 21284 10696 21358 10724
rect 21453 10727 21511 10733
rect 21284 10665 21312 10696
rect 21453 10693 21465 10727
rect 21499 10724 21511 10727
rect 23842 10724 23848 10736
rect 21499 10696 23848 10724
rect 21499 10693 21511 10696
rect 21453 10687 21511 10693
rect 23842 10684 23848 10696
rect 23900 10684 23906 10736
rect 23934 10684 23940 10736
rect 23992 10724 23998 10736
rect 25317 10727 25375 10733
rect 25317 10724 25329 10727
rect 23992 10696 25329 10724
rect 23992 10684 23998 10696
rect 25317 10693 25329 10696
rect 25363 10693 25375 10727
rect 25317 10687 25375 10693
rect 21269 10659 21327 10665
rect 20640 10628 21220 10656
rect 20088 10560 20300 10588
rect 18233 10551 18291 10557
rect 20272 10529 20300 10560
rect 20622 10548 20628 10600
rect 20680 10588 20686 10600
rect 20717 10591 20775 10597
rect 20717 10588 20729 10591
rect 20680 10560 20729 10588
rect 20680 10548 20686 10560
rect 20717 10557 20729 10560
rect 20763 10557 20775 10591
rect 20717 10551 20775 10557
rect 20901 10591 20959 10597
rect 20901 10557 20913 10591
rect 20947 10557 20959 10591
rect 21192 10588 21220 10628
rect 21269 10625 21281 10659
rect 21315 10625 21327 10659
rect 21269 10619 21327 10625
rect 21358 10616 21364 10668
rect 21416 10616 21422 10668
rect 21637 10659 21695 10665
rect 21637 10625 21649 10659
rect 21683 10625 21695 10659
rect 21637 10619 21695 10625
rect 21652 10588 21680 10619
rect 21726 10616 21732 10668
rect 21784 10656 21790 10668
rect 21821 10659 21879 10665
rect 21821 10656 21833 10659
rect 21784 10628 21833 10656
rect 21784 10616 21790 10628
rect 21821 10625 21833 10628
rect 21867 10656 21879 10659
rect 22189 10659 22247 10665
rect 22189 10656 22201 10659
rect 21867 10628 22201 10656
rect 21867 10625 21879 10628
rect 21821 10619 21879 10625
rect 22189 10625 22201 10628
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 22649 10659 22707 10665
rect 22649 10625 22661 10659
rect 22695 10656 22707 10659
rect 25590 10656 25596 10668
rect 22695 10628 25596 10656
rect 22695 10625 22707 10628
rect 22649 10619 22707 10625
rect 21192 10560 21680 10588
rect 20901 10551 20959 10557
rect 14461 10523 14519 10529
rect 14461 10489 14473 10523
rect 14507 10520 14519 10523
rect 17589 10523 17647 10529
rect 14507 10492 16896 10520
rect 14507 10489 14519 10492
rect 14461 10483 14519 10489
rect 5905 10455 5963 10461
rect 5905 10421 5917 10455
rect 5951 10452 5963 10455
rect 10042 10452 10048 10464
rect 5951 10424 10048 10452
rect 5951 10421 5963 10424
rect 5905 10415 5963 10421
rect 10042 10412 10048 10424
rect 10100 10452 10106 10464
rect 10778 10452 10784 10464
rect 10100 10424 10784 10452
rect 10100 10412 10106 10424
rect 10778 10412 10784 10424
rect 10836 10452 10842 10464
rect 11241 10455 11299 10461
rect 11241 10452 11253 10455
rect 10836 10424 11253 10452
rect 10836 10412 10842 10424
rect 11241 10421 11253 10424
rect 11287 10421 11299 10455
rect 11241 10415 11299 10421
rect 12158 10412 12164 10464
rect 12216 10452 12222 10464
rect 12805 10455 12863 10461
rect 12805 10452 12817 10455
rect 12216 10424 12817 10452
rect 12216 10412 12222 10424
rect 12805 10421 12817 10424
rect 12851 10452 12863 10455
rect 13814 10452 13820 10464
rect 12851 10424 13820 10452
rect 12851 10421 12863 10424
rect 12805 10415 12863 10421
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 16022 10412 16028 10464
rect 16080 10452 16086 10464
rect 16669 10455 16727 10461
rect 16669 10452 16681 10455
rect 16080 10424 16681 10452
rect 16080 10412 16086 10424
rect 16669 10421 16681 10424
rect 16715 10421 16727 10455
rect 16868 10452 16896 10492
rect 17589 10489 17601 10523
rect 17635 10489 17647 10523
rect 17589 10483 17647 10489
rect 20257 10523 20315 10529
rect 20257 10489 20269 10523
rect 20303 10489 20315 10523
rect 20916 10520 20944 10551
rect 21910 10548 21916 10600
rect 21968 10588 21974 10600
rect 22664 10588 22692 10619
rect 25590 10616 25596 10628
rect 25648 10616 25654 10668
rect 21968 10560 22692 10588
rect 21968 10548 21974 10560
rect 25498 10548 25504 10600
rect 25556 10588 25562 10600
rect 25777 10591 25835 10597
rect 25777 10588 25789 10591
rect 25556 10560 25789 10588
rect 25556 10548 25562 10560
rect 25777 10557 25789 10560
rect 25823 10557 25835 10591
rect 25777 10551 25835 10557
rect 27356 10520 27384 10764
rect 28994 10752 29000 10764
rect 29052 10792 29058 10804
rect 29638 10792 29644 10804
rect 29052 10764 29644 10792
rect 29052 10752 29058 10764
rect 29638 10752 29644 10764
rect 29696 10752 29702 10804
rect 29917 10795 29975 10801
rect 29917 10761 29929 10795
rect 29963 10761 29975 10795
rect 29917 10755 29975 10761
rect 29086 10724 29092 10736
rect 28368 10696 29092 10724
rect 27522 10616 27528 10668
rect 27580 10656 27586 10668
rect 28368 10665 28396 10696
rect 29086 10684 29092 10696
rect 29144 10684 29150 10736
rect 29558 10727 29616 10733
rect 29558 10693 29570 10727
rect 29604 10724 29616 10727
rect 29932 10724 29960 10755
rect 30282 10752 30288 10804
rect 30340 10792 30346 10804
rect 30377 10795 30435 10801
rect 30377 10792 30389 10795
rect 30340 10764 30389 10792
rect 30340 10752 30346 10764
rect 30377 10761 30389 10764
rect 30423 10761 30435 10795
rect 30377 10755 30435 10761
rect 34974 10752 34980 10804
rect 35032 10752 35038 10804
rect 29604 10696 29960 10724
rect 29604 10693 29616 10696
rect 29558 10687 29616 10693
rect 30190 10684 30196 10736
rect 30248 10724 30254 10736
rect 30248 10696 30512 10724
rect 30248 10684 30254 10696
rect 28086 10659 28144 10665
rect 28086 10656 28098 10659
rect 27580 10628 28098 10656
rect 27580 10616 27586 10628
rect 28086 10625 28098 10628
rect 28132 10625 28144 10659
rect 28086 10619 28144 10625
rect 28353 10659 28411 10665
rect 28353 10625 28365 10659
rect 28399 10625 28411 10659
rect 28994 10656 29000 10668
rect 28353 10619 28411 10625
rect 28828 10628 29000 10656
rect 28828 10520 28856 10628
rect 28994 10616 29000 10628
rect 29052 10656 29058 10668
rect 29270 10656 29276 10668
rect 29052 10628 29276 10656
rect 29052 10616 29058 10628
rect 29270 10616 29276 10628
rect 29328 10616 29334 10668
rect 30285 10659 30343 10665
rect 30285 10625 30297 10659
rect 30331 10625 30343 10659
rect 30285 10619 30343 10625
rect 29822 10548 29828 10600
rect 29880 10548 29886 10600
rect 20916 10492 27384 10520
rect 28368 10492 28856 10520
rect 20257 10483 20315 10489
rect 20806 10452 20812 10464
rect 16868 10424 20812 10452
rect 16669 10415 16727 10421
rect 20806 10412 20812 10424
rect 20864 10412 20870 10464
rect 21082 10412 21088 10464
rect 21140 10412 21146 10464
rect 21818 10412 21824 10464
rect 21876 10452 21882 10464
rect 22005 10455 22063 10461
rect 22005 10452 22017 10455
rect 21876 10424 22017 10452
rect 21876 10412 21882 10424
rect 22005 10421 22017 10424
rect 22051 10421 22063 10455
rect 22005 10415 22063 10421
rect 23842 10412 23848 10464
rect 23900 10452 23906 10464
rect 28368 10452 28396 10492
rect 23900 10424 28396 10452
rect 28445 10455 28503 10461
rect 23900 10412 23906 10424
rect 28445 10421 28457 10455
rect 28491 10452 28503 10455
rect 29178 10452 29184 10464
rect 28491 10424 29184 10452
rect 28491 10421 28503 10424
rect 28445 10415 28503 10421
rect 29178 10412 29184 10424
rect 29236 10452 29242 10464
rect 30300 10452 30328 10619
rect 30484 10597 30512 10696
rect 33502 10684 33508 10736
rect 33560 10684 33566 10736
rect 34514 10684 34520 10736
rect 34572 10684 34578 10736
rect 30469 10591 30527 10597
rect 30469 10557 30481 10591
rect 30515 10557 30527 10591
rect 30469 10551 30527 10557
rect 32766 10548 32772 10600
rect 32824 10588 32830 10600
rect 33229 10591 33287 10597
rect 33229 10588 33241 10591
rect 32824 10560 33241 10588
rect 32824 10548 32830 10560
rect 33229 10557 33241 10560
rect 33275 10557 33287 10591
rect 33229 10551 33287 10557
rect 29236 10424 30328 10452
rect 29236 10412 29242 10424
rect 1104 10362 35328 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 35328 10362
rect 1104 10288 35328 10310
rect 3237 10251 3295 10257
rect 3237 10217 3249 10251
rect 3283 10248 3295 10251
rect 3602 10248 3608 10260
rect 3283 10220 3608 10248
rect 3283 10217 3295 10220
rect 3237 10211 3295 10217
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 4890 10208 4896 10260
rect 4948 10248 4954 10260
rect 5626 10248 5632 10260
rect 4948 10220 5632 10248
rect 4948 10208 4954 10220
rect 5626 10208 5632 10220
rect 5684 10248 5690 10260
rect 6733 10251 6791 10257
rect 6733 10248 6745 10251
rect 5684 10220 6745 10248
rect 5684 10208 5690 10220
rect 6733 10217 6745 10220
rect 6779 10217 6791 10251
rect 6733 10211 6791 10217
rect 8662 10208 8668 10260
rect 8720 10208 8726 10260
rect 8754 10208 8760 10260
rect 8812 10248 8818 10260
rect 9861 10251 9919 10257
rect 9861 10248 9873 10251
rect 8812 10220 9873 10248
rect 8812 10208 8818 10220
rect 9861 10217 9873 10220
rect 9907 10248 9919 10251
rect 10410 10248 10416 10260
rect 9907 10220 10416 10248
rect 9907 10217 9919 10220
rect 9861 10211 9919 10217
rect 10410 10208 10416 10220
rect 10468 10248 10474 10260
rect 11514 10248 11520 10260
rect 10468 10220 11520 10248
rect 10468 10208 10474 10220
rect 11514 10208 11520 10220
rect 11572 10208 11578 10260
rect 11609 10251 11667 10257
rect 11609 10217 11621 10251
rect 11655 10248 11667 10251
rect 11790 10248 11796 10260
rect 11655 10220 11796 10248
rect 11655 10217 11667 10220
rect 11609 10211 11667 10217
rect 3620 9976 3648 10208
rect 4706 10180 4712 10192
rect 4448 10152 4712 10180
rect 4338 10072 4344 10124
rect 4396 10112 4402 10124
rect 4448 10121 4476 10152
rect 4706 10140 4712 10152
rect 4764 10140 4770 10192
rect 5261 10183 5319 10189
rect 5261 10149 5273 10183
rect 5307 10180 5319 10183
rect 8297 10183 8355 10189
rect 5307 10152 6592 10180
rect 5307 10149 5319 10152
rect 5261 10143 5319 10149
rect 4433 10115 4491 10121
rect 4433 10112 4445 10115
rect 4396 10084 4445 10112
rect 4396 10072 4402 10084
rect 4433 10081 4445 10084
rect 4479 10081 4491 10115
rect 4433 10075 4491 10081
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4246 10044 4252 10056
rect 4203 10016 4252 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 4246 10004 4252 10016
rect 4304 10004 4310 10056
rect 4706 10004 4712 10056
rect 4764 10044 4770 10056
rect 5074 10044 5080 10056
rect 4764 10016 5080 10044
rect 4764 10004 4770 10016
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 5368 10053 5396 10152
rect 6564 10112 6592 10152
rect 8297 10149 8309 10183
rect 8343 10180 8355 10183
rect 9950 10180 9956 10192
rect 8343 10152 9956 10180
rect 8343 10149 8355 10152
rect 8297 10143 8355 10149
rect 9950 10140 9956 10152
rect 10008 10140 10014 10192
rect 9766 10112 9772 10124
rect 5460 10084 6500 10112
rect 6564 10084 9772 10112
rect 5353 10047 5411 10053
rect 5353 10013 5365 10047
rect 5399 10013 5411 10047
rect 5353 10007 5411 10013
rect 3620 9948 4292 9976
rect 3786 9868 3792 9920
rect 3844 9868 3850 9920
rect 4264 9917 4292 9948
rect 4798 9936 4804 9988
rect 4856 9976 4862 9988
rect 5460 9976 5488 10084
rect 5718 10004 5724 10056
rect 5776 10044 5782 10056
rect 6472 10053 6500 10084
rect 7834 10053 7840 10056
rect 6089 10047 6147 10053
rect 6089 10044 6101 10047
rect 5776 10016 6101 10044
rect 5776 10004 5782 10016
rect 6089 10013 6101 10016
rect 6135 10013 6147 10047
rect 6089 10007 6147 10013
rect 6457 10047 6515 10053
rect 6457 10013 6469 10047
rect 6503 10013 6515 10047
rect 7653 10047 7711 10053
rect 7653 10044 7665 10047
rect 6457 10007 6515 10013
rect 6656 10016 7665 10044
rect 4856 9948 5488 9976
rect 4856 9936 4862 9948
rect 5626 9936 5632 9988
rect 5684 9976 5690 9988
rect 6273 9979 6331 9985
rect 6273 9976 6285 9979
rect 5684 9948 6285 9976
rect 5684 9936 5690 9948
rect 6273 9945 6285 9948
rect 6319 9945 6331 9979
rect 6273 9939 6331 9945
rect 6362 9936 6368 9988
rect 6420 9936 6426 9988
rect 4249 9911 4307 9917
rect 4249 9877 4261 9911
rect 4295 9877 4307 9911
rect 4249 9871 4307 9877
rect 5537 9911 5595 9917
rect 5537 9877 5549 9911
rect 5583 9908 5595 9911
rect 5902 9908 5908 9920
rect 5583 9880 5908 9908
rect 5583 9877 5595 9880
rect 5537 9871 5595 9877
rect 5902 9868 5908 9880
rect 5960 9868 5966 9920
rect 6656 9917 6684 10016
rect 7653 10013 7665 10016
rect 7699 10013 7711 10047
rect 7653 10007 7711 10013
rect 7801 10047 7840 10053
rect 7801 10013 7813 10047
rect 7801 10007 7840 10013
rect 7834 10004 7840 10007
rect 7892 10004 7898 10056
rect 8159 10047 8217 10053
rect 8159 10013 8171 10047
rect 8205 10044 8217 10047
rect 8662 10044 8668 10056
rect 8205 10016 8668 10044
rect 8205 10013 8217 10016
rect 8159 10007 8217 10013
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 9324 10053 9352 10084
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 10870 10072 10876 10124
rect 10928 10112 10934 10124
rect 11333 10115 11391 10121
rect 11333 10112 11345 10115
rect 10928 10084 11345 10112
rect 10928 10072 10934 10084
rect 11333 10081 11345 10084
rect 11379 10081 11391 10115
rect 11333 10075 11391 10081
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10013 9367 10047
rect 9309 10007 9367 10013
rect 10042 10004 10048 10056
rect 10100 10044 10106 10056
rect 10224 10047 10282 10053
rect 10224 10044 10236 10047
rect 10100 10016 10236 10044
rect 10100 10004 10106 10016
rect 10224 10013 10236 10016
rect 10270 10013 10282 10047
rect 10224 10007 10282 10013
rect 10410 10004 10416 10056
rect 10468 10004 10474 10056
rect 10502 10004 10508 10056
rect 10560 10053 10566 10056
rect 10560 10047 10599 10053
rect 10587 10013 10599 10047
rect 10560 10007 10599 10013
rect 10560 10004 10566 10007
rect 10686 10004 10692 10056
rect 10744 10004 10750 10056
rect 11149 10047 11207 10053
rect 11149 10013 11161 10047
rect 11195 10044 11207 10047
rect 11624 10044 11652 10211
rect 11790 10208 11796 10220
rect 11848 10208 11854 10260
rect 13906 10208 13912 10260
rect 13964 10248 13970 10260
rect 14458 10248 14464 10260
rect 13964 10220 14464 10248
rect 13964 10208 13970 10220
rect 14458 10208 14464 10220
rect 14516 10208 14522 10260
rect 17034 10208 17040 10260
rect 17092 10248 17098 10260
rect 17129 10251 17187 10257
rect 17129 10248 17141 10251
rect 17092 10220 17141 10248
rect 17092 10208 17098 10220
rect 17129 10217 17141 10220
rect 17175 10217 17187 10251
rect 17129 10211 17187 10217
rect 12158 10072 12164 10124
rect 12216 10072 12222 10124
rect 12250 10072 12256 10124
rect 12308 10072 12314 10124
rect 12526 10072 12532 10124
rect 12584 10072 12590 10124
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 14550 10112 14556 10124
rect 13872 10084 14556 10112
rect 13872 10072 13878 10084
rect 14550 10072 14556 10084
rect 14608 10072 14614 10124
rect 14737 10115 14795 10121
rect 14737 10081 14749 10115
rect 14783 10112 14795 10115
rect 14826 10112 14832 10124
rect 14783 10084 14832 10112
rect 14783 10081 14795 10084
rect 14737 10075 14795 10081
rect 14826 10072 14832 10084
rect 14884 10072 14890 10124
rect 15470 10072 15476 10124
rect 15528 10112 15534 10124
rect 15749 10115 15807 10121
rect 15749 10112 15761 10115
rect 15528 10084 15761 10112
rect 15528 10072 15534 10084
rect 15749 10081 15761 10084
rect 15795 10081 15807 10115
rect 15749 10075 15807 10081
rect 11195 10016 11652 10044
rect 11195 10013 11207 10016
rect 11149 10007 11207 10013
rect 13630 10004 13636 10056
rect 13688 10044 13694 10056
rect 13688 10016 14412 10044
rect 13688 10004 13694 10016
rect 7929 9979 7987 9985
rect 7929 9945 7941 9979
rect 7975 9945 7987 9979
rect 7929 9939 7987 9945
rect 6641 9911 6699 9917
rect 6641 9877 6653 9911
rect 6687 9877 6699 9911
rect 7944 9908 7972 9939
rect 8018 9936 8024 9988
rect 8076 9936 8082 9988
rect 8481 9979 8539 9985
rect 8481 9945 8493 9979
rect 8527 9976 8539 9979
rect 9398 9976 9404 9988
rect 8527 9948 9404 9976
rect 8527 9945 8539 9948
rect 8481 9939 8539 9945
rect 8496 9908 8524 9939
rect 9398 9936 9404 9948
rect 9456 9936 9462 9988
rect 10134 9936 10140 9988
rect 10192 9976 10198 9988
rect 10301 9979 10359 9985
rect 10301 9976 10313 9979
rect 10192 9948 10313 9976
rect 10192 9936 10198 9948
rect 10301 9945 10313 9948
rect 10347 9945 10359 9979
rect 10301 9939 10359 9945
rect 12069 9979 12127 9985
rect 12069 9945 12081 9979
rect 12115 9976 12127 9979
rect 12796 9979 12854 9985
rect 12115 9948 12434 9976
rect 12115 9945 12127 9948
rect 12069 9939 12127 9945
rect 7944 9880 8524 9908
rect 9493 9911 9551 9917
rect 6641 9871 6699 9877
rect 9493 9877 9505 9911
rect 9539 9908 9551 9911
rect 9582 9908 9588 9920
rect 9539 9880 9588 9908
rect 9539 9877 9551 9880
rect 9493 9871 9551 9877
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 10042 9868 10048 9920
rect 10100 9868 10106 9920
rect 11698 9868 11704 9920
rect 11756 9868 11762 9920
rect 12406 9908 12434 9948
rect 12796 9945 12808 9979
rect 12842 9976 12854 9979
rect 14384 9976 14412 10016
rect 14458 10004 14464 10056
rect 14516 10004 14522 10056
rect 16022 10053 16028 10056
rect 16016 10044 16028 10053
rect 15983 10016 16028 10044
rect 16016 10007 16028 10016
rect 16022 10004 16028 10007
rect 16080 10004 16086 10056
rect 17144 10044 17172 10211
rect 17770 10208 17776 10260
rect 17828 10248 17834 10260
rect 17828 10220 22094 10248
rect 17828 10208 17834 10220
rect 17402 10140 17408 10192
rect 17460 10180 17466 10192
rect 17865 10183 17923 10189
rect 17865 10180 17877 10183
rect 17460 10152 17877 10180
rect 17460 10140 17466 10152
rect 17865 10149 17877 10152
rect 17911 10149 17923 10183
rect 17865 10143 17923 10149
rect 18414 10140 18420 10192
rect 18472 10180 18478 10192
rect 18785 10183 18843 10189
rect 18785 10180 18797 10183
rect 18472 10152 18797 10180
rect 18472 10140 18478 10152
rect 18785 10149 18797 10152
rect 18831 10180 18843 10183
rect 22066 10180 22094 10220
rect 22278 10208 22284 10260
rect 22336 10248 22342 10260
rect 22925 10251 22983 10257
rect 22925 10248 22937 10251
rect 22336 10220 22937 10248
rect 22336 10208 22342 10220
rect 22925 10217 22937 10220
rect 22971 10217 22983 10251
rect 22925 10211 22983 10217
rect 23477 10251 23535 10257
rect 23477 10217 23489 10251
rect 23523 10248 23535 10251
rect 23566 10248 23572 10260
rect 23523 10220 23572 10248
rect 23523 10217 23535 10220
rect 23477 10211 23535 10217
rect 23566 10208 23572 10220
rect 23624 10208 23630 10260
rect 24581 10251 24639 10257
rect 24581 10217 24593 10251
rect 24627 10248 24639 10251
rect 24627 10220 25912 10248
rect 24627 10217 24639 10220
rect 24581 10211 24639 10217
rect 25498 10180 25504 10192
rect 18831 10152 19334 10180
rect 22066 10152 25504 10180
rect 18831 10149 18843 10152
rect 18785 10143 18843 10149
rect 18877 10115 18935 10121
rect 18877 10112 18889 10115
rect 17328 10084 18889 10112
rect 17221 10047 17279 10053
rect 17221 10044 17233 10047
rect 17144 10016 17233 10044
rect 17221 10013 17233 10016
rect 17267 10013 17279 10047
rect 17221 10007 17279 10013
rect 17328 9976 17356 10084
rect 17402 10004 17408 10056
rect 17460 10004 17466 10056
rect 17604 10053 17632 10084
rect 18877 10081 18889 10084
rect 18923 10081 18935 10115
rect 18877 10075 18935 10081
rect 17589 10047 17647 10053
rect 17589 10013 17601 10047
rect 17635 10013 17647 10047
rect 17589 10007 17647 10013
rect 18414 10004 18420 10056
rect 18472 10004 18478 10056
rect 12842 9948 14136 9976
rect 14384 9948 17356 9976
rect 17493 9979 17551 9985
rect 12842 9945 12854 9948
rect 12796 9939 12854 9945
rect 13354 9908 13360 9920
rect 12406 9880 13360 9908
rect 13354 9868 13360 9880
rect 13412 9868 13418 9920
rect 14108 9917 14136 9948
rect 17493 9945 17505 9979
rect 17539 9976 17551 9979
rect 18782 9976 18788 9988
rect 17539 9948 18788 9976
rect 17539 9945 17551 9948
rect 17493 9939 17551 9945
rect 18782 9936 18788 9948
rect 18840 9936 18846 9988
rect 14093 9911 14151 9917
rect 14093 9877 14105 9911
rect 14139 9877 14151 9911
rect 14093 9871 14151 9877
rect 17310 9868 17316 9920
rect 17368 9908 17374 9920
rect 17773 9911 17831 9917
rect 17773 9908 17785 9911
rect 17368 9880 17785 9908
rect 17368 9868 17374 9880
rect 17773 9877 17785 9880
rect 17819 9877 17831 9911
rect 17773 9871 17831 9877
rect 18233 9911 18291 9917
rect 18233 9877 18245 9911
rect 18279 9908 18291 9911
rect 18322 9908 18328 9920
rect 18279 9880 18328 9908
rect 18279 9877 18291 9880
rect 18233 9871 18291 9877
rect 18322 9868 18328 9880
rect 18380 9908 18386 9920
rect 18509 9911 18567 9917
rect 18509 9908 18521 9911
rect 18380 9880 18521 9908
rect 18380 9868 18386 9880
rect 18509 9877 18521 9880
rect 18555 9877 18567 9911
rect 18892 9908 18920 10075
rect 19306 10044 19334 10152
rect 25498 10140 25504 10152
rect 25556 10140 25562 10192
rect 25884 10180 25912 10220
rect 26786 10208 26792 10260
rect 26844 10248 26850 10260
rect 27154 10248 27160 10260
rect 26844 10220 27160 10248
rect 26844 10208 26850 10220
rect 27154 10208 27160 10220
rect 27212 10208 27218 10260
rect 27433 10251 27491 10257
rect 27433 10217 27445 10251
rect 27479 10248 27491 10251
rect 27522 10248 27528 10260
rect 27479 10220 27528 10248
rect 27479 10217 27491 10220
rect 27433 10211 27491 10217
rect 27522 10208 27528 10220
rect 27580 10208 27586 10260
rect 27706 10208 27712 10260
rect 27764 10208 27770 10260
rect 27798 10208 27804 10260
rect 27856 10248 27862 10260
rect 27893 10251 27951 10257
rect 27893 10248 27905 10251
rect 27856 10220 27905 10248
rect 27856 10208 27862 10220
rect 27893 10217 27905 10220
rect 27939 10248 27951 10251
rect 28077 10251 28135 10257
rect 28077 10248 28089 10251
rect 27939 10220 28089 10248
rect 27939 10217 27951 10220
rect 27893 10211 27951 10217
rect 28077 10217 28089 10220
rect 28123 10217 28135 10251
rect 28077 10211 28135 10217
rect 28353 10251 28411 10257
rect 28353 10217 28365 10251
rect 28399 10248 28411 10251
rect 28626 10248 28632 10260
rect 28399 10220 28632 10248
rect 28399 10217 28411 10220
rect 28353 10211 28411 10217
rect 28626 10208 28632 10220
rect 28684 10208 28690 10260
rect 29086 10208 29092 10260
rect 29144 10248 29150 10260
rect 29822 10248 29828 10260
rect 29144 10220 29828 10248
rect 29144 10208 29150 10220
rect 29822 10208 29828 10220
rect 29880 10208 29886 10260
rect 28166 10180 28172 10192
rect 25884 10152 28172 10180
rect 28166 10140 28172 10152
rect 28224 10140 28230 10192
rect 20346 10072 20352 10124
rect 20404 10072 20410 10124
rect 22462 10072 22468 10124
rect 22520 10112 22526 10124
rect 23109 10115 23167 10121
rect 23109 10112 23121 10115
rect 22520 10084 23121 10112
rect 22520 10072 22526 10084
rect 23109 10081 23121 10084
rect 23155 10081 23167 10115
rect 23109 10075 23167 10081
rect 23216 10084 23520 10112
rect 19794 10044 19800 10056
rect 19306 10016 19800 10044
rect 19794 10004 19800 10016
rect 19852 10044 19858 10056
rect 22370 10044 22376 10056
rect 19852 10016 22376 10044
rect 19852 10004 19858 10016
rect 22370 10004 22376 10016
rect 22428 10004 22434 10056
rect 22554 10004 22560 10056
rect 22612 10044 22618 10056
rect 22741 10047 22799 10053
rect 22741 10044 22753 10047
rect 22612 10016 22753 10044
rect 22612 10004 22618 10016
rect 22741 10013 22753 10016
rect 22787 10013 22799 10047
rect 22741 10007 22799 10013
rect 22925 10047 22983 10053
rect 22925 10013 22937 10047
rect 22971 10013 22983 10047
rect 22925 10007 22983 10013
rect 20622 9985 20628 9988
rect 20616 9939 20628 9985
rect 20622 9936 20628 9939
rect 20680 9936 20686 9988
rect 21910 9976 21916 9988
rect 20732 9948 21916 9976
rect 20732 9908 20760 9948
rect 21910 9936 21916 9948
rect 21968 9936 21974 9988
rect 18892 9880 20760 9908
rect 18509 9871 18567 9877
rect 20990 9868 20996 9920
rect 21048 9908 21054 9920
rect 21358 9908 21364 9920
rect 21048 9880 21364 9908
rect 21048 9868 21054 9880
rect 21358 9868 21364 9880
rect 21416 9908 21422 9920
rect 21729 9911 21787 9917
rect 21729 9908 21741 9911
rect 21416 9880 21741 9908
rect 21416 9868 21422 9880
rect 21729 9877 21741 9880
rect 21775 9877 21787 9911
rect 22940 9908 22968 10007
rect 23014 10004 23020 10056
rect 23072 10004 23078 10056
rect 23216 10053 23244 10084
rect 23492 10056 23520 10084
rect 26786 10072 26792 10124
rect 26844 10072 26850 10124
rect 30101 10115 30159 10121
rect 30101 10112 30113 10115
rect 28828 10084 30113 10112
rect 28828 10056 28856 10084
rect 30101 10081 30113 10084
rect 30147 10081 30159 10115
rect 30101 10075 30159 10081
rect 23201 10047 23259 10053
rect 23201 10013 23213 10047
rect 23247 10013 23259 10047
rect 23201 10007 23259 10013
rect 23290 10004 23296 10056
rect 23348 10004 23354 10056
rect 23474 10004 23480 10056
rect 23532 10004 23538 10056
rect 23569 10047 23627 10053
rect 23569 10013 23581 10047
rect 23615 10013 23627 10047
rect 23569 10007 23627 10013
rect 23753 10047 23811 10053
rect 23753 10013 23765 10047
rect 23799 10013 23811 10047
rect 23753 10007 23811 10013
rect 23032 9976 23060 10004
rect 23584 9976 23612 10007
rect 23032 9948 23612 9976
rect 23768 9976 23796 10007
rect 24394 10004 24400 10056
rect 24452 10004 24458 10056
rect 24581 10047 24639 10053
rect 24581 10013 24593 10047
rect 24627 10044 24639 10047
rect 24762 10044 24768 10056
rect 24627 10016 24768 10044
rect 24627 10013 24639 10016
rect 24581 10007 24639 10013
rect 24596 9976 24624 10007
rect 24762 10004 24768 10016
rect 24820 10004 24826 10056
rect 26970 10004 26976 10056
rect 27028 10044 27034 10056
rect 27065 10047 27123 10053
rect 27065 10044 27077 10047
rect 27028 10016 27077 10044
rect 27028 10004 27034 10016
rect 27065 10013 27077 10016
rect 27111 10013 27123 10047
rect 27065 10007 27123 10013
rect 27154 10004 27160 10056
rect 27212 10044 27218 10056
rect 27617 10047 27675 10053
rect 27617 10044 27629 10047
rect 27212 10016 27629 10044
rect 27212 10004 27218 10016
rect 27617 10013 27629 10016
rect 27663 10044 27675 10047
rect 28074 10044 28080 10056
rect 27663 10016 28080 10044
rect 27663 10013 27675 10016
rect 27617 10007 27675 10013
rect 28074 10004 28080 10016
rect 28132 10004 28138 10056
rect 28810 10053 28816 10056
rect 28808 10044 28816 10053
rect 28771 10016 28816 10044
rect 28808 10007 28816 10016
rect 28810 10004 28816 10007
rect 28868 10004 28874 10056
rect 28994 10004 29000 10056
rect 29052 10004 29058 10056
rect 29178 10044 29184 10056
rect 29139 10016 29184 10044
rect 29178 10004 29184 10016
rect 29236 10004 29242 10056
rect 29270 10004 29276 10056
rect 29328 10004 29334 10056
rect 29638 10004 29644 10056
rect 29696 10004 29702 10056
rect 29822 10004 29828 10056
rect 29880 10044 29886 10056
rect 31021 10047 31079 10053
rect 31021 10044 31033 10047
rect 29880 10016 31033 10044
rect 29880 10004 29886 10016
rect 31021 10013 31033 10016
rect 31067 10044 31079 10047
rect 31067 10016 32076 10044
rect 31067 10013 31079 10016
rect 31021 10007 31079 10013
rect 27890 9976 27896 9988
rect 23768 9948 24624 9976
rect 25792 9948 27896 9976
rect 23198 9908 23204 9920
rect 22940 9880 23204 9908
rect 21729 9871 21787 9877
rect 23198 9868 23204 9880
rect 23256 9868 23262 9920
rect 23661 9911 23719 9917
rect 23661 9877 23673 9911
rect 23707 9908 23719 9911
rect 25792 9908 25820 9948
rect 27890 9936 27896 9948
rect 27948 9936 27954 9988
rect 28902 9936 28908 9988
rect 28960 9936 28966 9988
rect 29656 9976 29684 10004
rect 30285 9979 30343 9985
rect 30285 9976 30297 9979
rect 29656 9948 30297 9976
rect 30285 9945 30297 9948
rect 30331 9945 30343 9979
rect 30285 9939 30343 9945
rect 31202 9936 31208 9988
rect 31260 9936 31266 9988
rect 32048 9985 32076 10016
rect 32033 9979 32091 9985
rect 32033 9945 32045 9979
rect 32079 9976 32091 9979
rect 32766 9976 32772 9988
rect 32079 9948 32772 9976
rect 32079 9945 32091 9948
rect 32033 9939 32091 9945
rect 32766 9936 32772 9948
rect 32824 9936 32830 9988
rect 23707 9880 25820 9908
rect 26973 9911 27031 9917
rect 23707 9877 23719 9880
rect 23661 9871 23719 9877
rect 26973 9877 26985 9911
rect 27019 9908 27031 9911
rect 27246 9908 27252 9920
rect 27019 9880 27252 9908
rect 27019 9877 27031 9880
rect 26973 9871 27031 9877
rect 27246 9868 27252 9880
rect 27304 9868 27310 9920
rect 28258 9868 28264 9920
rect 28316 9908 28322 9920
rect 28445 9911 28503 9917
rect 28445 9908 28457 9911
rect 28316 9880 28457 9908
rect 28316 9868 28322 9880
rect 28445 9877 28457 9880
rect 28491 9877 28503 9911
rect 28445 9871 28503 9877
rect 28534 9868 28540 9920
rect 28592 9908 28598 9920
rect 28629 9911 28687 9917
rect 28629 9908 28641 9911
rect 28592 9880 28641 9908
rect 28592 9868 28598 9880
rect 28629 9877 28641 9880
rect 28675 9877 28687 9911
rect 28629 9871 28687 9877
rect 29730 9868 29736 9920
rect 29788 9908 29794 9920
rect 30466 9908 30472 9920
rect 29788 9880 30472 9908
rect 29788 9868 29794 9880
rect 30466 9868 30472 9880
rect 30524 9868 30530 9920
rect 1104 9818 35328 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35328 9818
rect 1104 9744 35328 9766
rect 4338 9664 4344 9716
rect 4396 9664 4402 9716
rect 5626 9664 5632 9716
rect 5684 9704 5690 9716
rect 5684 9676 6868 9704
rect 5684 9664 5690 9676
rect 3636 9639 3694 9645
rect 3636 9605 3648 9639
rect 3682 9636 3694 9639
rect 3786 9636 3792 9648
rect 3682 9608 3792 9636
rect 3682 9605 3694 9608
rect 3636 9599 3694 9605
rect 3786 9596 3792 9608
rect 3844 9596 3850 9648
rect 3970 9528 3976 9580
rect 4028 9568 4034 9580
rect 4157 9571 4215 9577
rect 4157 9568 4169 9571
rect 4028 9540 4169 9568
rect 4028 9528 4034 9540
rect 4157 9537 4169 9540
rect 4203 9537 4215 9571
rect 4356 9568 4384 9664
rect 4893 9639 4951 9645
rect 4893 9605 4905 9639
rect 4939 9636 4951 9639
rect 5534 9636 5540 9648
rect 4939 9608 5540 9636
rect 4939 9605 4951 9608
rect 4893 9599 4951 9605
rect 5534 9596 5540 9608
rect 5592 9636 5598 9648
rect 5718 9636 5724 9648
rect 5592 9608 5724 9636
rect 5592 9596 5598 9608
rect 5718 9596 5724 9608
rect 5776 9596 5782 9648
rect 5813 9639 5871 9645
rect 5813 9605 5825 9639
rect 5859 9636 5871 9639
rect 6840 9636 6868 9676
rect 7834 9664 7840 9716
rect 7892 9704 7898 9716
rect 8205 9707 8263 9713
rect 8205 9704 8217 9707
rect 7892 9676 8217 9704
rect 7892 9664 7898 9676
rect 8205 9673 8217 9676
rect 8251 9673 8263 9707
rect 8205 9667 8263 9673
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 10502 9704 10508 9716
rect 9824 9676 10508 9704
rect 9824 9664 9830 9676
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 12989 9707 13047 9713
rect 12989 9673 13001 9707
rect 13035 9704 13047 9707
rect 13354 9704 13360 9716
rect 13035 9676 13360 9704
rect 13035 9673 13047 9676
rect 12989 9667 13047 9673
rect 13354 9664 13360 9676
rect 13412 9664 13418 9716
rect 14001 9707 14059 9713
rect 14001 9673 14013 9707
rect 14047 9704 14059 9707
rect 14826 9704 14832 9716
rect 14047 9676 14832 9704
rect 14047 9673 14059 9676
rect 14001 9667 14059 9673
rect 14826 9664 14832 9676
rect 14884 9664 14890 9716
rect 20622 9664 20628 9716
rect 20680 9664 20686 9716
rect 20990 9664 20996 9716
rect 21048 9664 21054 9716
rect 21376 9676 22048 9704
rect 5859 9608 6040 9636
rect 6840 9608 11192 9636
rect 5859 9605 5871 9608
rect 5813 9599 5871 9605
rect 4614 9568 4620 9580
rect 4356 9540 4620 9568
rect 4157 9531 4215 9537
rect 4614 9528 4620 9540
rect 4672 9568 4678 9580
rect 6012 9568 6040 9608
rect 6362 9568 6368 9580
rect 4672 9540 5120 9568
rect 6012 9540 6368 9568
rect 4672 9528 4678 9540
rect 3878 9460 3884 9512
rect 3936 9460 3942 9512
rect 4246 9500 4252 9512
rect 3988 9472 4252 9500
rect 3988 9432 4016 9472
rect 4246 9460 4252 9472
rect 4304 9460 4310 9512
rect 5092 9509 5120 9540
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 6638 9528 6644 9580
rect 6696 9528 6702 9580
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 6825 9571 6883 9577
rect 6825 9568 6837 9571
rect 6788 9540 6837 9568
rect 6788 9528 6794 9540
rect 6825 9537 6837 9540
rect 6871 9537 6883 9571
rect 6825 9531 6883 9537
rect 7092 9571 7150 9577
rect 7092 9537 7104 9571
rect 7138 9568 7150 9571
rect 7374 9568 7380 9580
rect 7138 9540 7380 9568
rect 7138 9537 7150 9540
rect 7092 9531 7150 9537
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 8656 9571 8714 9577
rect 8656 9537 8668 9571
rect 8702 9568 8714 9571
rect 8938 9568 8944 9580
rect 8702 9540 8944 9568
rect 8702 9537 8714 9540
rect 8656 9531 8714 9537
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 11054 9528 11060 9580
rect 11112 9577 11118 9580
rect 11112 9531 11124 9577
rect 11164 9568 11192 9608
rect 11698 9596 11704 9648
rect 11756 9636 11762 9648
rect 11854 9639 11912 9645
rect 11854 9636 11866 9639
rect 11756 9608 11866 9636
rect 11756 9596 11762 9608
rect 11854 9605 11866 9608
rect 11900 9605 11912 9639
rect 11854 9599 11912 9605
rect 14366 9596 14372 9648
rect 14424 9636 14430 9648
rect 20346 9636 20352 9648
rect 14424 9608 20352 9636
rect 14424 9596 14430 9608
rect 20346 9596 20352 9608
rect 20404 9596 20410 9648
rect 20714 9596 20720 9648
rect 20772 9636 20778 9648
rect 21376 9636 21404 9676
rect 20772 9608 21404 9636
rect 22020 9636 22048 9676
rect 22554 9664 22560 9716
rect 22612 9704 22618 9716
rect 23290 9704 23296 9716
rect 22612 9676 23296 9704
rect 22612 9664 22618 9676
rect 23290 9664 23296 9676
rect 23348 9664 23354 9716
rect 24302 9704 24308 9716
rect 23400 9676 24308 9704
rect 22462 9636 22468 9648
rect 22020 9608 22468 9636
rect 20772 9596 20778 9608
rect 22462 9596 22468 9608
rect 22520 9596 22526 9648
rect 22646 9596 22652 9648
rect 22704 9636 22710 9648
rect 23400 9636 23428 9676
rect 24302 9664 24308 9676
rect 24360 9664 24366 9716
rect 25685 9707 25743 9713
rect 25685 9704 25697 9707
rect 25148 9676 25697 9704
rect 22704 9608 23428 9636
rect 22704 9596 22710 9608
rect 23474 9596 23480 9648
rect 23532 9636 23538 9648
rect 23532 9608 24164 9636
rect 23532 9596 23538 9608
rect 24136 9580 24164 9608
rect 24210 9596 24216 9648
rect 24268 9596 24274 9648
rect 25148 9636 25176 9676
rect 25685 9673 25697 9676
rect 25731 9704 25743 9707
rect 26697 9707 26755 9713
rect 26697 9704 26709 9707
rect 25731 9676 26709 9704
rect 25731 9673 25743 9676
rect 25685 9667 25743 9673
rect 26697 9673 26709 9676
rect 26743 9704 26755 9707
rect 28445 9707 28503 9713
rect 26743 9676 26832 9704
rect 26743 9673 26755 9676
rect 26697 9667 26755 9673
rect 24964 9608 25176 9636
rect 14829 9571 14887 9577
rect 11164 9540 13676 9568
rect 11112 9528 11118 9531
rect 4985 9503 5043 9509
rect 4985 9469 4997 9503
rect 5031 9469 5043 9503
rect 4985 9463 5043 9469
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9469 5135 9503
rect 5077 9463 5135 9469
rect 3896 9404 4016 9432
rect 2501 9367 2559 9373
rect 2501 9333 2513 9367
rect 2547 9364 2559 9367
rect 3896 9364 3924 9404
rect 4062 9392 4068 9444
rect 4120 9432 4126 9444
rect 4525 9435 4583 9441
rect 4525 9432 4537 9435
rect 4120 9404 4537 9432
rect 4120 9392 4126 9404
rect 4525 9401 4537 9404
rect 4571 9401 4583 9435
rect 5000 9432 5028 9463
rect 5902 9460 5908 9512
rect 5960 9460 5966 9512
rect 6086 9460 6092 9512
rect 6144 9500 6150 9512
rect 6144 9472 6500 9500
rect 6144 9460 6150 9472
rect 5920 9432 5948 9460
rect 6472 9441 6500 9472
rect 8202 9460 8208 9512
rect 8260 9500 8266 9512
rect 8389 9503 8447 9509
rect 8389 9500 8401 9503
rect 8260 9472 8401 9500
rect 8260 9460 8266 9472
rect 8389 9469 8401 9472
rect 8435 9469 8447 9503
rect 8389 9463 8447 9469
rect 11333 9503 11391 9509
rect 11333 9469 11345 9503
rect 11379 9500 11391 9503
rect 11514 9500 11520 9512
rect 11379 9472 11520 9500
rect 11379 9469 11391 9472
rect 11333 9463 11391 9469
rect 11514 9460 11520 9472
rect 11572 9500 11578 9512
rect 11609 9503 11667 9509
rect 11609 9500 11621 9503
rect 11572 9472 11621 9500
rect 11572 9460 11578 9472
rect 11609 9469 11621 9472
rect 11655 9469 11667 9503
rect 13648 9500 13676 9540
rect 14829 9537 14841 9571
rect 14875 9568 14887 9571
rect 15194 9568 15200 9580
rect 14875 9540 15200 9568
rect 14875 9537 14887 9540
rect 14829 9531 14887 9537
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 15470 9528 15476 9580
rect 15528 9568 15534 9580
rect 17678 9577 17684 9580
rect 17405 9571 17463 9577
rect 17405 9568 17417 9571
rect 15528 9540 17417 9568
rect 15528 9528 15534 9540
rect 17405 9537 17417 9540
rect 17451 9537 17463 9571
rect 17405 9531 17463 9537
rect 17672 9531 17684 9577
rect 17678 9528 17684 9531
rect 17736 9528 17742 9580
rect 19886 9528 19892 9580
rect 19944 9568 19950 9580
rect 20073 9571 20131 9577
rect 20073 9568 20085 9571
rect 19944 9540 20085 9568
rect 19944 9528 19950 9540
rect 20073 9537 20085 9540
rect 20119 9537 20131 9571
rect 20073 9531 20131 9537
rect 20441 9571 20499 9577
rect 20441 9537 20453 9571
rect 20487 9537 20499 9571
rect 20441 9531 20499 9537
rect 14921 9503 14979 9509
rect 14921 9500 14933 9503
rect 13648 9472 14933 9500
rect 11609 9463 11667 9469
rect 14921 9469 14933 9472
rect 14967 9469 14979 9503
rect 16758 9500 16764 9512
rect 14921 9463 14979 9469
rect 15028 9472 16764 9500
rect 5000 9404 5948 9432
rect 4525 9395 4583 9401
rect 2547 9336 3924 9364
rect 2547 9333 2559 9336
rect 2501 9327 2559 9333
rect 3970 9324 3976 9376
rect 4028 9324 4034 9376
rect 5442 9324 5448 9376
rect 5500 9324 5506 9376
rect 5920 9364 5948 9404
rect 6457 9435 6515 9441
rect 6457 9401 6469 9435
rect 6503 9401 6515 9435
rect 6457 9395 6515 9401
rect 9398 9392 9404 9444
rect 9456 9432 9462 9444
rect 15028 9432 15056 9472
rect 16758 9460 16764 9472
rect 16816 9460 16822 9512
rect 9456 9404 10272 9432
rect 9456 9392 9462 9404
rect 7466 9364 7472 9376
rect 5920 9336 7472 9364
rect 7466 9324 7472 9336
rect 7524 9324 7530 9376
rect 9953 9367 10011 9373
rect 9953 9333 9965 9367
rect 9999 9364 10011 9367
rect 10134 9364 10140 9376
rect 9999 9336 10140 9364
rect 9999 9333 10011 9336
rect 9953 9327 10011 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10244 9364 10272 9404
rect 12728 9404 15056 9432
rect 12728 9364 12756 9404
rect 18782 9392 18788 9444
rect 18840 9392 18846 9444
rect 10244 9336 12756 9364
rect 14918 9324 14924 9376
rect 14976 9324 14982 9376
rect 15197 9367 15255 9373
rect 15197 9333 15209 9367
rect 15243 9364 15255 9367
rect 19978 9364 19984 9376
rect 15243 9336 19984 9364
rect 15243 9333 15255 9336
rect 15197 9327 15255 9333
rect 19978 9324 19984 9336
rect 20036 9324 20042 9376
rect 20088 9364 20116 9531
rect 20456 9432 20484 9531
rect 22370 9528 22376 9580
rect 22428 9568 22434 9580
rect 22925 9571 22983 9577
rect 22925 9568 22937 9571
rect 22428 9540 22937 9568
rect 22428 9528 22434 9540
rect 22925 9537 22937 9540
rect 22971 9568 22983 9571
rect 23014 9568 23020 9580
rect 22971 9540 23020 9568
rect 22971 9537 22983 9540
rect 22925 9531 22983 9537
rect 23014 9528 23020 9540
rect 23072 9528 23078 9580
rect 23198 9528 23204 9580
rect 23256 9528 23262 9580
rect 23566 9528 23572 9580
rect 23624 9568 23630 9580
rect 24029 9571 24087 9577
rect 24029 9568 24041 9571
rect 23624 9540 24041 9568
rect 23624 9528 23630 9540
rect 24029 9537 24041 9540
rect 24075 9537 24087 9571
rect 24029 9531 24087 9537
rect 24118 9528 24124 9580
rect 24176 9528 24182 9580
rect 24305 9571 24363 9577
rect 24305 9537 24317 9571
rect 24351 9568 24363 9571
rect 24394 9568 24400 9580
rect 24351 9540 24400 9568
rect 24351 9537 24363 9540
rect 24305 9531 24363 9537
rect 24394 9528 24400 9540
rect 24452 9528 24458 9580
rect 24581 9571 24639 9577
rect 24581 9537 24593 9571
rect 24627 9568 24639 9571
rect 24857 9571 24915 9577
rect 24857 9568 24869 9571
rect 24627 9540 24869 9568
rect 24627 9537 24639 9540
rect 24581 9531 24639 9537
rect 24857 9537 24869 9540
rect 24903 9537 24915 9571
rect 24857 9531 24915 9537
rect 20530 9460 20536 9512
rect 20588 9500 20594 9512
rect 20990 9500 20996 9512
rect 20588 9472 20996 9500
rect 20588 9460 20594 9472
rect 20990 9460 20996 9472
rect 21048 9500 21054 9512
rect 21085 9503 21143 9509
rect 21085 9500 21097 9503
rect 21048 9472 21097 9500
rect 21048 9460 21054 9472
rect 21085 9469 21097 9472
rect 21131 9469 21143 9503
rect 21085 9463 21143 9469
rect 21269 9503 21327 9509
rect 21269 9469 21281 9503
rect 21315 9500 21327 9503
rect 21818 9500 21824 9512
rect 21315 9472 21824 9500
rect 21315 9469 21327 9472
rect 21269 9463 21327 9469
rect 21818 9460 21824 9472
rect 21876 9460 21882 9512
rect 23216 9500 23244 9528
rect 24596 9500 24624 9531
rect 24964 9500 24992 9608
rect 25222 9596 25228 9648
rect 25280 9596 25286 9648
rect 25501 9639 25559 9645
rect 25501 9605 25513 9639
rect 25547 9636 25559 9639
rect 26602 9636 26608 9648
rect 25547 9608 26608 9636
rect 25547 9605 25559 9608
rect 25501 9599 25559 9605
rect 26602 9596 26608 9608
rect 26660 9596 26666 9648
rect 25041 9571 25099 9577
rect 25041 9537 25053 9571
rect 25087 9537 25099 9571
rect 25041 9531 25099 9537
rect 23216 9472 24624 9500
rect 24688 9472 24992 9500
rect 25056 9500 25084 9531
rect 25130 9528 25136 9580
rect 25188 9528 25194 9580
rect 25314 9528 25320 9580
rect 25372 9568 25378 9580
rect 25409 9571 25467 9577
rect 25409 9568 25421 9571
rect 25372 9540 25421 9568
rect 25372 9528 25378 9540
rect 25409 9537 25421 9540
rect 25455 9537 25467 9571
rect 25409 9531 25467 9537
rect 25593 9571 25651 9577
rect 25593 9537 25605 9571
rect 25639 9537 25651 9571
rect 25593 9531 25651 9537
rect 25332 9500 25360 9528
rect 25056 9472 25360 9500
rect 23106 9432 23112 9444
rect 20456 9404 23112 9432
rect 23106 9392 23112 9404
rect 23164 9392 23170 9444
rect 23201 9435 23259 9441
rect 23201 9401 23213 9435
rect 23247 9401 23259 9435
rect 23201 9395 23259 9401
rect 21453 9367 21511 9373
rect 21453 9364 21465 9367
rect 20088 9336 21465 9364
rect 21453 9333 21465 9336
rect 21499 9364 21511 9367
rect 22094 9364 22100 9376
rect 21499 9336 22100 9364
rect 21499 9333 21511 9336
rect 21453 9327 21511 9333
rect 22094 9324 22100 9336
rect 22152 9324 22158 9376
rect 22646 9324 22652 9376
rect 22704 9364 22710 9376
rect 23216 9364 23244 9395
rect 24026 9392 24032 9444
rect 24084 9432 24090 9444
rect 24688 9441 24716 9472
rect 25498 9460 25504 9512
rect 25556 9500 25562 9512
rect 25608 9500 25636 9531
rect 26510 9528 26516 9580
rect 26568 9528 26574 9580
rect 26804 9568 26832 9676
rect 28445 9673 28457 9707
rect 28491 9673 28503 9707
rect 28445 9667 28503 9673
rect 31113 9707 31171 9713
rect 31113 9673 31125 9707
rect 31159 9704 31171 9707
rect 31202 9704 31208 9716
rect 31159 9676 31208 9704
rect 31159 9673 31171 9676
rect 31113 9667 31171 9673
rect 26878 9596 26884 9648
rect 26936 9636 26942 9648
rect 27614 9636 27620 9648
rect 26936 9608 27620 9636
rect 26936 9596 26942 9608
rect 27614 9596 27620 9608
rect 27672 9596 27678 9648
rect 28460 9636 28488 9667
rect 31202 9664 31208 9676
rect 31260 9664 31266 9716
rect 28902 9636 28908 9648
rect 28460 9608 28908 9636
rect 28902 9596 28908 9608
rect 28960 9636 28966 9648
rect 30285 9639 30343 9645
rect 30285 9636 30297 9639
rect 28960 9608 30297 9636
rect 28960 9596 28966 9608
rect 30285 9605 30297 9608
rect 30331 9605 30343 9639
rect 30285 9599 30343 9605
rect 27065 9571 27123 9577
rect 27065 9568 27077 9571
rect 26804 9540 27077 9568
rect 27065 9537 27077 9540
rect 27111 9537 27123 9571
rect 27065 9531 27123 9537
rect 27525 9571 27583 9577
rect 27525 9537 27537 9571
rect 27571 9537 27583 9571
rect 27525 9531 27583 9537
rect 28169 9571 28227 9577
rect 28169 9537 28181 9571
rect 28215 9568 28227 9571
rect 28258 9568 28264 9580
rect 28215 9540 28264 9568
rect 28215 9537 28227 9540
rect 28169 9531 28227 9537
rect 25556 9472 25636 9500
rect 26528 9500 26556 9528
rect 27540 9500 27568 9531
rect 28258 9528 28264 9540
rect 28316 9528 28322 9580
rect 29569 9571 29627 9577
rect 29569 9537 29581 9571
rect 29615 9568 29627 9571
rect 29615 9540 29776 9568
rect 29615 9537 29627 9540
rect 29569 9531 29627 9537
rect 26528 9472 27568 9500
rect 25556 9460 25562 9472
rect 27798 9460 27804 9512
rect 27856 9500 27862 9512
rect 28353 9503 28411 9509
rect 28353 9500 28365 9503
rect 27856 9472 28365 9500
rect 27856 9460 27862 9472
rect 28353 9469 28365 9472
rect 28399 9469 28411 9503
rect 29748 9500 29776 9540
rect 29822 9528 29828 9580
rect 29880 9528 29886 9580
rect 34054 9528 34060 9580
rect 34112 9528 34118 9580
rect 34238 9528 34244 9580
rect 34296 9528 34302 9580
rect 34333 9571 34391 9577
rect 34333 9537 34345 9571
rect 34379 9568 34391 9571
rect 34422 9568 34428 9580
rect 34379 9540 34428 9568
rect 34379 9537 34391 9540
rect 34333 9531 34391 9537
rect 34422 9528 34428 9540
rect 34480 9528 34486 9580
rect 29748 9472 29960 9500
rect 28353 9463 28411 9469
rect 24673 9435 24731 9441
rect 24673 9432 24685 9435
rect 24084 9404 24685 9432
rect 24084 9392 24090 9404
rect 24673 9401 24685 9404
rect 24719 9401 24731 9435
rect 24673 9395 24731 9401
rect 24857 9435 24915 9441
rect 24857 9401 24869 9435
rect 24903 9432 24915 9435
rect 25406 9432 25412 9444
rect 24903 9404 25412 9432
rect 24903 9401 24915 9404
rect 24857 9395 24915 9401
rect 25406 9392 25412 9404
rect 25464 9392 25470 9444
rect 26326 9392 26332 9444
rect 26384 9432 26390 9444
rect 27709 9435 27767 9441
rect 27709 9432 27721 9435
rect 26384 9404 27721 9432
rect 26384 9392 26390 9404
rect 27709 9401 27721 9404
rect 27755 9432 27767 9435
rect 28166 9432 28172 9444
rect 27755 9404 28172 9432
rect 27755 9401 27767 9404
rect 27709 9395 27767 9401
rect 28166 9392 28172 9404
rect 28224 9392 28230 9444
rect 29932 9441 29960 9472
rect 30282 9460 30288 9512
rect 30340 9500 30346 9512
rect 30377 9503 30435 9509
rect 30377 9500 30389 9503
rect 30340 9472 30389 9500
rect 30340 9460 30346 9472
rect 30377 9469 30389 9472
rect 30423 9469 30435 9503
rect 30377 9463 30435 9469
rect 30466 9460 30472 9512
rect 30524 9500 30530 9512
rect 30745 9503 30803 9509
rect 30745 9500 30757 9503
rect 30524 9472 30757 9500
rect 30524 9460 30530 9472
rect 30745 9469 30757 9472
rect 30791 9469 30803 9503
rect 30745 9463 30803 9469
rect 29917 9435 29975 9441
rect 29917 9401 29929 9435
rect 29963 9401 29975 9435
rect 29917 9395 29975 9401
rect 23477 9367 23535 9373
rect 23477 9364 23489 9367
rect 22704 9336 23489 9364
rect 22704 9324 22710 9336
rect 23477 9333 23489 9336
rect 23523 9364 23535 9367
rect 23750 9364 23756 9376
rect 23523 9336 23756 9364
rect 23523 9333 23535 9336
rect 23477 9327 23535 9333
rect 23750 9324 23756 9336
rect 23808 9324 23814 9376
rect 23842 9324 23848 9376
rect 23900 9324 23906 9376
rect 24118 9324 24124 9376
rect 24176 9364 24182 9376
rect 25498 9364 25504 9376
rect 24176 9336 25504 9364
rect 24176 9324 24182 9336
rect 25498 9324 25504 9336
rect 25556 9324 25562 9376
rect 26786 9324 26792 9376
rect 26844 9364 26850 9376
rect 27157 9367 27215 9373
rect 27157 9364 27169 9367
rect 26844 9336 27169 9364
rect 26844 9324 26850 9336
rect 27157 9333 27169 9336
rect 27203 9364 27215 9367
rect 27798 9364 27804 9376
rect 27203 9336 27804 9364
rect 27203 9333 27215 9336
rect 27157 9327 27215 9333
rect 27798 9324 27804 9336
rect 27856 9324 27862 9376
rect 27985 9367 28043 9373
rect 27985 9333 27997 9367
rect 28031 9364 28043 9367
rect 28074 9364 28080 9376
rect 28031 9336 28080 9364
rect 28031 9333 28043 9336
rect 27985 9327 28043 9333
rect 28074 9324 28080 9336
rect 28132 9324 28138 9376
rect 33042 9324 33048 9376
rect 33100 9364 33106 9376
rect 33873 9367 33931 9373
rect 33873 9364 33885 9367
rect 33100 9336 33885 9364
rect 33100 9324 33106 9336
rect 33873 9333 33885 9336
rect 33919 9333 33931 9367
rect 33873 9327 33931 9333
rect 1104 9274 35328 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 35328 9274
rect 1104 9200 35328 9222
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 4706 9160 4712 9172
rect 1627 9132 4712 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 5169 9163 5227 9169
rect 5169 9129 5181 9163
rect 5215 9160 5227 9163
rect 5534 9160 5540 9172
rect 5215 9132 5540 9160
rect 5215 9129 5227 9132
rect 5169 9123 5227 9129
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 6362 9120 6368 9172
rect 6420 9160 6426 9172
rect 6641 9163 6699 9169
rect 6641 9160 6653 9163
rect 6420 9132 6653 9160
rect 6420 9120 6426 9132
rect 6641 9129 6653 9132
rect 6687 9129 6699 9163
rect 6641 9123 6699 9129
rect 7374 9120 7380 9172
rect 7432 9120 7438 9172
rect 8938 9120 8944 9172
rect 8996 9120 9002 9172
rect 10042 9120 10048 9172
rect 10100 9120 10106 9172
rect 10321 9163 10379 9169
rect 10321 9129 10333 9163
rect 10367 9160 10379 9163
rect 10367 9132 11008 9160
rect 10367 9129 10379 9132
rect 10321 9123 10379 9129
rect 8297 9095 8355 9101
rect 8297 9092 8309 9095
rect 8036 9064 8309 9092
rect 6638 8984 6644 9036
rect 6696 9024 6702 9036
rect 8036 9033 8064 9064
rect 8297 9061 8309 9064
rect 8343 9092 8355 9095
rect 9398 9092 9404 9104
rect 8343 9064 9404 9092
rect 8343 9061 8355 9064
rect 8297 9055 8355 9061
rect 9398 9052 9404 9064
rect 9456 9052 9462 9104
rect 10980 9092 11008 9132
rect 11054 9120 11060 9172
rect 11112 9160 11118 9172
rect 11149 9163 11207 9169
rect 11149 9160 11161 9163
rect 11112 9132 11161 9160
rect 11112 9120 11118 9132
rect 11149 9129 11161 9132
rect 11195 9129 11207 9163
rect 11149 9123 11207 9129
rect 13078 9120 13084 9172
rect 13136 9160 13142 9172
rect 13630 9160 13636 9172
rect 13136 9132 13636 9160
rect 13136 9120 13142 9132
rect 13630 9120 13636 9132
rect 13688 9120 13694 9172
rect 14918 9120 14924 9172
rect 14976 9120 14982 9172
rect 17678 9120 17684 9172
rect 17736 9160 17742 9172
rect 17773 9163 17831 9169
rect 17773 9160 17785 9163
rect 17736 9132 17785 9160
rect 17736 9120 17742 9132
rect 17773 9129 17785 9132
rect 17819 9129 17831 9163
rect 17773 9123 17831 9129
rect 19978 9120 19984 9172
rect 20036 9160 20042 9172
rect 21818 9160 21824 9172
rect 20036 9132 21824 9160
rect 20036 9120 20042 9132
rect 21818 9120 21824 9132
rect 21876 9120 21882 9172
rect 22002 9120 22008 9172
rect 22060 9160 22066 9172
rect 22646 9160 22652 9172
rect 22060 9132 22652 9160
rect 22060 9120 22066 9132
rect 22646 9120 22652 9132
rect 22704 9120 22710 9172
rect 23017 9163 23075 9169
rect 23017 9160 23029 9163
rect 22756 9132 23029 9160
rect 15562 9092 15568 9104
rect 10980 9064 15568 9092
rect 15562 9052 15568 9064
rect 15620 9052 15626 9104
rect 20625 9095 20683 9101
rect 20625 9061 20637 9095
rect 20671 9061 20683 9095
rect 22756 9092 22784 9132
rect 23017 9129 23029 9132
rect 23063 9129 23075 9163
rect 23017 9123 23075 9129
rect 25225 9163 25283 9169
rect 25225 9129 25237 9163
rect 25271 9160 25283 9163
rect 25314 9160 25320 9172
rect 25271 9132 25320 9160
rect 25271 9129 25283 9132
rect 25225 9123 25283 9129
rect 25314 9120 25320 9132
rect 25372 9120 25378 9172
rect 28537 9163 28595 9169
rect 28537 9129 28549 9163
rect 28583 9160 28595 9163
rect 29270 9160 29276 9172
rect 28583 9132 29276 9160
rect 28583 9129 28595 9132
rect 28537 9123 28595 9129
rect 29270 9120 29276 9132
rect 29328 9120 29334 9172
rect 34238 9120 34244 9172
rect 34296 9160 34302 9172
rect 34517 9163 34575 9169
rect 34517 9160 34529 9163
rect 34296 9132 34529 9160
rect 34296 9120 34302 9132
rect 34517 9129 34529 9132
rect 34563 9129 34575 9163
rect 34517 9123 34575 9129
rect 20625 9055 20683 9061
rect 22020 9064 22784 9092
rect 22848 9064 23152 9092
rect 8021 9027 8079 9033
rect 6696 8996 6868 9024
rect 6696 8984 6702 8996
rect 6840 8968 6868 8996
rect 8021 8993 8033 9027
rect 8067 8993 8079 9027
rect 8021 8987 8079 8993
rect 9585 9027 9643 9033
rect 9585 8993 9597 9027
rect 9631 9024 9643 9027
rect 9674 9024 9680 9036
rect 9631 8996 9680 9024
rect 9631 8993 9643 8996
rect 9585 8987 9643 8993
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 10226 9024 10232 9036
rect 9968 8996 10232 9024
rect 1302 8916 1308 8968
rect 1360 8956 1366 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 1360 8928 1409 8956
rect 1360 8916 1366 8928
rect 1397 8925 1409 8928
rect 1443 8956 1455 8959
rect 1673 8959 1731 8965
rect 1673 8956 1685 8959
rect 1443 8928 1685 8956
rect 1443 8925 1455 8928
rect 1397 8919 1455 8925
rect 1673 8925 1685 8928
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8956 3847 8959
rect 3878 8956 3884 8968
rect 3835 8928 3884 8956
rect 3835 8925 3847 8928
rect 3789 8919 3847 8925
rect 3878 8916 3884 8928
rect 3936 8916 3942 8968
rect 4062 8965 4068 8968
rect 4056 8956 4068 8965
rect 4023 8928 4068 8956
rect 4056 8919 4068 8928
rect 4062 8916 4068 8919
rect 4120 8916 4126 8968
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8925 5319 8959
rect 5261 8919 5319 8925
rect 5528 8959 5586 8965
rect 5528 8925 5540 8959
rect 5574 8925 5586 8959
rect 5528 8919 5586 8925
rect 5276 8820 5304 8919
rect 5442 8848 5448 8900
rect 5500 8888 5506 8900
rect 5552 8888 5580 8919
rect 6822 8916 6828 8968
rect 6880 8916 6886 8968
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8956 7803 8959
rect 7834 8956 7840 8968
rect 7791 8928 7840 8956
rect 7791 8925 7803 8928
rect 7745 8919 7803 8925
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 9309 8959 9367 8965
rect 9309 8925 9321 8959
rect 9355 8956 9367 8959
rect 9766 8956 9772 8968
rect 9355 8928 9772 8956
rect 9355 8925 9367 8928
rect 9309 8919 9367 8925
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 9968 8965 9996 8996
rect 10226 8984 10232 8996
rect 10284 8984 10290 9036
rect 10502 8984 10508 9036
rect 10560 8984 10566 9036
rect 13449 9027 13507 9033
rect 13449 9024 13461 9027
rect 13188 8996 13461 9024
rect 9953 8959 10011 8965
rect 9953 8925 9965 8959
rect 9999 8925 10011 8959
rect 9953 8919 10011 8925
rect 10042 8916 10048 8968
rect 10100 8916 10106 8968
rect 10134 8916 10140 8968
rect 10192 8956 10198 8968
rect 10781 8959 10839 8965
rect 10781 8956 10793 8959
rect 10192 8928 10793 8956
rect 10192 8916 10198 8928
rect 10781 8925 10793 8928
rect 10827 8925 10839 8959
rect 10781 8919 10839 8925
rect 12710 8916 12716 8968
rect 12768 8916 12774 8968
rect 12802 8916 12808 8968
rect 12860 8956 12866 8968
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 12860 8928 13001 8956
rect 12860 8916 12866 8928
rect 12989 8925 13001 8928
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 13078 8916 13084 8968
rect 13136 8916 13142 8968
rect 10689 8891 10747 8897
rect 10689 8888 10701 8891
rect 5500 8860 5580 8888
rect 9600 8860 10701 8888
rect 5500 8848 5506 8860
rect 9600 8832 9628 8860
rect 10689 8857 10701 8860
rect 10735 8857 10747 8891
rect 10689 8851 10747 8857
rect 10870 8848 10876 8900
rect 10928 8888 10934 8900
rect 12897 8891 12955 8897
rect 12897 8888 12909 8891
rect 10928 8860 12909 8888
rect 10928 8848 10934 8860
rect 12897 8857 12909 8860
rect 12943 8888 12955 8891
rect 13188 8888 13216 8996
rect 13449 8993 13461 8996
rect 13495 9024 13507 9027
rect 16390 9024 16396 9036
rect 13495 8996 16396 9024
rect 13495 8993 13507 8996
rect 13449 8987 13507 8993
rect 16390 8984 16396 8996
rect 16448 8984 16454 9036
rect 16850 8984 16856 9036
rect 16908 9024 16914 9036
rect 18322 9024 18328 9036
rect 16908 8996 18328 9024
rect 16908 8984 16914 8996
rect 18322 8984 18328 8996
rect 18380 9024 18386 9036
rect 18601 9027 18659 9033
rect 18601 9024 18613 9027
rect 18380 8996 18613 9024
rect 18380 8984 18386 8996
rect 18601 8993 18613 8996
rect 18647 8993 18659 9027
rect 20640 9024 20668 9055
rect 22020 9036 22048 9064
rect 20806 9024 20812 9036
rect 20640 8996 20812 9024
rect 18601 8987 18659 8993
rect 20806 8984 20812 8996
rect 20864 9024 20870 9036
rect 20864 8996 20944 9024
rect 20864 8984 20870 8996
rect 14458 8965 14464 8968
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 12943 8860 13216 8888
rect 13372 8928 14289 8956
rect 12943 8857 12955 8860
rect 12897 8851 12955 8857
rect 6730 8820 6736 8832
rect 5276 8792 6736 8820
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 7466 8780 7472 8832
rect 7524 8820 7530 8832
rect 7742 8820 7748 8832
rect 7524 8792 7748 8820
rect 7524 8780 7530 8792
rect 7742 8780 7748 8792
rect 7800 8820 7806 8832
rect 7837 8823 7895 8829
rect 7837 8820 7849 8823
rect 7800 8792 7849 8820
rect 7800 8780 7806 8792
rect 7837 8789 7849 8792
rect 7883 8789 7895 8823
rect 7837 8783 7895 8789
rect 9401 8823 9459 8829
rect 9401 8789 9413 8823
rect 9447 8820 9459 8823
rect 9582 8820 9588 8832
rect 9447 8792 9588 8820
rect 9447 8789 9459 8792
rect 9401 8783 9459 8789
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 9861 8823 9919 8829
rect 9861 8820 9873 8823
rect 9732 8792 9873 8820
rect 9732 8780 9738 8792
rect 9861 8789 9873 8792
rect 9907 8820 9919 8823
rect 10318 8820 10324 8832
rect 9907 8792 10324 8820
rect 9907 8789 9919 8792
rect 9861 8783 9919 8789
rect 10318 8780 10324 8792
rect 10376 8780 10382 8832
rect 10502 8780 10508 8832
rect 10560 8820 10566 8832
rect 10778 8820 10784 8832
rect 10560 8792 10784 8820
rect 10560 8780 10566 8792
rect 10778 8780 10784 8792
rect 10836 8820 10842 8832
rect 11241 8823 11299 8829
rect 11241 8820 11253 8823
rect 10836 8792 11253 8820
rect 10836 8780 10842 8792
rect 11241 8789 11253 8792
rect 11287 8789 11299 8823
rect 11241 8783 11299 8789
rect 11330 8780 11336 8832
rect 11388 8820 11394 8832
rect 13170 8820 13176 8832
rect 11388 8792 13176 8820
rect 11388 8780 11394 8792
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 13265 8823 13323 8829
rect 13265 8789 13277 8823
rect 13311 8820 13323 8823
rect 13372 8820 13400 8928
rect 14277 8925 14289 8928
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 14425 8959 14464 8965
rect 14425 8925 14437 8959
rect 14425 8919 14464 8925
rect 14458 8916 14464 8919
rect 14516 8916 14522 8968
rect 14642 8916 14648 8968
rect 14700 8916 14706 8968
rect 14781 8959 14839 8965
rect 14781 8925 14793 8959
rect 14827 8956 14839 8959
rect 15010 8956 15016 8968
rect 14827 8928 15016 8956
rect 14827 8925 14839 8928
rect 14781 8919 14839 8925
rect 15010 8916 15016 8928
rect 15068 8956 15074 8968
rect 15105 8959 15163 8965
rect 15105 8956 15117 8959
rect 15068 8928 15117 8956
rect 15068 8916 15074 8928
rect 15105 8925 15117 8928
rect 15151 8956 15163 8959
rect 17862 8956 17868 8968
rect 15151 8928 17868 8956
rect 15151 8925 15163 8928
rect 15105 8919 15163 8925
rect 17862 8916 17868 8928
rect 17920 8916 17926 8968
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8956 18291 8959
rect 18782 8956 18788 8968
rect 18279 8928 18788 8956
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 18782 8916 18788 8928
rect 18840 8916 18846 8968
rect 18874 8916 18880 8968
rect 18932 8956 18938 8968
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 18932 8928 19257 8956
rect 18932 8916 18938 8928
rect 19245 8925 19257 8928
rect 19291 8925 19303 8959
rect 20714 8956 20720 8968
rect 19245 8919 19303 8925
rect 19444 8928 20720 8956
rect 13998 8848 14004 8900
rect 14056 8888 14062 8900
rect 14553 8891 14611 8897
rect 14553 8888 14565 8891
rect 14056 8860 14565 8888
rect 14056 8848 14062 8860
rect 14553 8857 14565 8860
rect 14599 8888 14611 8891
rect 15289 8891 15347 8897
rect 15289 8888 15301 8891
rect 14599 8860 15301 8888
rect 14599 8857 14611 8860
rect 14553 8851 14611 8857
rect 15289 8857 15301 8860
rect 15335 8888 15347 8891
rect 19444 8888 19472 8928
rect 20714 8916 20720 8928
rect 20772 8916 20778 8968
rect 20916 8956 20944 8996
rect 20990 8984 20996 9036
rect 21048 9024 21054 9036
rect 21177 9027 21235 9033
rect 21177 9024 21189 9027
rect 21048 8996 21189 9024
rect 21048 8984 21054 8996
rect 21177 8993 21189 8996
rect 21223 8993 21235 9027
rect 21177 8987 21235 8993
rect 21266 8984 21272 9036
rect 21324 8984 21330 9036
rect 21818 8984 21824 9036
rect 21876 8984 21882 9036
rect 21913 9027 21971 9033
rect 21913 8993 21925 9027
rect 21959 9024 21971 9027
rect 22002 9024 22008 9036
rect 21959 8996 22008 9024
rect 21959 8993 21971 8996
rect 21913 8987 21971 8993
rect 22002 8984 22008 8996
rect 22060 8984 22066 9036
rect 22370 8984 22376 9036
rect 22428 9024 22434 9036
rect 22557 9027 22615 9033
rect 22557 9024 22569 9027
rect 22428 8996 22569 9024
rect 22428 8984 22434 8996
rect 22557 8993 22569 8996
rect 22603 8993 22615 9027
rect 22557 8987 22615 8993
rect 21085 8959 21143 8965
rect 21085 8956 21097 8959
rect 20916 8928 21097 8956
rect 21085 8925 21097 8928
rect 21131 8925 21143 8959
rect 21085 8919 21143 8925
rect 21545 8959 21603 8965
rect 21545 8925 21557 8959
rect 21591 8956 21603 8959
rect 21634 8956 21640 8968
rect 21591 8928 21640 8956
rect 21591 8925 21603 8928
rect 21545 8919 21603 8925
rect 21634 8916 21640 8928
rect 21692 8916 21698 8968
rect 21726 8916 21732 8968
rect 21784 8916 21790 8968
rect 22848 8965 22876 9064
rect 23124 9024 23152 9064
rect 24394 9052 24400 9104
rect 24452 9052 24458 9104
rect 24578 9052 24584 9104
rect 24636 9052 24642 9104
rect 27065 9095 27123 9101
rect 27065 9061 27077 9095
rect 27111 9061 27123 9095
rect 27065 9055 27123 9061
rect 24596 9024 24624 9052
rect 23124 8996 24808 9024
rect 22097 8959 22155 8965
rect 22097 8925 22109 8959
rect 22143 8925 22155 8959
rect 22097 8919 22155 8925
rect 22832 8959 22890 8965
rect 22832 8925 22844 8959
rect 22878 8925 22890 8959
rect 22832 8919 22890 8925
rect 22925 8959 22983 8965
rect 22925 8925 22937 8959
rect 22971 8958 22983 8959
rect 22971 8956 23060 8958
rect 23842 8956 23848 8968
rect 22971 8930 23848 8956
rect 22971 8925 22983 8930
rect 22925 8919 22983 8925
rect 23032 8928 23848 8930
rect 15335 8860 19472 8888
rect 19512 8891 19570 8897
rect 15335 8857 15347 8860
rect 15289 8851 15347 8857
rect 19512 8857 19524 8891
rect 19558 8888 19570 8891
rect 19558 8860 20760 8888
rect 19558 8857 19570 8860
rect 19512 8851 19570 8857
rect 13311 8792 13400 8820
rect 13311 8789 13323 8792
rect 13265 8783 13323 8789
rect 13446 8780 13452 8832
rect 13504 8820 13510 8832
rect 16850 8820 16856 8832
rect 13504 8792 16856 8820
rect 13504 8780 13510 8792
rect 16850 8780 16856 8792
rect 16908 8780 16914 8832
rect 16942 8780 16948 8832
rect 17000 8820 17006 8832
rect 18141 8823 18199 8829
rect 18141 8820 18153 8823
rect 17000 8792 18153 8820
rect 17000 8780 17006 8792
rect 18141 8789 18153 8792
rect 18187 8789 18199 8823
rect 18141 8783 18199 8789
rect 19150 8780 19156 8832
rect 19208 8820 19214 8832
rect 20622 8820 20628 8832
rect 19208 8792 20628 8820
rect 19208 8780 19214 8792
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 20732 8829 20760 8860
rect 21266 8848 21272 8900
rect 21324 8888 21330 8900
rect 22112 8888 22140 8919
rect 21324 8860 22140 8888
rect 22204 8860 22600 8888
rect 21324 8848 21330 8860
rect 20717 8823 20775 8829
rect 20717 8789 20729 8823
rect 20763 8789 20775 8823
rect 20717 8783 20775 8789
rect 21542 8780 21548 8832
rect 21600 8820 21606 8832
rect 22094 8820 22100 8832
rect 21600 8792 22100 8820
rect 21600 8780 21606 8792
rect 22094 8780 22100 8792
rect 22152 8820 22158 8832
rect 22204 8820 22232 8860
rect 22152 8792 22232 8820
rect 22152 8780 22158 8792
rect 22278 8780 22284 8832
rect 22336 8780 22342 8832
rect 22462 8780 22468 8832
rect 22520 8780 22526 8832
rect 22572 8820 22600 8860
rect 22646 8848 22652 8900
rect 22704 8888 22710 8900
rect 23032 8888 23060 8928
rect 23842 8916 23848 8928
rect 23900 8956 23906 8968
rect 24780 8965 24808 8996
rect 24854 8984 24860 9036
rect 24912 9024 24918 9036
rect 25685 9027 25743 9033
rect 25685 9024 25697 9027
rect 24912 8996 25697 9024
rect 24912 8984 24918 8996
rect 25685 8993 25697 8996
rect 25731 8993 25743 9027
rect 25685 8987 25743 8993
rect 24611 8959 24669 8965
rect 24611 8956 24623 8959
rect 23900 8928 24623 8956
rect 23900 8916 23906 8928
rect 24611 8925 24623 8928
rect 24657 8925 24669 8959
rect 24611 8919 24669 8925
rect 24758 8959 24816 8965
rect 24758 8925 24770 8959
rect 24804 8956 24816 8959
rect 27080 8956 27108 9055
rect 27154 9052 27160 9104
rect 27212 9092 27218 9104
rect 27212 9064 28672 9092
rect 27212 9052 27218 9064
rect 27246 8984 27252 9036
rect 27304 9024 27310 9036
rect 27617 9027 27675 9033
rect 27617 9024 27629 9027
rect 27304 8996 27629 9024
rect 27304 8984 27310 8996
rect 27617 8993 27629 8996
rect 27663 8993 27675 9027
rect 27617 8987 27675 8993
rect 27798 8984 27804 9036
rect 27856 8984 27862 9036
rect 27525 8959 27583 8965
rect 27525 8956 27537 8959
rect 24804 8928 24906 8956
rect 27080 8928 27537 8956
rect 24804 8925 24816 8928
rect 24758 8919 24816 8925
rect 22704 8860 23060 8888
rect 22704 8848 22710 8860
rect 24486 8820 24492 8832
rect 22572 8792 24492 8820
rect 24486 8780 24492 8792
rect 24544 8780 24550 8832
rect 24626 8820 24654 8919
rect 24872 8897 24900 8928
rect 27525 8925 27537 8928
rect 27571 8956 27583 8959
rect 27985 8959 28043 8965
rect 27985 8956 27997 8959
rect 27571 8928 27997 8956
rect 27571 8925 27583 8928
rect 27525 8919 27583 8925
rect 27985 8925 27997 8928
rect 28031 8925 28043 8959
rect 27985 8919 28043 8925
rect 28074 8916 28080 8968
rect 28132 8956 28138 8968
rect 28644 8965 28672 9064
rect 28718 9052 28724 9104
rect 28776 9092 28782 9104
rect 28813 9095 28871 9101
rect 28813 9092 28825 9095
rect 28776 9064 28825 9092
rect 28776 9052 28782 9064
rect 28813 9061 28825 9064
rect 28859 9092 28871 9095
rect 29549 9095 29607 9101
rect 29549 9092 29561 9095
rect 28859 9064 29561 9092
rect 28859 9061 28871 9064
rect 28813 9055 28871 9061
rect 29549 9061 29561 9064
rect 29595 9061 29607 9095
rect 29549 9055 29607 9061
rect 33042 8984 33048 9036
rect 33100 8984 33106 9036
rect 28353 8959 28411 8965
rect 28353 8956 28365 8959
rect 28132 8928 28365 8956
rect 28132 8916 28138 8928
rect 28353 8925 28365 8928
rect 28399 8956 28411 8959
rect 28629 8959 28687 8965
rect 28399 8928 28488 8956
rect 28399 8925 28411 8928
rect 28353 8919 28411 8925
rect 24857 8891 24915 8897
rect 24857 8857 24869 8891
rect 24903 8857 24915 8891
rect 24857 8851 24915 8857
rect 25041 8891 25099 8897
rect 25041 8857 25053 8891
rect 25087 8857 25099 8891
rect 25041 8851 25099 8857
rect 25952 8891 26010 8897
rect 25952 8857 25964 8891
rect 25998 8888 26010 8891
rect 25998 8860 27200 8888
rect 25998 8857 26010 8860
rect 25952 8851 26010 8857
rect 25056 8820 25084 8851
rect 27172 8829 27200 8860
rect 28166 8848 28172 8900
rect 28224 8848 28230 8900
rect 28261 8891 28319 8897
rect 28261 8857 28273 8891
rect 28307 8888 28319 8891
rect 28460 8888 28488 8928
rect 28629 8925 28641 8959
rect 28675 8925 28687 8959
rect 28629 8919 28687 8925
rect 32766 8916 32772 8968
rect 32824 8916 32830 8968
rect 28997 8891 29055 8897
rect 28997 8888 29009 8891
rect 28307 8860 28396 8888
rect 28460 8860 29009 8888
rect 28307 8857 28319 8860
rect 28261 8851 28319 8857
rect 28368 8832 28396 8860
rect 28997 8857 29009 8860
rect 29043 8888 29055 8891
rect 29181 8891 29239 8897
rect 29181 8888 29193 8891
rect 29043 8860 29193 8888
rect 29043 8857 29055 8860
rect 28997 8851 29055 8857
rect 29181 8857 29193 8860
rect 29227 8857 29239 8891
rect 29181 8851 29239 8857
rect 33134 8848 33140 8900
rect 33192 8888 33198 8900
rect 33192 8860 33534 8888
rect 33192 8848 33198 8860
rect 24626 8792 25084 8820
rect 27157 8823 27215 8829
rect 27157 8789 27169 8823
rect 27203 8789 27215 8823
rect 27157 8783 27215 8789
rect 28350 8780 28356 8832
rect 28408 8780 28414 8832
rect 1104 8730 35328 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35328 8730
rect 1104 8656 35328 8678
rect 4433 8619 4491 8625
rect 4433 8585 4445 8619
rect 4479 8616 4491 8619
rect 4614 8616 4620 8628
rect 4479 8588 4620 8616
rect 4479 8585 4491 8588
rect 4433 8579 4491 8585
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 9858 8576 9864 8628
rect 9916 8576 9922 8628
rect 10413 8619 10471 8625
rect 10413 8585 10425 8619
rect 10459 8616 10471 8619
rect 10686 8616 10692 8628
rect 10459 8588 10692 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 10870 8616 10876 8628
rect 10827 8588 10876 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 5994 8508 6000 8560
rect 6052 8548 6058 8560
rect 6457 8551 6515 8557
rect 6457 8548 6469 8551
rect 6052 8520 6469 8548
rect 6052 8508 6058 8520
rect 6457 8517 6469 8520
rect 6503 8548 6515 8551
rect 7469 8551 7527 8557
rect 7469 8548 7481 8551
rect 6503 8520 7481 8548
rect 6503 8517 6515 8520
rect 6457 8511 6515 8517
rect 7469 8517 7481 8520
rect 7515 8517 7527 8551
rect 9876 8548 9904 8576
rect 10045 8551 10103 8557
rect 10045 8548 10057 8551
rect 9876 8520 10057 8548
rect 7469 8511 7527 8517
rect 10045 8517 10057 8520
rect 10091 8548 10103 8551
rect 10505 8551 10563 8557
rect 10505 8548 10517 8551
rect 10091 8520 10517 8548
rect 10091 8517 10103 8520
rect 10045 8511 10103 8517
rect 10505 8517 10517 8520
rect 10551 8517 10563 8551
rect 10505 8511 10563 8517
rect 3878 8440 3884 8492
rect 3936 8480 3942 8492
rect 6914 8480 6920 8492
rect 3936 8452 6920 8480
rect 3936 8440 3942 8452
rect 6914 8440 6920 8452
rect 6972 8480 6978 8492
rect 7193 8483 7251 8489
rect 7193 8480 7205 8483
rect 6972 8452 7205 8480
rect 6972 8440 6978 8452
rect 7193 8449 7205 8452
rect 7239 8480 7251 8483
rect 8202 8480 8208 8492
rect 7239 8452 8208 8480
rect 7239 8449 7251 8452
rect 7193 8443 7251 8449
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 10134 8440 10140 8492
rect 10192 8440 10198 8492
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8480 10287 8483
rect 10796 8480 10824 8579
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 14366 8616 14372 8628
rect 11440 8588 14372 8616
rect 10275 8452 10824 8480
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 5258 8372 5264 8424
rect 5316 8412 5322 8424
rect 11330 8412 11336 8424
rect 5316 8384 11336 8412
rect 5316 8372 5322 8384
rect 11330 8372 11336 8384
rect 11388 8372 11394 8424
rect 3970 8304 3976 8356
rect 4028 8344 4034 8356
rect 11440 8344 11468 8588
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 14458 8576 14464 8628
rect 14516 8616 14522 8628
rect 15013 8619 15071 8625
rect 15013 8616 15025 8619
rect 14516 8588 15025 8616
rect 14516 8576 14522 8588
rect 15013 8585 15025 8588
rect 15059 8585 15071 8619
rect 15013 8579 15071 8585
rect 16485 8619 16543 8625
rect 16485 8585 16497 8619
rect 16531 8616 16543 8619
rect 17129 8619 17187 8625
rect 17129 8616 17141 8619
rect 16531 8588 17141 8616
rect 16531 8585 16543 8588
rect 16485 8579 16543 8585
rect 17129 8585 17141 8588
rect 17175 8616 17187 8619
rect 17402 8616 17408 8628
rect 17175 8588 17408 8616
rect 17175 8585 17187 8588
rect 17129 8579 17187 8585
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 17494 8576 17500 8628
rect 17552 8616 17558 8628
rect 17770 8616 17776 8628
rect 17552 8588 17776 8616
rect 17552 8576 17558 8588
rect 17770 8576 17776 8588
rect 17828 8576 17834 8628
rect 18969 8619 19027 8625
rect 18969 8616 18981 8619
rect 18248 8588 18981 8616
rect 15470 8548 15476 8560
rect 11808 8520 13124 8548
rect 11514 8372 11520 8424
rect 11572 8412 11578 8424
rect 11808 8421 11836 8520
rect 12060 8483 12118 8489
rect 12060 8449 12072 8483
rect 12106 8480 12118 8483
rect 12342 8480 12348 8492
rect 12106 8452 12348 8480
rect 12106 8449 12118 8452
rect 12060 8443 12118 8449
rect 12342 8440 12348 8452
rect 12400 8440 12406 8492
rect 11793 8415 11851 8421
rect 11793 8412 11805 8415
rect 11572 8384 11805 8412
rect 11572 8372 11578 8384
rect 11793 8381 11805 8384
rect 11839 8381 11851 8415
rect 13096 8412 13124 8520
rect 13832 8520 15056 8548
rect 13170 8440 13176 8492
rect 13228 8480 13234 8492
rect 13832 8480 13860 8520
rect 13228 8452 13860 8480
rect 13900 8483 13958 8489
rect 13228 8440 13234 8452
rect 13900 8449 13912 8483
rect 13946 8480 13958 8483
rect 14182 8480 14188 8492
rect 13946 8452 14188 8480
rect 13946 8449 13958 8452
rect 13900 8443 13958 8449
rect 14182 8440 14188 8452
rect 14240 8440 14246 8492
rect 13630 8412 13636 8424
rect 13096 8384 13636 8412
rect 11793 8375 11851 8381
rect 13630 8372 13636 8384
rect 13688 8372 13694 8424
rect 4028 8316 11468 8344
rect 15028 8344 15056 8520
rect 15120 8520 15476 8548
rect 15120 8489 15148 8520
rect 15470 8508 15476 8520
rect 15528 8508 15534 8560
rect 15562 8508 15568 8560
rect 15620 8548 15626 8560
rect 15620 8520 18184 8548
rect 15620 8508 15626 8520
rect 15105 8483 15163 8489
rect 15105 8449 15117 8483
rect 15151 8449 15163 8483
rect 15105 8443 15163 8449
rect 15372 8483 15430 8489
rect 15372 8449 15384 8483
rect 15418 8480 15430 8483
rect 15418 8452 16712 8480
rect 15418 8449 15430 8452
rect 15372 8443 15430 8449
rect 16684 8353 16712 8452
rect 16942 8440 16948 8492
rect 17000 8480 17006 8492
rect 17037 8483 17095 8489
rect 17037 8480 17049 8483
rect 17000 8452 17049 8480
rect 17000 8440 17006 8452
rect 17037 8449 17049 8452
rect 17083 8449 17095 8483
rect 17037 8443 17095 8449
rect 17865 8483 17923 8489
rect 17865 8449 17877 8483
rect 17911 8449 17923 8483
rect 17865 8443 17923 8449
rect 17221 8415 17279 8421
rect 17221 8412 17233 8415
rect 16776 8384 17233 8412
rect 16669 8347 16727 8353
rect 15028 8316 15148 8344
rect 4028 8304 4034 8316
rect 12802 8236 12808 8288
rect 12860 8276 12866 8288
rect 13173 8279 13231 8285
rect 13173 8276 13185 8279
rect 12860 8248 13185 8276
rect 12860 8236 12866 8248
rect 13173 8245 13185 8248
rect 13219 8245 13231 8279
rect 13173 8239 13231 8245
rect 14274 8236 14280 8288
rect 14332 8276 14338 8288
rect 14918 8276 14924 8288
rect 14332 8248 14924 8276
rect 14332 8236 14338 8248
rect 14918 8236 14924 8248
rect 14976 8236 14982 8288
rect 15120 8276 15148 8316
rect 16040 8316 16620 8344
rect 16040 8276 16068 8316
rect 15120 8248 16068 8276
rect 16592 8276 16620 8316
rect 16669 8313 16681 8347
rect 16715 8313 16727 8347
rect 16669 8307 16727 8313
rect 16776 8276 16804 8384
rect 17221 8381 17233 8384
rect 17267 8412 17279 8415
rect 17497 8415 17555 8421
rect 17497 8412 17509 8415
rect 17267 8384 17509 8412
rect 17267 8381 17279 8384
rect 17221 8375 17279 8381
rect 17497 8381 17509 8384
rect 17543 8381 17555 8415
rect 17880 8412 17908 8443
rect 18046 8440 18052 8492
rect 18104 8440 18110 8492
rect 18156 8489 18184 8520
rect 18248 8489 18276 8588
rect 18969 8585 18981 8588
rect 19015 8616 19027 8619
rect 19150 8616 19156 8628
rect 19015 8588 19156 8616
rect 19015 8585 19027 8588
rect 18969 8579 19027 8585
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 21085 8619 21143 8625
rect 19996 8588 20944 8616
rect 18785 8551 18843 8557
rect 18785 8517 18797 8551
rect 18831 8548 18843 8551
rect 19242 8548 19248 8560
rect 18831 8520 19248 8548
rect 18831 8517 18843 8520
rect 18785 8511 18843 8517
rect 18141 8483 18199 8489
rect 18141 8449 18153 8483
rect 18187 8449 18199 8483
rect 18141 8443 18199 8449
rect 18233 8483 18291 8489
rect 18233 8449 18245 8483
rect 18279 8449 18291 8483
rect 18233 8443 18291 8449
rect 18414 8440 18420 8492
rect 18472 8440 18478 8492
rect 18800 8412 18828 8511
rect 19242 8508 19248 8520
rect 19300 8508 19306 8560
rect 19886 8508 19892 8560
rect 19944 8548 19950 8560
rect 19996 8557 20024 8588
rect 19981 8551 20039 8557
rect 19981 8548 19993 8551
rect 19944 8520 19993 8548
rect 19944 8508 19950 8520
rect 19981 8517 19993 8520
rect 20027 8517 20039 8551
rect 19981 8511 20039 8517
rect 20806 8508 20812 8560
rect 20864 8508 20870 8560
rect 20916 8548 20944 8588
rect 21085 8585 21097 8619
rect 21131 8616 21143 8619
rect 21726 8616 21732 8628
rect 21131 8588 21732 8616
rect 21131 8585 21143 8588
rect 21085 8579 21143 8585
rect 21726 8576 21732 8588
rect 21784 8576 21790 8628
rect 21913 8619 21971 8625
rect 21913 8585 21925 8619
rect 21959 8616 21971 8619
rect 22094 8616 22100 8628
rect 21959 8588 22100 8616
rect 21959 8585 21971 8588
rect 21913 8579 21971 8585
rect 22094 8576 22100 8588
rect 22152 8576 22158 8628
rect 22738 8576 22744 8628
rect 22796 8576 22802 8628
rect 22830 8576 22836 8628
rect 22888 8576 22894 8628
rect 23106 8576 23112 8628
rect 23164 8576 23170 8628
rect 23382 8576 23388 8628
rect 23440 8616 23446 8628
rect 26786 8616 26792 8628
rect 23440 8588 26792 8616
rect 23440 8576 23446 8588
rect 26786 8576 26792 8588
rect 26844 8576 26850 8628
rect 28074 8616 28080 8628
rect 26896 8588 28080 8616
rect 21361 8551 21419 8557
rect 21361 8548 21373 8551
rect 20916 8520 21373 8548
rect 21361 8517 21373 8520
rect 21407 8517 21419 8551
rect 26896 8548 26924 8588
rect 28074 8576 28080 8588
rect 28132 8576 28138 8628
rect 28166 8576 28172 8628
rect 28224 8616 28230 8628
rect 28445 8619 28503 8625
rect 28445 8616 28457 8619
rect 28224 8588 28457 8616
rect 28224 8576 28230 8588
rect 28445 8585 28457 8588
rect 28491 8585 28503 8619
rect 28445 8579 28503 8585
rect 21361 8511 21419 8517
rect 22066 8520 26924 8548
rect 27240 8551 27298 8557
rect 20622 8489 20628 8492
rect 20441 8483 20499 8489
rect 20441 8449 20453 8483
rect 20487 8449 20499 8483
rect 20441 8443 20499 8449
rect 20589 8483 20628 8489
rect 20589 8449 20601 8483
rect 20589 8443 20628 8449
rect 19978 8412 19984 8424
rect 17880 8384 18828 8412
rect 19168 8384 19984 8412
rect 17497 8375 17555 8381
rect 17512 8344 17540 8375
rect 17512 8316 18557 8344
rect 16592 8248 16804 8276
rect 18529 8276 18557 8316
rect 18598 8304 18604 8356
rect 18656 8304 18662 8356
rect 19168 8344 19196 8384
rect 19978 8372 19984 8384
rect 20036 8372 20042 8424
rect 20456 8412 20484 8443
rect 20622 8440 20628 8443
rect 20680 8440 20686 8492
rect 20714 8440 20720 8492
rect 20772 8440 20778 8492
rect 20947 8483 21005 8489
rect 20947 8449 20959 8483
rect 20993 8480 21005 8483
rect 21542 8480 21548 8492
rect 20993 8452 21548 8480
rect 20993 8449 21005 8452
rect 20947 8443 21005 8449
rect 21542 8440 21548 8452
rect 21600 8440 21606 8492
rect 21910 8440 21916 8492
rect 21968 8480 21974 8492
rect 22066 8480 22094 8520
rect 27240 8517 27252 8551
rect 27286 8548 27298 8551
rect 27430 8548 27436 8560
rect 27286 8520 27436 8548
rect 27286 8517 27298 8520
rect 27240 8511 27298 8517
rect 27430 8508 27436 8520
rect 27488 8508 27494 8560
rect 27798 8508 27804 8560
rect 27856 8548 27862 8560
rect 28629 8551 28687 8557
rect 28629 8548 28641 8551
rect 27856 8520 28641 8548
rect 27856 8508 27862 8520
rect 28629 8517 28641 8520
rect 28675 8517 28687 8551
rect 28629 8511 28687 8517
rect 33134 8508 33140 8560
rect 33192 8508 33198 8560
rect 34790 8508 34796 8560
rect 34848 8508 34854 8560
rect 21968 8452 22094 8480
rect 21968 8440 21974 8452
rect 22554 8440 22560 8492
rect 22612 8480 22618 8492
rect 23017 8483 23075 8489
rect 23017 8480 23029 8483
rect 22612 8452 23029 8480
rect 22612 8440 22618 8452
rect 23017 8449 23029 8452
rect 23063 8480 23075 8483
rect 23106 8480 23112 8492
rect 23063 8452 23112 8480
rect 23063 8449 23075 8452
rect 23017 8443 23075 8449
rect 23106 8440 23112 8452
rect 23164 8440 23170 8492
rect 23201 8483 23259 8489
rect 23201 8449 23213 8483
rect 23247 8480 23259 8483
rect 23382 8480 23388 8492
rect 23247 8452 23388 8480
rect 23247 8449 23259 8452
rect 23201 8443 23259 8449
rect 23382 8440 23388 8452
rect 23440 8440 23446 8492
rect 23474 8440 23480 8492
rect 23532 8440 23538 8492
rect 26878 8440 26884 8492
rect 26936 8480 26942 8492
rect 26973 8483 27031 8489
rect 26973 8480 26985 8483
rect 26936 8452 26985 8480
rect 26936 8440 26942 8452
rect 26973 8449 26985 8452
rect 27019 8449 27031 8483
rect 30374 8480 30380 8492
rect 26973 8443 27031 8449
rect 27080 8452 30380 8480
rect 21082 8412 21088 8424
rect 20456 8384 21088 8412
rect 21082 8372 21088 8384
rect 21140 8372 21146 8424
rect 21174 8372 21180 8424
rect 21232 8412 21238 8424
rect 21637 8415 21695 8421
rect 21637 8412 21649 8415
rect 21232 8384 21649 8412
rect 21232 8372 21238 8384
rect 21637 8381 21649 8384
rect 21683 8381 21695 8415
rect 21637 8375 21695 8381
rect 22186 8372 22192 8424
rect 22244 8412 22250 8424
rect 22465 8415 22523 8421
rect 22465 8412 22477 8415
rect 22244 8384 22477 8412
rect 22244 8372 22250 8384
rect 22465 8381 22477 8384
rect 22511 8412 22523 8415
rect 22922 8412 22928 8424
rect 22511 8384 22928 8412
rect 22511 8381 22523 8384
rect 22465 8375 22523 8381
rect 22922 8372 22928 8384
rect 22980 8372 22986 8424
rect 27080 8412 27108 8452
rect 30374 8440 30380 8452
rect 30432 8440 30438 8492
rect 30653 8483 30711 8489
rect 30653 8449 30665 8483
rect 30699 8480 30711 8483
rect 31294 8480 31300 8492
rect 30699 8452 31300 8480
rect 30699 8449 30711 8452
rect 30653 8443 30711 8449
rect 31294 8440 31300 8452
rect 31352 8440 31358 8492
rect 34238 8440 34244 8492
rect 34296 8480 34302 8492
rect 34517 8483 34575 8489
rect 34517 8480 34529 8483
rect 34296 8452 34529 8480
rect 34296 8440 34302 8452
rect 34517 8449 34529 8452
rect 34563 8449 34575 8483
rect 34517 8443 34575 8449
rect 29638 8412 29644 8424
rect 23676 8384 27108 8412
rect 28000 8384 29644 8412
rect 18708 8316 19196 8344
rect 18708 8276 18736 8316
rect 19242 8304 19248 8356
rect 19300 8344 19306 8356
rect 21542 8344 21548 8356
rect 19300 8316 21548 8344
rect 19300 8304 19306 8316
rect 21542 8304 21548 8316
rect 21600 8304 21606 8356
rect 21910 8304 21916 8356
rect 21968 8344 21974 8356
rect 22097 8347 22155 8353
rect 22097 8344 22109 8347
rect 21968 8316 22109 8344
rect 21968 8304 21974 8316
rect 22097 8313 22109 8316
rect 22143 8344 22155 8347
rect 23676 8344 23704 8384
rect 22143 8316 23704 8344
rect 22143 8313 22155 8316
rect 22097 8307 22155 8313
rect 23750 8304 23756 8356
rect 23808 8344 23814 8356
rect 28000 8344 28028 8384
rect 29638 8372 29644 8384
rect 29696 8372 29702 8424
rect 30745 8415 30803 8421
rect 30745 8381 30757 8415
rect 30791 8412 30803 8415
rect 31110 8412 31116 8424
rect 30791 8384 31116 8412
rect 30791 8381 30803 8384
rect 30745 8375 30803 8381
rect 31110 8372 31116 8384
rect 31168 8372 31174 8424
rect 32125 8415 32183 8421
rect 32125 8381 32137 8415
rect 32171 8381 32183 8415
rect 32125 8375 32183 8381
rect 23808 8316 27016 8344
rect 23808 8304 23814 8316
rect 18529 8248 18736 8276
rect 19610 8236 19616 8288
rect 19668 8276 19674 8288
rect 20073 8279 20131 8285
rect 20073 8276 20085 8279
rect 19668 8248 20085 8276
rect 19668 8236 19674 8248
rect 20073 8245 20085 8248
rect 20119 8276 20131 8279
rect 21177 8279 21235 8285
rect 21177 8276 21189 8279
rect 20119 8248 21189 8276
rect 20119 8245 20131 8248
rect 20073 8239 20131 8245
rect 21177 8245 21189 8248
rect 21223 8276 21235 8279
rect 21358 8276 21364 8288
rect 21223 8248 21364 8276
rect 21223 8245 21235 8248
rect 21177 8239 21235 8245
rect 21358 8236 21364 8248
rect 21416 8236 21422 8288
rect 23290 8236 23296 8288
rect 23348 8236 23354 8288
rect 23382 8236 23388 8288
rect 23440 8276 23446 8288
rect 25130 8276 25136 8288
rect 23440 8248 25136 8276
rect 23440 8236 23446 8248
rect 25130 8236 25136 8248
rect 25188 8236 25194 8288
rect 26988 8276 27016 8316
rect 27908 8316 28028 8344
rect 27908 8276 27936 8316
rect 28350 8304 28356 8356
rect 28408 8304 28414 8356
rect 26988 8248 27936 8276
rect 29822 8236 29828 8288
rect 29880 8276 29886 8288
rect 30285 8279 30343 8285
rect 30285 8276 30297 8279
rect 29880 8248 30297 8276
rect 29880 8236 29886 8248
rect 30285 8245 30297 8248
rect 30331 8245 30343 8279
rect 32140 8276 32168 8375
rect 32398 8372 32404 8424
rect 32456 8372 32462 8424
rect 32490 8372 32496 8424
rect 32548 8412 32554 8424
rect 33873 8415 33931 8421
rect 33873 8412 33885 8415
rect 32548 8384 33885 8412
rect 32548 8372 32554 8384
rect 33873 8381 33885 8384
rect 33919 8381 33931 8415
rect 33873 8375 33931 8381
rect 32766 8276 32772 8288
rect 32140 8248 32772 8276
rect 30285 8239 30343 8245
rect 32766 8236 32772 8248
rect 32824 8236 32830 8288
rect 1104 8186 35328 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 35328 8186
rect 1104 8112 35328 8134
rect 9861 8075 9919 8081
rect 9861 8041 9873 8075
rect 9907 8072 9919 8075
rect 13538 8072 13544 8084
rect 9907 8044 13544 8072
rect 9907 8041 9919 8044
rect 9861 8035 9919 8041
rect 7742 7896 7748 7948
rect 7800 7896 7806 7948
rect 7929 7939 7987 7945
rect 7929 7905 7941 7939
rect 7975 7936 7987 7939
rect 9585 7939 9643 7945
rect 7975 7908 8248 7936
rect 7975 7905 7987 7908
rect 7929 7899 7987 7905
rect 6914 7828 6920 7880
rect 6972 7828 6978 7880
rect 7653 7871 7711 7877
rect 7653 7837 7665 7871
rect 7699 7868 7711 7871
rect 8018 7868 8024 7880
rect 7699 7840 8024 7868
rect 7699 7837 7711 7840
rect 7653 7831 7711 7837
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 8220 7809 8248 7908
rect 9585 7905 9597 7939
rect 9631 7936 9643 7939
rect 9876 7936 9904 8035
rect 13538 8032 13544 8044
rect 13596 8072 13602 8084
rect 17957 8075 18015 8081
rect 13596 8044 17908 8072
rect 13596 8032 13602 8044
rect 12342 7964 12348 8016
rect 12400 7964 12406 8016
rect 17880 8004 17908 8044
rect 17957 8041 17969 8075
rect 18003 8072 18015 8075
rect 18046 8072 18052 8084
rect 18003 8044 18052 8072
rect 18003 8041 18015 8044
rect 17957 8035 18015 8041
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 19978 8032 19984 8084
rect 20036 8032 20042 8084
rect 20254 8032 20260 8084
rect 20312 8072 20318 8084
rect 20312 8044 22094 8072
rect 20312 8032 20318 8044
rect 19610 8004 19616 8016
rect 17880 7976 19616 8004
rect 19610 7964 19616 7976
rect 19668 7964 19674 8016
rect 19702 7964 19708 8016
rect 19760 8004 19766 8016
rect 19760 7976 21404 8004
rect 19760 7964 19766 7976
rect 9631 7908 9904 7936
rect 9631 7905 9643 7908
rect 9585 7899 9643 7905
rect 12802 7896 12808 7948
rect 12860 7896 12866 7948
rect 12989 7939 13047 7945
rect 12989 7905 13001 7939
rect 13035 7936 13047 7939
rect 13446 7936 13452 7948
rect 13035 7908 13452 7936
rect 13035 7905 13047 7908
rect 12989 7899 13047 7905
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 15102 7936 15108 7948
rect 13556 7908 15108 7936
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7868 9367 7871
rect 9858 7868 9864 7880
rect 9355 7840 9864 7868
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 8205 7803 8263 7809
rect 8205 7769 8217 7803
rect 8251 7800 8263 7803
rect 13556 7800 13584 7908
rect 15102 7896 15108 7908
rect 15160 7896 15166 7948
rect 17129 7939 17187 7945
rect 17129 7936 17141 7939
rect 15212 7908 17141 7936
rect 13630 7828 13636 7880
rect 13688 7868 13694 7880
rect 13725 7871 13783 7877
rect 13725 7868 13737 7871
rect 13688 7840 13737 7868
rect 13688 7828 13694 7840
rect 13725 7837 13737 7840
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 8251 7772 13584 7800
rect 13740 7800 13768 7831
rect 13998 7828 14004 7880
rect 14056 7868 14062 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 14056 7840 14105 7868
rect 14056 7828 14062 7840
rect 14093 7837 14105 7840
rect 14139 7868 14151 7871
rect 14734 7868 14740 7880
rect 14139 7840 14740 7868
rect 14139 7837 14151 7840
rect 14093 7831 14151 7837
rect 14734 7828 14740 7840
rect 14792 7828 14798 7880
rect 15010 7828 15016 7880
rect 15068 7868 15074 7880
rect 15212 7868 15240 7908
rect 17129 7905 17141 7908
rect 17175 7936 17187 7939
rect 17494 7936 17500 7948
rect 17175 7908 17500 7936
rect 17175 7905 17187 7908
rect 17129 7899 17187 7905
rect 17494 7896 17500 7908
rect 17552 7896 17558 7948
rect 17678 7896 17684 7948
rect 17736 7936 17742 7948
rect 18049 7939 18107 7945
rect 18049 7936 18061 7939
rect 17736 7908 18061 7936
rect 17736 7896 17742 7908
rect 18049 7905 18061 7908
rect 18095 7936 18107 7939
rect 18095 7908 19932 7936
rect 18095 7905 18107 7908
rect 18049 7899 18107 7905
rect 15068 7840 15240 7868
rect 16853 7871 16911 7877
rect 15068 7828 15074 7840
rect 16853 7837 16865 7871
rect 16899 7868 16911 7871
rect 16942 7868 16948 7880
rect 16899 7840 16948 7868
rect 16899 7837 16911 7840
rect 16853 7831 16911 7837
rect 16942 7828 16948 7840
rect 17000 7828 17006 7880
rect 17310 7828 17316 7880
rect 17368 7828 17374 7880
rect 17402 7828 17408 7880
rect 17460 7868 17466 7880
rect 17862 7877 17868 7880
rect 17819 7871 17868 7877
rect 17460 7840 17505 7868
rect 17460 7828 17466 7840
rect 17819 7837 17831 7871
rect 17865 7837 17868 7871
rect 17819 7831 17868 7837
rect 17862 7828 17868 7831
rect 17920 7868 17926 7880
rect 18233 7871 18291 7877
rect 18233 7868 18245 7871
rect 17920 7840 18245 7868
rect 17920 7828 17926 7840
rect 18233 7837 18245 7840
rect 18279 7837 18291 7871
rect 18233 7831 18291 7837
rect 14921 7803 14979 7809
rect 14921 7800 14933 7803
rect 13740 7772 14933 7800
rect 8251 7769 8263 7772
rect 8205 7763 8263 7769
rect 14921 7769 14933 7772
rect 14967 7800 14979 7803
rect 15930 7800 15936 7812
rect 14967 7772 15936 7800
rect 14967 7769 14979 7772
rect 14921 7763 14979 7769
rect 15930 7760 15936 7772
rect 15988 7760 15994 7812
rect 17586 7760 17592 7812
rect 17644 7760 17650 7812
rect 17681 7803 17739 7809
rect 17681 7769 17693 7803
rect 17727 7769 17739 7803
rect 19904 7800 19932 7908
rect 19978 7896 19984 7948
rect 20036 7936 20042 7948
rect 20438 7936 20444 7948
rect 20036 7908 20444 7936
rect 20036 7896 20042 7908
rect 20438 7896 20444 7908
rect 20496 7936 20502 7948
rect 20625 7939 20683 7945
rect 20625 7936 20637 7939
rect 20496 7908 20637 7936
rect 20496 7896 20502 7908
rect 20625 7905 20637 7908
rect 20671 7905 20683 7939
rect 20625 7899 20683 7905
rect 21266 7896 21272 7948
rect 21324 7896 21330 7948
rect 21376 7945 21404 7976
rect 21910 7964 21916 8016
rect 21968 7964 21974 8016
rect 22066 8004 22094 8044
rect 22186 8032 22192 8084
rect 22244 8032 22250 8084
rect 22922 8032 22928 8084
rect 22980 8072 22986 8084
rect 23290 8072 23296 8084
rect 22980 8044 23296 8072
rect 22980 8032 22986 8044
rect 23290 8032 23296 8044
rect 23348 8072 23354 8084
rect 23477 8075 23535 8081
rect 23477 8072 23489 8075
rect 23348 8044 23489 8072
rect 23348 8032 23354 8044
rect 23477 8041 23489 8044
rect 23523 8041 23535 8075
rect 23477 8035 23535 8041
rect 27065 8075 27123 8081
rect 27065 8041 27077 8075
rect 27111 8072 27123 8075
rect 27430 8072 27436 8084
rect 27111 8044 27436 8072
rect 27111 8041 27123 8044
rect 27065 8035 27123 8041
rect 27430 8032 27436 8044
rect 27488 8032 27494 8084
rect 27985 8075 28043 8081
rect 27985 8041 27997 8075
rect 28031 8072 28043 8075
rect 28718 8072 28724 8084
rect 28031 8044 28724 8072
rect 28031 8041 28043 8044
rect 27985 8035 28043 8041
rect 23017 8007 23075 8013
rect 23017 8004 23029 8007
rect 22066 7976 23029 8004
rect 23017 7973 23029 7976
rect 23063 8004 23075 8007
rect 23937 8007 23995 8013
rect 23937 8004 23949 8007
rect 23063 7976 23949 8004
rect 23063 7973 23075 7976
rect 23017 7967 23075 7973
rect 23937 7973 23949 7976
rect 23983 7973 23995 8007
rect 23937 7967 23995 7973
rect 21361 7939 21419 7945
rect 21361 7905 21373 7939
rect 21407 7905 21419 7939
rect 21361 7899 21419 7905
rect 20165 7871 20223 7877
rect 20165 7837 20177 7871
rect 20211 7868 20223 7871
rect 20254 7868 20260 7880
rect 20211 7840 20260 7868
rect 20211 7837 20223 7840
rect 20165 7831 20223 7837
rect 20254 7828 20260 7840
rect 20312 7828 20318 7880
rect 20346 7828 20352 7880
rect 20404 7868 20410 7880
rect 21177 7871 21235 7877
rect 21177 7868 21189 7871
rect 20404 7840 21189 7868
rect 20404 7828 20410 7840
rect 21177 7837 21189 7840
rect 21223 7837 21235 7871
rect 21177 7831 21235 7837
rect 20714 7800 20720 7812
rect 19904 7772 20720 7800
rect 17681 7763 17739 7769
rect 7282 7692 7288 7744
rect 7340 7692 7346 7744
rect 8938 7692 8944 7744
rect 8996 7692 9002 7744
rect 9401 7735 9459 7741
rect 9401 7701 9413 7735
rect 9447 7732 9459 7735
rect 9582 7732 9588 7744
rect 9447 7704 9588 7732
rect 9447 7701 9459 7704
rect 9401 7695 9459 7701
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 12713 7735 12771 7741
rect 12713 7701 12725 7735
rect 12759 7732 12771 7735
rect 13814 7732 13820 7744
rect 12759 7704 13820 7732
rect 12759 7701 12771 7704
rect 12713 7695 12771 7701
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 16482 7692 16488 7744
rect 16540 7692 16546 7744
rect 16945 7735 17003 7741
rect 16945 7701 16957 7735
rect 16991 7732 17003 7735
rect 17310 7732 17316 7744
rect 16991 7704 17316 7732
rect 16991 7701 17003 7704
rect 16945 7695 17003 7701
rect 17310 7692 17316 7704
rect 17368 7732 17374 7744
rect 17696 7732 17724 7763
rect 20714 7760 20720 7772
rect 20772 7760 20778 7812
rect 17368 7704 17724 7732
rect 17368 7692 17374 7704
rect 19610 7692 19616 7744
rect 19668 7732 19674 7744
rect 20441 7735 20499 7741
rect 20441 7732 20453 7735
rect 19668 7704 20453 7732
rect 19668 7692 19674 7704
rect 20441 7701 20453 7704
rect 20487 7701 20499 7735
rect 20441 7695 20499 7701
rect 20806 7692 20812 7744
rect 20864 7692 20870 7744
rect 21376 7732 21404 7899
rect 21928 7868 21956 7964
rect 27709 7939 27767 7945
rect 27709 7905 27721 7939
rect 27755 7936 27767 7939
rect 28000 7936 28028 8035
rect 28718 8032 28724 8044
rect 28776 8032 28782 8084
rect 31294 8032 31300 8084
rect 31352 8032 31358 8084
rect 32398 8032 32404 8084
rect 32456 8072 32462 8084
rect 32585 8075 32643 8081
rect 32585 8072 32597 8075
rect 32456 8044 32597 8072
rect 32456 8032 32462 8044
rect 32585 8041 32597 8044
rect 32631 8041 32643 8075
rect 32585 8035 32643 8041
rect 27755 7908 28028 7936
rect 29549 7939 29607 7945
rect 27755 7905 27767 7908
rect 27709 7899 27767 7905
rect 29549 7905 29561 7939
rect 29595 7936 29607 7939
rect 29914 7936 29920 7948
rect 29595 7908 29920 7936
rect 29595 7905 29607 7908
rect 29549 7899 29607 7905
rect 29914 7896 29920 7908
rect 29972 7896 29978 7948
rect 31018 7896 31024 7948
rect 31076 7896 31082 7948
rect 31110 7896 31116 7948
rect 31168 7936 31174 7948
rect 31941 7939 31999 7945
rect 31941 7936 31953 7939
rect 31168 7908 31953 7936
rect 31168 7896 31174 7908
rect 31941 7905 31953 7908
rect 31987 7905 31999 7939
rect 33134 7936 33140 7948
rect 31941 7899 31999 7905
rect 32140 7908 33140 7936
rect 22005 7871 22063 7877
rect 22005 7868 22017 7871
rect 21928 7840 22017 7868
rect 22005 7837 22017 7840
rect 22051 7837 22063 7871
rect 22005 7831 22063 7837
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7868 22891 7871
rect 22922 7868 22928 7880
rect 22879 7840 22928 7868
rect 22879 7837 22891 7840
rect 22833 7831 22891 7837
rect 22922 7828 22928 7840
rect 22980 7828 22986 7880
rect 23014 7828 23020 7880
rect 23072 7828 23078 7880
rect 23109 7871 23167 7877
rect 23109 7837 23121 7871
rect 23155 7868 23167 7871
rect 23477 7871 23535 7877
rect 23477 7868 23489 7871
rect 23155 7840 23489 7868
rect 23155 7837 23167 7840
rect 23109 7831 23167 7837
rect 23477 7837 23489 7840
rect 23523 7868 23535 7871
rect 23750 7868 23756 7880
rect 23523 7840 23756 7868
rect 23523 7837 23535 7840
rect 23477 7831 23535 7837
rect 23750 7828 23756 7840
rect 23808 7828 23814 7880
rect 23842 7828 23848 7880
rect 23900 7828 23906 7880
rect 27246 7828 27252 7880
rect 27304 7868 27310 7880
rect 27433 7871 27491 7877
rect 27433 7868 27445 7871
rect 27304 7840 27445 7868
rect 27304 7828 27310 7840
rect 27433 7837 27445 7840
rect 27479 7837 27491 7871
rect 27433 7831 27491 7837
rect 27525 7871 27583 7877
rect 27525 7837 27537 7871
rect 27571 7868 27583 7871
rect 28350 7868 28356 7880
rect 27571 7840 28356 7868
rect 27571 7837 27583 7840
rect 27525 7831 27583 7837
rect 28350 7828 28356 7840
rect 28408 7828 28414 7880
rect 31036 7868 31064 7896
rect 32140 7868 32168 7908
rect 33134 7896 33140 7908
rect 33192 7896 33198 7948
rect 30958 7840 32168 7868
rect 32217 7871 32275 7877
rect 32217 7837 32229 7871
rect 32263 7868 32275 7871
rect 32490 7868 32496 7880
rect 32263 7840 32496 7868
rect 32263 7837 32275 7840
rect 32217 7831 32275 7837
rect 32490 7828 32496 7840
rect 32548 7828 32554 7880
rect 34330 7828 34336 7880
rect 34388 7868 34394 7880
rect 34517 7871 34575 7877
rect 34517 7868 34529 7871
rect 34388 7840 34529 7868
rect 34388 7828 34394 7840
rect 34517 7837 34529 7840
rect 34563 7837 34575 7871
rect 34517 7831 34575 7837
rect 21729 7803 21787 7809
rect 21729 7769 21741 7803
rect 21775 7800 21787 7803
rect 21775 7772 22416 7800
rect 21775 7769 21787 7772
rect 21729 7763 21787 7769
rect 21818 7732 21824 7744
rect 21376 7704 21824 7732
rect 21818 7692 21824 7704
rect 21876 7732 21882 7744
rect 22186 7732 22192 7744
rect 21876 7704 22192 7732
rect 21876 7692 21882 7704
rect 22186 7692 22192 7704
rect 22244 7692 22250 7744
rect 22388 7732 22416 7772
rect 22462 7760 22468 7812
rect 22520 7800 22526 7812
rect 22520 7772 28994 7800
rect 22520 7760 22526 7772
rect 23293 7735 23351 7741
rect 23293 7732 23305 7735
rect 22388 7704 23305 7732
rect 23293 7701 23305 7704
rect 23339 7701 23351 7735
rect 23293 7695 23351 7701
rect 23382 7692 23388 7744
rect 23440 7732 23446 7744
rect 27154 7732 27160 7744
rect 23440 7704 27160 7732
rect 23440 7692 23446 7704
rect 27154 7692 27160 7704
rect 27212 7692 27218 7744
rect 28966 7732 28994 7772
rect 29822 7760 29828 7812
rect 29880 7760 29886 7812
rect 32582 7800 32588 7812
rect 31128 7772 32588 7800
rect 31128 7732 31156 7772
rect 32582 7760 32588 7772
rect 32640 7800 32646 7812
rect 32861 7803 32919 7809
rect 32861 7800 32873 7803
rect 32640 7772 32873 7800
rect 32640 7760 32646 7772
rect 32861 7769 32873 7772
rect 32907 7769 32919 7803
rect 32861 7763 32919 7769
rect 34241 7803 34299 7809
rect 34241 7769 34253 7803
rect 34287 7800 34299 7803
rect 34698 7800 34704 7812
rect 34287 7772 34704 7800
rect 34287 7769 34299 7772
rect 34241 7763 34299 7769
rect 34698 7760 34704 7772
rect 34756 7760 34762 7812
rect 28966 7704 31156 7732
rect 31570 7692 31576 7744
rect 31628 7732 31634 7744
rect 32125 7735 32183 7741
rect 32125 7732 32137 7735
rect 31628 7704 32137 7732
rect 31628 7692 31634 7704
rect 32125 7701 32137 7704
rect 32171 7701 32183 7735
rect 32125 7695 32183 7701
rect 32674 7692 32680 7744
rect 32732 7692 32738 7744
rect 33042 7692 33048 7744
rect 33100 7732 33106 7744
rect 33229 7735 33287 7741
rect 33229 7732 33241 7735
rect 33100 7704 33241 7732
rect 33100 7692 33106 7704
rect 33229 7701 33241 7704
rect 33275 7701 33287 7735
rect 33229 7695 33287 7701
rect 1104 7642 35328 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35328 7642
rect 1104 7568 35328 7590
rect 7837 7531 7895 7537
rect 7837 7497 7849 7531
rect 7883 7528 7895 7531
rect 8018 7528 8024 7540
rect 7883 7500 8024 7528
rect 7883 7497 7895 7500
rect 7837 7491 7895 7497
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 9309 7531 9367 7537
rect 9309 7497 9321 7531
rect 9355 7528 9367 7531
rect 9858 7528 9864 7540
rect 9355 7500 9864 7528
rect 9355 7497 9367 7500
rect 9309 7491 9367 7497
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 10134 7488 10140 7540
rect 10192 7528 10198 7540
rect 10781 7531 10839 7537
rect 10781 7528 10793 7531
rect 10192 7500 10793 7528
rect 10192 7488 10198 7500
rect 10781 7497 10793 7500
rect 10827 7497 10839 7531
rect 10781 7491 10839 7497
rect 12710 7488 12716 7540
rect 12768 7528 12774 7540
rect 12897 7531 12955 7537
rect 12897 7528 12909 7531
rect 12768 7500 12909 7528
rect 12768 7488 12774 7500
rect 12897 7497 12909 7500
rect 12943 7497 12955 7531
rect 12897 7491 12955 7497
rect 13265 7531 13323 7537
rect 13265 7497 13277 7531
rect 13311 7528 13323 7531
rect 13446 7528 13452 7540
rect 13311 7500 13452 7528
rect 13311 7497 13323 7500
rect 13265 7491 13323 7497
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 13998 7488 14004 7540
rect 14056 7488 14062 7540
rect 14182 7488 14188 7540
rect 14240 7488 14246 7540
rect 14458 7488 14464 7540
rect 14516 7528 14522 7540
rect 14553 7531 14611 7537
rect 14553 7528 14565 7531
rect 14516 7500 14565 7528
rect 14516 7488 14522 7500
rect 14553 7497 14565 7500
rect 14599 7497 14611 7531
rect 14553 7491 14611 7497
rect 15102 7488 15108 7540
rect 15160 7488 15166 7540
rect 18414 7488 18420 7540
rect 18472 7528 18478 7540
rect 18785 7531 18843 7537
rect 18785 7528 18797 7531
rect 18472 7500 18797 7528
rect 18472 7488 18478 7500
rect 18785 7497 18797 7500
rect 18831 7497 18843 7531
rect 18785 7491 18843 7497
rect 20349 7531 20407 7537
rect 20349 7497 20361 7531
rect 20395 7497 20407 7531
rect 20349 7491 20407 7497
rect 6914 7460 6920 7472
rect 6472 7432 6920 7460
rect 1302 7352 1308 7404
rect 1360 7392 1366 7404
rect 6472 7401 6500 7432
rect 6914 7420 6920 7432
rect 6972 7460 6978 7472
rect 6972 7432 9444 7460
rect 6972 7420 6978 7432
rect 1489 7395 1547 7401
rect 1489 7392 1501 7395
rect 1360 7364 1501 7392
rect 1360 7352 1366 7364
rect 1489 7361 1501 7364
rect 1535 7392 1547 7395
rect 1949 7395 2007 7401
rect 1949 7392 1961 7395
rect 1535 7364 1961 7392
rect 1535 7361 1547 7364
rect 1489 7355 1547 7361
rect 1949 7361 1961 7364
rect 1995 7361 2007 7395
rect 1949 7355 2007 7361
rect 6457 7395 6515 7401
rect 6457 7361 6469 7395
rect 6503 7361 6515 7395
rect 6457 7355 6515 7361
rect 6724 7395 6782 7401
rect 6724 7361 6736 7395
rect 6770 7392 6782 7395
rect 7282 7392 7288 7404
rect 6770 7364 7288 7392
rect 6770 7361 6782 7364
rect 6724 7355 6782 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7944 7401 7972 7432
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 8196 7395 8254 7401
rect 8196 7361 8208 7395
rect 8242 7392 8254 7395
rect 8938 7392 8944 7404
rect 8242 7364 8944 7392
rect 8242 7361 8254 7364
rect 8196 7355 8254 7361
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 9416 7401 9444 7432
rect 13814 7420 13820 7472
rect 13872 7460 13878 7472
rect 14645 7463 14703 7469
rect 14645 7460 14657 7463
rect 13872 7432 14657 7460
rect 13872 7420 13878 7432
rect 14568 7404 14596 7432
rect 14645 7429 14657 7432
rect 14691 7429 14703 7463
rect 14645 7423 14703 7429
rect 19144 7463 19202 7469
rect 19144 7429 19156 7463
rect 19190 7460 19202 7463
rect 20364 7460 20392 7491
rect 20622 7488 20628 7540
rect 20680 7528 20686 7540
rect 20809 7531 20867 7537
rect 20809 7528 20821 7531
rect 20680 7500 20821 7528
rect 20680 7488 20686 7500
rect 20809 7497 20821 7500
rect 20855 7497 20867 7531
rect 20809 7491 20867 7497
rect 21818 7488 21824 7540
rect 21876 7488 21882 7540
rect 21910 7488 21916 7540
rect 21968 7528 21974 7540
rect 22005 7531 22063 7537
rect 22005 7528 22017 7531
rect 21968 7500 22017 7528
rect 21968 7488 21974 7500
rect 22005 7497 22017 7500
rect 22051 7497 22063 7531
rect 22005 7491 22063 7497
rect 22465 7531 22523 7537
rect 22465 7497 22477 7531
rect 22511 7528 22523 7531
rect 22738 7528 22744 7540
rect 22511 7500 22744 7528
rect 22511 7497 22523 7500
rect 22465 7491 22523 7497
rect 22738 7488 22744 7500
rect 22796 7488 22802 7540
rect 22922 7488 22928 7540
rect 22980 7488 22986 7540
rect 23109 7531 23167 7537
rect 23109 7497 23121 7531
rect 23155 7528 23167 7531
rect 23382 7528 23388 7540
rect 23155 7500 23388 7528
rect 23155 7497 23167 7500
rect 23109 7491 23167 7497
rect 23382 7488 23388 7500
rect 23440 7488 23446 7540
rect 23569 7531 23627 7537
rect 23569 7497 23581 7531
rect 23615 7528 23627 7531
rect 23658 7528 23664 7540
rect 23615 7500 23664 7528
rect 23615 7497 23627 7500
rect 23569 7491 23627 7497
rect 23658 7488 23664 7500
rect 23716 7488 23722 7540
rect 23753 7531 23811 7537
rect 23753 7497 23765 7531
rect 23799 7528 23811 7531
rect 23842 7528 23848 7540
rect 23799 7500 23848 7528
rect 23799 7497 23811 7500
rect 23753 7491 23811 7497
rect 22940 7460 22968 7488
rect 19190 7432 20392 7460
rect 22756 7432 22968 7460
rect 19190 7429 19202 7432
rect 19144 7423 19202 7429
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7361 9459 7395
rect 9401 7355 9459 7361
rect 9668 7395 9726 7401
rect 9668 7361 9680 7395
rect 9714 7392 9726 7395
rect 10042 7392 10048 7404
rect 9714 7364 10048 7392
rect 9714 7361 9726 7364
rect 9668 7355 9726 7361
rect 10042 7352 10048 7364
rect 10100 7352 10106 7404
rect 11514 7352 11520 7404
rect 11572 7352 11578 7404
rect 11606 7352 11612 7404
rect 11664 7392 11670 7404
rect 11773 7395 11831 7401
rect 11773 7392 11785 7395
rect 11664 7364 11785 7392
rect 11664 7352 11670 7364
rect 11773 7361 11785 7364
rect 11819 7361 11831 7395
rect 11773 7355 11831 7361
rect 14550 7352 14556 7404
rect 14608 7352 14614 7404
rect 17678 7401 17684 7404
rect 17672 7355 17684 7401
rect 17678 7352 17684 7355
rect 17736 7352 17742 7404
rect 18874 7352 18880 7404
rect 18932 7352 18938 7404
rect 20346 7352 20352 7404
rect 20404 7392 20410 7404
rect 20717 7395 20775 7401
rect 20717 7392 20729 7395
rect 20404 7364 20729 7392
rect 20404 7352 20410 7364
rect 20717 7361 20729 7364
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 21542 7352 21548 7404
rect 21600 7392 21606 7404
rect 22756 7401 22784 7432
rect 23014 7420 23020 7472
rect 23072 7460 23078 7472
rect 23768 7460 23796 7491
rect 23842 7488 23848 7500
rect 23900 7488 23906 7540
rect 24762 7488 24768 7540
rect 24820 7528 24826 7540
rect 24820 7500 25636 7528
rect 24820 7488 24826 7500
rect 23072 7432 23796 7460
rect 24121 7463 24179 7469
rect 23072 7420 23078 7432
rect 22373 7395 22431 7401
rect 22373 7392 22385 7395
rect 21600 7364 22385 7392
rect 21600 7352 21606 7364
rect 22373 7361 22385 7364
rect 22419 7361 22431 7395
rect 22373 7355 22431 7361
rect 22741 7395 22799 7401
rect 22741 7361 22753 7395
rect 22787 7361 22799 7395
rect 22741 7355 22799 7361
rect 22833 7395 22891 7401
rect 22833 7361 22845 7395
rect 22879 7361 22891 7395
rect 22833 7355 22891 7361
rect 22925 7395 22983 7401
rect 22925 7361 22937 7395
rect 22971 7392 22983 7395
rect 23032 7392 23060 7420
rect 22971 7364 23060 7392
rect 22971 7361 22983 7364
rect 22925 7355 22983 7361
rect 14829 7327 14887 7333
rect 14829 7293 14841 7327
rect 14875 7324 14887 7327
rect 15102 7324 15108 7336
rect 14875 7296 15108 7324
rect 14875 7293 14887 7296
rect 14829 7287 14887 7293
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 15930 7284 15936 7336
rect 15988 7324 15994 7336
rect 17405 7327 17463 7333
rect 17405 7324 17417 7327
rect 15988 7296 17417 7324
rect 15988 7284 15994 7296
rect 17405 7293 17417 7296
rect 17451 7293 17463 7327
rect 17405 7287 17463 7293
rect 20438 7284 20444 7336
rect 20496 7324 20502 7336
rect 20901 7327 20959 7333
rect 20901 7324 20913 7327
rect 20496 7296 20913 7324
rect 20496 7284 20502 7296
rect 20901 7293 20913 7296
rect 20947 7293 20959 7327
rect 20901 7287 20959 7293
rect 22646 7284 22652 7336
rect 22704 7324 22710 7336
rect 22848 7324 22876 7355
rect 23106 7352 23112 7404
rect 23164 7392 23170 7404
rect 23309 7401 23337 7432
rect 24121 7429 24133 7463
rect 24167 7460 24179 7463
rect 25222 7460 25228 7472
rect 24167 7432 25228 7460
rect 24167 7429 24179 7432
rect 24121 7423 24179 7429
rect 23201 7395 23259 7401
rect 23201 7392 23213 7395
rect 23164 7364 23213 7392
rect 23164 7352 23170 7364
rect 23201 7361 23213 7364
rect 23247 7361 23259 7395
rect 23201 7355 23259 7361
rect 23294 7395 23352 7401
rect 23294 7361 23306 7395
rect 23340 7361 23352 7395
rect 23294 7355 23352 7361
rect 23912 7395 23970 7401
rect 23912 7361 23924 7395
rect 23958 7392 23970 7395
rect 24302 7392 24308 7404
rect 23958 7364 24308 7392
rect 23958 7361 23970 7364
rect 23912 7355 23970 7361
rect 24302 7352 24308 7364
rect 24360 7352 24366 7404
rect 24486 7352 24492 7404
rect 24544 7352 24550 7404
rect 24762 7352 24768 7404
rect 24820 7352 24826 7404
rect 25056 7401 25084 7432
rect 25222 7420 25228 7432
rect 25280 7420 25286 7472
rect 25041 7395 25099 7401
rect 25041 7361 25053 7395
rect 25087 7392 25099 7395
rect 25087 7364 25121 7392
rect 25087 7361 25099 7364
rect 25041 7355 25099 7361
rect 25314 7352 25320 7404
rect 25372 7352 25378 7404
rect 25406 7352 25412 7404
rect 25464 7352 25470 7404
rect 25498 7352 25504 7404
rect 25556 7352 25562 7404
rect 25608 7392 25636 7500
rect 31570 7488 31576 7540
rect 31628 7488 31634 7540
rect 31938 7488 31944 7540
rect 31996 7528 32002 7540
rect 32309 7531 32367 7537
rect 32309 7528 32321 7531
rect 31996 7500 32321 7528
rect 31996 7488 32002 7500
rect 32309 7497 32321 7500
rect 32355 7497 32367 7531
rect 32309 7491 32367 7497
rect 28813 7463 28871 7469
rect 26068 7432 26372 7460
rect 26068 7404 26096 7432
rect 25685 7395 25743 7401
rect 25685 7392 25697 7395
rect 25608 7364 25697 7392
rect 25685 7361 25697 7364
rect 25731 7361 25743 7395
rect 25685 7355 25743 7361
rect 26050 7352 26056 7404
rect 26108 7352 26114 7404
rect 26142 7352 26148 7404
rect 26200 7352 26206 7404
rect 26344 7401 26372 7432
rect 28813 7429 28825 7463
rect 28859 7460 28871 7463
rect 29089 7463 29147 7469
rect 29089 7460 29101 7463
rect 28859 7432 29101 7460
rect 28859 7429 28871 7432
rect 28813 7423 28871 7429
rect 29089 7429 29101 7432
rect 29135 7429 29147 7463
rect 31294 7460 31300 7472
rect 29089 7423 29147 7429
rect 31220 7432 31300 7460
rect 26329 7395 26387 7401
rect 26329 7361 26341 7395
rect 26375 7361 26387 7395
rect 26329 7355 26387 7361
rect 28718 7352 28724 7404
rect 28776 7352 28782 7404
rect 28905 7395 28963 7401
rect 28905 7361 28917 7395
rect 28951 7361 28963 7395
rect 28905 7355 28963 7361
rect 29273 7395 29331 7401
rect 29273 7361 29285 7395
rect 29319 7392 29331 7395
rect 30466 7392 30472 7404
rect 29319 7364 30472 7392
rect 29319 7361 29331 7364
rect 29273 7355 29331 7361
rect 22704 7296 22876 7324
rect 24029 7327 24087 7333
rect 22704 7284 22710 7296
rect 24029 7293 24041 7327
rect 24075 7293 24087 7327
rect 24029 7287 24087 7293
rect 24397 7327 24455 7333
rect 24397 7293 24409 7327
rect 24443 7324 24455 7327
rect 24780 7324 24808 7352
rect 24443 7296 24808 7324
rect 24443 7293 24455 7296
rect 24397 7287 24455 7293
rect 1673 7259 1731 7265
rect 1673 7225 1685 7259
rect 1719 7256 1731 7259
rect 1765 7259 1823 7265
rect 1765 7256 1777 7259
rect 1719 7228 1777 7256
rect 1719 7225 1731 7228
rect 1673 7219 1731 7225
rect 1765 7225 1777 7228
rect 1811 7256 1823 7259
rect 1854 7256 1860 7268
rect 1811 7228 1860 7256
rect 1811 7225 1823 7228
rect 1765 7219 1823 7225
rect 1854 7216 1860 7228
rect 1912 7216 1918 7268
rect 20257 7259 20315 7265
rect 20257 7225 20269 7259
rect 20303 7256 20315 7259
rect 20622 7256 20628 7268
rect 20303 7228 20628 7256
rect 20303 7225 20315 7228
rect 20257 7219 20315 7225
rect 20622 7216 20628 7228
rect 20680 7216 20686 7268
rect 24044 7256 24072 7287
rect 25130 7284 25136 7336
rect 25188 7284 25194 7336
rect 25314 7256 25320 7268
rect 24044 7228 25320 7256
rect 25314 7216 25320 7228
rect 25372 7216 25378 7268
rect 28920 7256 28948 7355
rect 30466 7352 30472 7364
rect 30524 7352 30530 7404
rect 31220 7401 31248 7432
rect 31294 7420 31300 7432
rect 31352 7420 31358 7472
rect 31205 7395 31263 7401
rect 31205 7361 31217 7395
rect 31251 7361 31263 7395
rect 31205 7355 31263 7361
rect 32214 7352 32220 7404
rect 32272 7352 32278 7404
rect 32324 7392 32352 7491
rect 32582 7488 32588 7540
rect 32640 7528 32646 7540
rect 32677 7531 32735 7537
rect 32677 7528 32689 7531
rect 32640 7500 32689 7528
rect 32640 7488 32646 7500
rect 32677 7497 32689 7500
rect 32723 7528 32735 7531
rect 32858 7528 32864 7540
rect 32723 7500 32864 7528
rect 32723 7497 32735 7500
rect 32677 7491 32735 7497
rect 32858 7488 32864 7500
rect 32916 7488 32922 7540
rect 33134 7488 33140 7540
rect 33192 7488 33198 7540
rect 33152 7460 33180 7488
rect 33152 7432 33994 7460
rect 32585 7395 32643 7401
rect 32585 7392 32597 7395
rect 32324 7364 32597 7392
rect 32585 7361 32597 7364
rect 32631 7392 32643 7395
rect 32674 7392 32680 7404
rect 32631 7364 32680 7392
rect 32631 7361 32643 7364
rect 32585 7355 32643 7361
rect 32674 7352 32680 7364
rect 32732 7352 32738 7404
rect 33045 7395 33103 7401
rect 33045 7361 33057 7395
rect 33091 7392 33103 7395
rect 33134 7392 33140 7404
rect 33091 7364 33140 7392
rect 33091 7361 33103 7364
rect 33045 7355 33103 7361
rect 33134 7352 33140 7364
rect 33192 7352 33198 7404
rect 31294 7284 31300 7336
rect 31352 7284 31358 7336
rect 32766 7284 32772 7336
rect 32824 7324 32830 7336
rect 33229 7327 33287 7333
rect 33229 7324 33241 7327
rect 32824 7296 33241 7324
rect 32824 7284 32830 7296
rect 33229 7293 33241 7296
rect 33275 7293 33287 7327
rect 33229 7287 33287 7293
rect 33502 7284 33508 7336
rect 33560 7284 33566 7336
rect 31846 7256 31852 7268
rect 28920 7228 31852 7256
rect 31846 7216 31852 7228
rect 31904 7216 31910 7268
rect 21542 7148 21548 7200
rect 21600 7148 21606 7200
rect 25222 7148 25228 7200
rect 25280 7188 25286 7200
rect 26421 7191 26479 7197
rect 26421 7188 26433 7191
rect 25280 7160 26433 7188
rect 25280 7148 25286 7160
rect 26421 7157 26433 7160
rect 26467 7157 26479 7191
rect 26421 7151 26479 7157
rect 29362 7148 29368 7200
rect 29420 7188 29426 7200
rect 31110 7188 31116 7200
rect 29420 7160 31116 7188
rect 29420 7148 29426 7160
rect 31110 7148 31116 7160
rect 31168 7148 31174 7200
rect 32953 7191 33011 7197
rect 32953 7157 32965 7191
rect 32999 7188 33011 7191
rect 33042 7188 33048 7200
rect 32999 7160 33048 7188
rect 32999 7157 33011 7160
rect 32953 7151 33011 7157
rect 33042 7148 33048 7160
rect 33100 7148 33106 7200
rect 34238 7148 34244 7200
rect 34296 7188 34302 7200
rect 34977 7191 35035 7197
rect 34977 7188 34989 7191
rect 34296 7160 34989 7188
rect 34296 7148 34302 7160
rect 34977 7157 34989 7160
rect 35023 7157 35035 7191
rect 34977 7151 35035 7157
rect 1104 7098 35328 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 35328 7098
rect 1104 7024 35328 7046
rect 10042 6944 10048 6996
rect 10100 6944 10106 6996
rect 11517 6987 11575 6993
rect 11517 6953 11529 6987
rect 11563 6984 11575 6987
rect 11606 6984 11612 6996
rect 11563 6956 11612 6984
rect 11563 6953 11575 6956
rect 11517 6947 11575 6953
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 17310 6944 17316 6996
rect 17368 6944 17374 6996
rect 17678 6944 17684 6996
rect 17736 6984 17742 6996
rect 17865 6987 17923 6993
rect 17865 6984 17877 6987
rect 17736 6956 17877 6984
rect 17736 6944 17742 6956
rect 17865 6953 17877 6956
rect 17911 6953 17923 6987
rect 17865 6947 17923 6953
rect 20257 6987 20315 6993
rect 20257 6953 20269 6987
rect 20303 6984 20315 6987
rect 20346 6984 20352 6996
rect 20303 6956 20352 6984
rect 20303 6953 20315 6956
rect 20257 6947 20315 6953
rect 20346 6944 20352 6956
rect 20404 6944 20410 6996
rect 21266 6944 21272 6996
rect 21324 6984 21330 6996
rect 21729 6987 21787 6993
rect 21729 6984 21741 6987
rect 21324 6956 21741 6984
rect 21324 6944 21330 6956
rect 21729 6953 21741 6956
rect 21775 6953 21787 6987
rect 21729 6947 21787 6953
rect 22738 6944 22744 6996
rect 22796 6984 22802 6996
rect 23658 6984 23664 6996
rect 22796 6956 23664 6984
rect 22796 6944 22802 6956
rect 23658 6944 23664 6956
rect 23716 6984 23722 6996
rect 24029 6987 24087 6993
rect 24029 6984 24041 6987
rect 23716 6956 24041 6984
rect 23716 6944 23722 6956
rect 24029 6953 24041 6956
rect 24075 6953 24087 6987
rect 24029 6947 24087 6953
rect 24857 6987 24915 6993
rect 24857 6953 24869 6987
rect 24903 6984 24915 6987
rect 25222 6984 25228 6996
rect 24903 6956 25228 6984
rect 24903 6953 24915 6956
rect 24857 6947 24915 6953
rect 25222 6944 25228 6956
rect 25280 6944 25286 6996
rect 26050 6944 26056 6996
rect 26108 6944 26114 6996
rect 26142 6944 26148 6996
rect 26200 6984 26206 6996
rect 27537 6987 27595 6993
rect 27537 6984 27549 6987
rect 26200 6956 27549 6984
rect 26200 6944 26206 6956
rect 27537 6953 27549 6956
rect 27583 6953 27595 6987
rect 27537 6947 27595 6953
rect 31846 6944 31852 6996
rect 31904 6984 31910 6996
rect 32217 6987 32275 6993
rect 32217 6984 32229 6987
rect 31904 6956 32229 6984
rect 31904 6944 31910 6956
rect 32217 6953 32229 6956
rect 32263 6984 32275 6987
rect 32263 6956 32996 6984
rect 32263 6953 32275 6956
rect 32217 6947 32275 6953
rect 25038 6876 25044 6928
rect 25096 6916 25102 6928
rect 25314 6916 25320 6928
rect 25096 6888 25320 6916
rect 25096 6876 25102 6888
rect 25314 6876 25320 6888
rect 25372 6916 25378 6928
rect 25372 6888 25544 6916
rect 25372 6876 25378 6888
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 10505 6851 10563 6857
rect 10505 6848 10517 6851
rect 9732 6820 10517 6848
rect 9732 6808 9738 6820
rect 10505 6817 10517 6820
rect 10551 6817 10563 6851
rect 10505 6811 10563 6817
rect 10689 6851 10747 6857
rect 10689 6817 10701 6851
rect 10735 6848 10747 6851
rect 11425 6851 11483 6857
rect 10735 6820 11008 6848
rect 10735 6817 10747 6820
rect 10689 6811 10747 6817
rect 10134 6740 10140 6792
rect 10192 6780 10198 6792
rect 10413 6783 10471 6789
rect 10413 6780 10425 6783
rect 10192 6752 10425 6780
rect 10192 6740 10198 6752
rect 10413 6749 10425 6752
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 10980 6721 11008 6820
rect 11425 6817 11437 6851
rect 11471 6848 11483 6851
rect 11974 6848 11980 6860
rect 11471 6820 11980 6848
rect 11471 6817 11483 6820
rect 11425 6811 11483 6817
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6848 12219 6851
rect 12434 6848 12440 6860
rect 12207 6820 12440 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 12434 6808 12440 6820
rect 12492 6808 12498 6860
rect 15930 6808 15936 6860
rect 15988 6808 15994 6860
rect 18509 6851 18567 6857
rect 18509 6817 18521 6851
rect 18555 6817 18567 6851
rect 18509 6811 18567 6817
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6780 11943 6783
rect 12710 6780 12716 6792
rect 11931 6752 12716 6780
rect 11931 6749 11943 6752
rect 11885 6743 11943 6749
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 14093 6783 14151 6789
rect 14093 6749 14105 6783
rect 14139 6780 14151 6783
rect 15948 6780 15976 6808
rect 14139 6752 15976 6780
rect 16200 6783 16258 6789
rect 14139 6749 14151 6752
rect 14093 6743 14151 6749
rect 16200 6749 16212 6783
rect 16246 6780 16258 6783
rect 16482 6780 16488 6792
rect 16246 6752 16488 6780
rect 16246 6749 16258 6752
rect 16200 6743 16258 6749
rect 16482 6740 16488 6752
rect 16540 6740 16546 6792
rect 16942 6740 16948 6792
rect 17000 6780 17006 6792
rect 18233 6783 18291 6789
rect 18233 6780 18245 6783
rect 17000 6752 18245 6780
rect 17000 6740 17006 6752
rect 18233 6749 18245 6752
rect 18279 6749 18291 6783
rect 18524 6780 18552 6811
rect 18874 6808 18880 6860
rect 18932 6848 18938 6860
rect 20349 6851 20407 6857
rect 20349 6848 20361 6851
rect 18932 6820 20361 6848
rect 18932 6808 18938 6820
rect 20349 6817 20361 6820
rect 20395 6817 20407 6851
rect 20349 6811 20407 6817
rect 18785 6783 18843 6789
rect 18785 6780 18797 6783
rect 18524 6752 18797 6780
rect 18233 6743 18291 6749
rect 18785 6749 18797 6752
rect 18831 6780 18843 6783
rect 19702 6780 19708 6792
rect 18831 6752 19708 6780
rect 18831 6749 18843 6752
rect 18785 6743 18843 6749
rect 19702 6740 19708 6752
rect 19760 6740 19766 6792
rect 20364 6780 20392 6811
rect 23198 6808 23204 6860
rect 23256 6848 23262 6860
rect 24555 6851 24613 6857
rect 24555 6848 24567 6851
rect 23256 6820 24567 6848
rect 23256 6808 23262 6820
rect 24555 6817 24567 6820
rect 24601 6817 24613 6851
rect 25516 6848 25544 6888
rect 27798 6876 27804 6928
rect 27856 6916 27862 6928
rect 28718 6916 28724 6928
rect 27856 6888 28724 6916
rect 27856 6876 27862 6888
rect 28718 6876 28724 6888
rect 28776 6916 28782 6928
rect 28776 6888 30972 6916
rect 28776 6876 28782 6888
rect 25958 6848 25964 6860
rect 24555 6811 24613 6817
rect 24780 6820 25452 6848
rect 24780 6792 24808 6820
rect 21913 6783 21971 6789
rect 21913 6780 21925 6783
rect 20364 6752 21925 6780
rect 21913 6749 21925 6752
rect 21959 6780 21971 6783
rect 22278 6780 22284 6792
rect 21959 6752 22284 6780
rect 21959 6749 21971 6752
rect 21913 6743 21971 6749
rect 22278 6740 22284 6752
rect 22336 6740 22342 6792
rect 22741 6783 22799 6789
rect 22741 6749 22753 6783
rect 22787 6780 22799 6783
rect 22830 6780 22836 6792
rect 22787 6752 22836 6780
rect 22787 6749 22799 6752
rect 22741 6743 22799 6749
rect 22830 6740 22836 6752
rect 22888 6740 22894 6792
rect 23382 6740 23388 6792
rect 23440 6740 23446 6792
rect 23658 6740 23664 6792
rect 23716 6740 23722 6792
rect 23753 6783 23811 6789
rect 23753 6749 23765 6783
rect 23799 6749 23811 6783
rect 23753 6743 23811 6749
rect 10965 6715 11023 6721
rect 10965 6681 10977 6715
rect 11011 6712 11023 6715
rect 12434 6712 12440 6724
rect 11011 6684 12440 6712
rect 11011 6681 11023 6684
rect 10965 6675 11023 6681
rect 12434 6672 12440 6684
rect 12492 6672 12498 6724
rect 14182 6672 14188 6724
rect 14240 6712 14246 6724
rect 14338 6715 14396 6721
rect 14338 6712 14350 6715
rect 14240 6684 14350 6712
rect 14240 6672 14246 6684
rect 14338 6681 14350 6684
rect 14384 6681 14396 6715
rect 14338 6675 14396 6681
rect 18325 6715 18383 6721
rect 18325 6681 18337 6715
rect 18371 6712 18383 6715
rect 18414 6712 18420 6724
rect 18371 6684 18420 6712
rect 18371 6681 18383 6684
rect 18325 6675 18383 6681
rect 18414 6672 18420 6684
rect 18472 6672 18478 6724
rect 20616 6715 20674 6721
rect 20616 6681 20628 6715
rect 20662 6712 20674 6715
rect 20806 6712 20812 6724
rect 20662 6684 20812 6712
rect 20662 6681 20674 6684
rect 20616 6675 20674 6681
rect 20806 6672 20812 6684
rect 20864 6672 20870 6724
rect 23474 6672 23480 6724
rect 23532 6712 23538 6724
rect 23768 6712 23796 6743
rect 24394 6740 24400 6792
rect 24452 6740 24458 6792
rect 24762 6740 24768 6792
rect 24820 6740 24826 6792
rect 25041 6783 25099 6789
rect 25041 6749 25053 6783
rect 25087 6780 25099 6783
rect 25222 6780 25228 6792
rect 25087 6752 25228 6780
rect 25087 6749 25099 6752
rect 25041 6743 25099 6749
rect 25222 6740 25228 6752
rect 25280 6740 25286 6792
rect 25424 6789 25452 6820
rect 25516 6820 25964 6848
rect 25516 6789 25544 6820
rect 25958 6808 25964 6820
rect 26016 6848 26022 6860
rect 27890 6848 27896 6860
rect 26016 6820 27896 6848
rect 26016 6808 26022 6820
rect 27890 6808 27896 6820
rect 27948 6808 27954 6860
rect 28629 6851 28687 6857
rect 28629 6817 28641 6851
rect 28675 6848 28687 6851
rect 28810 6848 28816 6860
rect 28675 6820 28816 6848
rect 28675 6817 28687 6820
rect 28629 6811 28687 6817
rect 28810 6808 28816 6820
rect 28868 6808 28874 6860
rect 29089 6851 29147 6857
rect 29089 6817 29101 6851
rect 29135 6848 29147 6851
rect 30190 6848 30196 6860
rect 29135 6820 30196 6848
rect 29135 6817 29147 6820
rect 29089 6811 29147 6817
rect 30190 6808 30196 6820
rect 30248 6848 30254 6860
rect 30837 6851 30895 6857
rect 30837 6848 30849 6851
rect 30248 6820 30849 6848
rect 30248 6808 30254 6820
rect 30837 6817 30849 6820
rect 30883 6817 30895 6851
rect 30944 6848 30972 6888
rect 31662 6876 31668 6928
rect 31720 6876 31726 6928
rect 31754 6876 31760 6928
rect 31812 6916 31818 6928
rect 32398 6916 32404 6928
rect 31812 6888 32404 6916
rect 31812 6876 31818 6888
rect 32398 6876 32404 6888
rect 32456 6876 32462 6928
rect 32968 6925 32996 6956
rect 33502 6944 33508 6996
rect 33560 6984 33566 6996
rect 33873 6987 33931 6993
rect 33873 6984 33885 6987
rect 33560 6956 33885 6984
rect 33560 6944 33566 6956
rect 33873 6953 33885 6956
rect 33919 6953 33931 6987
rect 33873 6947 33931 6953
rect 32953 6919 33011 6925
rect 32953 6885 32965 6919
rect 32999 6885 33011 6919
rect 32953 6879 33011 6885
rect 33042 6876 33048 6928
rect 33100 6916 33106 6928
rect 33100 6888 33456 6916
rect 33100 6876 33106 6888
rect 31570 6848 31576 6860
rect 30944 6820 31576 6848
rect 30837 6811 30895 6817
rect 31570 6808 31576 6820
rect 31628 6808 31634 6860
rect 31680 6848 31708 6876
rect 33428 6860 33456 6888
rect 31680 6820 32536 6848
rect 25409 6783 25467 6789
rect 25409 6749 25421 6783
rect 25455 6749 25467 6783
rect 25409 6743 25467 6749
rect 25501 6783 25559 6789
rect 25501 6749 25513 6783
rect 25547 6749 25559 6783
rect 25501 6743 25559 6749
rect 27801 6783 27859 6789
rect 27801 6749 27813 6783
rect 27847 6749 27859 6783
rect 27801 6743 27859 6749
rect 24578 6712 24584 6724
rect 23532 6684 23796 6712
rect 23952 6684 24584 6712
rect 23532 6672 23538 6684
rect 14642 6604 14648 6656
rect 14700 6644 14706 6656
rect 15473 6647 15531 6653
rect 15473 6644 15485 6647
rect 14700 6616 15485 6644
rect 14700 6604 14706 6616
rect 15473 6613 15485 6616
rect 15519 6613 15531 6647
rect 15473 6607 15531 6613
rect 21082 6604 21088 6656
rect 21140 6644 21146 6656
rect 23952 6653 23980 6684
rect 24578 6672 24584 6684
rect 24636 6672 24642 6724
rect 24946 6672 24952 6724
rect 25004 6712 25010 6724
rect 25133 6715 25191 6721
rect 25133 6712 25145 6715
rect 25004 6684 25145 6712
rect 25004 6672 25010 6684
rect 25133 6681 25145 6684
rect 25179 6681 25191 6715
rect 26050 6712 26056 6724
rect 25133 6675 25191 6681
rect 25240 6684 26056 6712
rect 23937 6647 23995 6653
rect 23937 6644 23949 6647
rect 21140 6616 23949 6644
rect 21140 6604 21146 6616
rect 23937 6613 23949 6616
rect 23983 6613 23995 6647
rect 23937 6607 23995 6613
rect 24486 6604 24492 6656
rect 24544 6644 24550 6656
rect 25240 6644 25268 6684
rect 26050 6672 26056 6684
rect 26108 6712 26114 6724
rect 27816 6712 27844 6743
rect 28994 6740 29000 6792
rect 29052 6740 29058 6792
rect 29914 6740 29920 6792
rect 29972 6740 29978 6792
rect 31021 6783 31079 6789
rect 31021 6749 31033 6783
rect 31067 6749 31079 6783
rect 31021 6743 31079 6749
rect 29932 6712 29960 6740
rect 26108 6684 26358 6712
rect 27816 6684 29960 6712
rect 31036 6712 31064 6743
rect 31110 6740 31116 6792
rect 31168 6780 31174 6792
rect 31297 6783 31355 6789
rect 31297 6780 31309 6783
rect 31168 6752 31309 6780
rect 31168 6740 31174 6752
rect 31297 6749 31309 6752
rect 31343 6780 31355 6783
rect 31481 6783 31539 6789
rect 31481 6780 31493 6783
rect 31343 6752 31493 6780
rect 31343 6749 31355 6752
rect 31297 6743 31355 6749
rect 31481 6749 31493 6752
rect 31527 6749 31539 6783
rect 31481 6743 31539 6749
rect 31665 6783 31723 6789
rect 31665 6749 31677 6783
rect 31711 6780 31723 6783
rect 31754 6780 31760 6792
rect 31711 6752 31760 6780
rect 31711 6749 31723 6752
rect 31665 6743 31723 6749
rect 31754 6740 31760 6752
rect 31812 6740 31818 6792
rect 31846 6740 31852 6792
rect 31904 6740 31910 6792
rect 31938 6740 31944 6792
rect 31996 6780 32002 6792
rect 32508 6789 32536 6820
rect 33410 6808 33416 6860
rect 33468 6808 33474 6860
rect 32493 6783 32551 6789
rect 31996 6752 32168 6780
rect 31996 6740 32002 6752
rect 32140 6712 32168 6752
rect 32493 6749 32505 6783
rect 32539 6749 32551 6783
rect 32493 6743 32551 6749
rect 32582 6740 32588 6792
rect 32640 6740 32646 6792
rect 32769 6783 32827 6789
rect 32769 6749 32781 6783
rect 32815 6749 32827 6783
rect 32769 6743 32827 6749
rect 32196 6715 32254 6721
rect 32196 6712 32208 6715
rect 31036 6684 32076 6712
rect 32140 6684 32208 6712
rect 26108 6672 26114 6684
rect 24544 6616 25268 6644
rect 24544 6604 24550 6616
rect 25314 6604 25320 6656
rect 25372 6604 25378 6656
rect 25682 6604 25688 6656
rect 25740 6604 25746 6656
rect 26878 6604 26884 6656
rect 26936 6644 26942 6656
rect 27338 6644 27344 6656
rect 26936 6616 27344 6644
rect 26936 6604 26942 6616
rect 27338 6604 27344 6616
rect 27396 6644 27402 6656
rect 27816 6644 27844 6684
rect 27396 6616 27844 6644
rect 27396 6604 27402 6616
rect 27890 6604 27896 6656
rect 27948 6644 27954 6656
rect 30834 6644 30840 6656
rect 27948 6616 30840 6644
rect 27948 6604 27954 6616
rect 30834 6604 30840 6616
rect 30892 6604 30898 6656
rect 31205 6647 31263 6653
rect 31205 6613 31217 6647
rect 31251 6644 31263 6647
rect 31386 6644 31392 6656
rect 31251 6616 31392 6644
rect 31251 6613 31263 6616
rect 31205 6607 31263 6613
rect 31386 6604 31392 6616
rect 31444 6604 31450 6656
rect 31570 6604 31576 6656
rect 31628 6644 31634 6656
rect 31938 6644 31944 6656
rect 31628 6616 31944 6644
rect 31628 6604 31634 6616
rect 31938 6604 31944 6616
rect 31996 6604 32002 6656
rect 32048 6653 32076 6684
rect 32196 6681 32208 6684
rect 32242 6712 32254 6715
rect 32306 6712 32312 6724
rect 32242 6684 32312 6712
rect 32242 6681 32254 6684
rect 32196 6675 32254 6681
rect 32306 6672 32312 6684
rect 32364 6672 32370 6724
rect 32398 6672 32404 6724
rect 32456 6672 32462 6724
rect 32033 6647 32091 6653
rect 32033 6613 32045 6647
rect 32079 6613 32091 6647
rect 32784 6644 32812 6743
rect 32858 6740 32864 6792
rect 32916 6780 32922 6792
rect 33137 6783 33195 6789
rect 33137 6780 33149 6783
rect 32916 6752 33149 6780
rect 32916 6740 32922 6752
rect 33137 6749 33149 6752
rect 33183 6780 33195 6783
rect 33689 6783 33747 6789
rect 33689 6780 33701 6783
rect 33183 6752 33701 6780
rect 33183 6749 33195 6752
rect 33137 6743 33195 6749
rect 33689 6749 33701 6752
rect 33735 6749 33747 6783
rect 33689 6743 33747 6749
rect 34054 6740 34060 6792
rect 34112 6740 34118 6792
rect 34238 6740 34244 6792
rect 34296 6740 34302 6792
rect 34333 6783 34391 6789
rect 34333 6749 34345 6783
rect 34379 6780 34391 6783
rect 34422 6780 34428 6792
rect 34379 6752 34428 6780
rect 34379 6749 34391 6752
rect 34333 6743 34391 6749
rect 33410 6672 33416 6724
rect 33468 6672 33474 6724
rect 33597 6715 33655 6721
rect 33597 6681 33609 6715
rect 33643 6712 33655 6715
rect 34348 6712 34376 6743
rect 34422 6740 34428 6752
rect 34480 6740 34486 6792
rect 33643 6684 34376 6712
rect 33643 6681 33655 6684
rect 33597 6675 33655 6681
rect 33612 6644 33640 6675
rect 32784 6616 33640 6644
rect 32033 6607 32091 6613
rect 1104 6554 35328 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35328 6554
rect 1104 6480 35328 6502
rect 14182 6400 14188 6452
rect 14240 6400 14246 6452
rect 14550 6400 14556 6452
rect 14608 6400 14614 6452
rect 14642 6400 14648 6452
rect 14700 6400 14706 6452
rect 15010 6400 15016 6452
rect 15068 6400 15074 6452
rect 21269 6443 21327 6449
rect 21269 6409 21281 6443
rect 21315 6440 21327 6443
rect 23106 6440 23112 6452
rect 21315 6412 23112 6440
rect 21315 6409 21327 6412
rect 21269 6403 21327 6409
rect 23106 6400 23112 6412
rect 23164 6400 23170 6452
rect 23750 6440 23756 6452
rect 23216 6412 23756 6440
rect 23216 6372 23244 6412
rect 23750 6400 23756 6412
rect 23808 6400 23814 6452
rect 24578 6400 24584 6452
rect 24636 6440 24642 6452
rect 25314 6440 25320 6452
rect 24636 6412 25320 6440
rect 24636 6400 24642 6412
rect 25314 6400 25320 6412
rect 25372 6400 25378 6452
rect 25777 6443 25835 6449
rect 25777 6409 25789 6443
rect 25823 6440 25835 6443
rect 26142 6440 26148 6452
rect 25823 6412 26148 6440
rect 25823 6409 25835 6412
rect 25777 6403 25835 6409
rect 26142 6400 26148 6412
rect 26200 6400 26206 6452
rect 26234 6400 26240 6452
rect 26292 6440 26298 6452
rect 26292 6412 28028 6440
rect 26292 6400 26298 6412
rect 28000 6372 28028 6412
rect 28810 6400 28816 6452
rect 28868 6400 28874 6452
rect 29454 6440 29460 6452
rect 28966 6412 29460 6440
rect 28966 6372 28994 6412
rect 29454 6400 29460 6412
rect 29512 6400 29518 6452
rect 31202 6400 31208 6452
rect 31260 6400 31266 6452
rect 31294 6400 31300 6452
rect 31352 6400 31358 6452
rect 32125 6443 32183 6449
rect 32125 6409 32137 6443
rect 32171 6440 32183 6443
rect 32214 6440 32220 6452
rect 32171 6412 32220 6440
rect 32171 6409 32183 6412
rect 32125 6403 32183 6409
rect 32214 6400 32220 6412
rect 32272 6400 32278 6452
rect 32306 6400 32312 6452
rect 32364 6440 32370 6452
rect 32769 6443 32827 6449
rect 32769 6440 32781 6443
rect 32364 6412 32781 6440
rect 32364 6400 32370 6412
rect 32769 6409 32781 6412
rect 32815 6409 32827 6443
rect 32769 6403 32827 6409
rect 33410 6400 33416 6452
rect 33468 6400 33474 6452
rect 21284 6344 23244 6372
rect 23492 6344 27936 6372
rect 28000 6344 28994 6372
rect 21082 6264 21088 6316
rect 21140 6264 21146 6316
rect 21284 6313 21312 6344
rect 21269 6307 21327 6313
rect 21269 6273 21281 6307
rect 21315 6273 21327 6307
rect 21269 6267 21327 6273
rect 21453 6307 21511 6313
rect 21453 6273 21465 6307
rect 21499 6304 21511 6307
rect 21499 6276 22232 6304
rect 21499 6273 21511 6276
rect 21453 6267 21511 6273
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6236 14887 6239
rect 15010 6236 15016 6248
rect 14875 6208 15016 6236
rect 14875 6205 14887 6208
rect 14829 6199 14887 6205
rect 15010 6196 15016 6208
rect 15068 6196 15074 6248
rect 22204 6236 22232 6276
rect 22278 6264 22284 6316
rect 22336 6264 22342 6316
rect 23492 6313 23520 6344
rect 23109 6307 23167 6313
rect 23109 6273 23121 6307
rect 23155 6304 23167 6307
rect 23477 6307 23535 6313
rect 23477 6304 23489 6307
rect 23155 6276 23489 6304
rect 23155 6273 23167 6276
rect 23109 6267 23167 6273
rect 23477 6273 23489 6276
rect 23523 6273 23535 6307
rect 23477 6267 23535 6273
rect 23658 6264 23664 6316
rect 23716 6304 23722 6316
rect 23753 6307 23811 6313
rect 23753 6304 23765 6307
rect 23716 6276 23765 6304
rect 23716 6264 23722 6276
rect 23753 6273 23765 6276
rect 23799 6304 23811 6307
rect 24486 6304 24492 6316
rect 23799 6276 24492 6304
rect 23799 6273 23811 6276
rect 23753 6267 23811 6273
rect 24486 6264 24492 6276
rect 24544 6264 24550 6316
rect 24578 6264 24584 6316
rect 24636 6264 24642 6316
rect 24765 6307 24823 6313
rect 24765 6273 24777 6307
rect 24811 6273 24823 6307
rect 24765 6267 24823 6273
rect 24857 6307 24915 6313
rect 24857 6273 24869 6307
rect 24903 6304 24915 6307
rect 25038 6304 25044 6316
rect 24903 6276 25044 6304
rect 24903 6273 24915 6276
rect 24857 6267 24915 6273
rect 22204 6208 22692 6236
rect 21545 6103 21603 6109
rect 21545 6069 21557 6103
rect 21591 6100 21603 6103
rect 22462 6100 22468 6112
rect 21591 6072 22468 6100
rect 21591 6069 21603 6072
rect 21545 6063 21603 6069
rect 22462 6060 22468 6072
rect 22520 6060 22526 6112
rect 22664 6100 22692 6208
rect 23382 6196 23388 6248
rect 23440 6236 23446 6248
rect 23440 6208 23796 6236
rect 23440 6196 23446 6208
rect 23768 6168 23796 6208
rect 23842 6196 23848 6248
rect 23900 6236 23906 6248
rect 24780 6236 24808 6267
rect 25038 6264 25044 6276
rect 25096 6264 25102 6316
rect 25130 6264 25136 6316
rect 25188 6304 25194 6316
rect 25409 6307 25467 6313
rect 25409 6304 25421 6307
rect 25188 6276 25421 6304
rect 25188 6264 25194 6276
rect 25409 6273 25421 6276
rect 25455 6273 25467 6307
rect 25409 6267 25467 6273
rect 24946 6236 24952 6248
rect 23900 6208 24952 6236
rect 23900 6196 23906 6208
rect 24946 6196 24952 6208
rect 25004 6196 25010 6248
rect 25501 6239 25559 6245
rect 25501 6205 25513 6239
rect 25547 6236 25559 6239
rect 25682 6236 25688 6248
rect 25547 6208 25688 6236
rect 25547 6205 25559 6208
rect 25501 6199 25559 6205
rect 25682 6196 25688 6208
rect 25740 6196 25746 6248
rect 23768 6140 25084 6168
rect 25056 6112 25084 6140
rect 25222 6128 25228 6180
rect 25280 6168 25286 6180
rect 27798 6168 27804 6180
rect 25280 6140 27804 6168
rect 25280 6128 25286 6140
rect 27798 6128 27804 6140
rect 27856 6128 27862 6180
rect 27908 6168 27936 6344
rect 29086 6332 29092 6384
rect 29144 6372 29150 6384
rect 29181 6375 29239 6381
rect 29181 6372 29193 6375
rect 29144 6344 29193 6372
rect 29144 6332 29150 6344
rect 29181 6341 29193 6344
rect 29227 6372 29239 6375
rect 31220 6372 31248 6400
rect 31573 6375 31631 6381
rect 31573 6372 31585 6375
rect 29227 6344 31248 6372
rect 31404 6344 31585 6372
rect 29227 6341 29239 6344
rect 29181 6335 29239 6341
rect 28721 6307 28779 6313
rect 28721 6273 28733 6307
rect 28767 6304 28779 6307
rect 28810 6304 28816 6316
rect 28767 6276 28816 6304
rect 28767 6273 28779 6276
rect 28721 6267 28779 6273
rect 28810 6264 28816 6276
rect 28868 6264 28874 6316
rect 28994 6264 29000 6316
rect 29052 6304 29058 6316
rect 30006 6304 30012 6316
rect 29052 6276 30012 6304
rect 29052 6264 29058 6276
rect 30006 6264 30012 6276
rect 30064 6304 30070 6316
rect 30561 6307 30619 6313
rect 30064 6276 30236 6304
rect 30064 6264 30070 6276
rect 28905 6239 28963 6245
rect 28905 6205 28917 6239
rect 28951 6236 28963 6239
rect 29362 6236 29368 6248
rect 28951 6208 29368 6236
rect 28951 6205 28963 6208
rect 28905 6199 28963 6205
rect 29362 6196 29368 6208
rect 29420 6236 29426 6248
rect 29730 6236 29736 6248
rect 29420 6208 29736 6236
rect 29420 6196 29426 6208
rect 29730 6196 29736 6208
rect 29788 6196 29794 6248
rect 29914 6196 29920 6248
rect 29972 6196 29978 6248
rect 30208 6245 30236 6276
rect 30561 6273 30573 6307
rect 30607 6304 30619 6307
rect 30742 6304 30748 6316
rect 30607 6276 30748 6304
rect 30607 6273 30619 6276
rect 30561 6267 30619 6273
rect 30742 6264 30748 6276
rect 30800 6264 30806 6316
rect 31110 6264 31116 6316
rect 31168 6304 31174 6316
rect 31404 6313 31432 6344
rect 31573 6341 31585 6344
rect 31619 6341 31631 6375
rect 33042 6372 33048 6384
rect 31573 6335 31631 6341
rect 32324 6344 33048 6372
rect 31205 6307 31263 6313
rect 31205 6304 31217 6307
rect 31168 6276 31217 6304
rect 31168 6264 31174 6276
rect 31205 6273 31217 6276
rect 31251 6273 31263 6307
rect 31205 6267 31263 6273
rect 31389 6307 31447 6313
rect 31389 6273 31401 6307
rect 31435 6273 31447 6307
rect 31389 6267 31447 6273
rect 31478 6264 31484 6316
rect 31536 6264 31542 6316
rect 31662 6264 31668 6316
rect 31720 6264 31726 6316
rect 32324 6313 32352 6344
rect 33042 6332 33048 6344
rect 33100 6372 33106 6384
rect 33597 6375 33655 6381
rect 33597 6372 33609 6375
rect 33100 6344 33609 6372
rect 33100 6332 33106 6344
rect 33597 6341 33609 6344
rect 33643 6341 33655 6375
rect 33597 6335 33655 6341
rect 32309 6307 32367 6313
rect 32309 6304 32321 6307
rect 31864 6276 32321 6304
rect 30193 6239 30251 6245
rect 30193 6205 30205 6239
rect 30239 6205 30251 6239
rect 30193 6199 30251 6205
rect 30466 6196 30472 6248
rect 30524 6236 30530 6248
rect 31680 6236 31708 6264
rect 30524 6208 31708 6236
rect 30524 6196 30530 6208
rect 27908 6140 28994 6168
rect 23658 6100 23664 6112
rect 22664 6072 23664 6100
rect 23658 6060 23664 6072
rect 23716 6060 23722 6112
rect 23750 6060 23756 6112
rect 23808 6100 23814 6112
rect 24397 6103 24455 6109
rect 24397 6100 24409 6103
rect 23808 6072 24409 6100
rect 23808 6060 23814 6072
rect 24397 6069 24409 6072
rect 24443 6069 24455 6103
rect 24397 6063 24455 6069
rect 25038 6060 25044 6112
rect 25096 6100 25102 6112
rect 26234 6100 26240 6112
rect 25096 6072 26240 6100
rect 25096 6060 25102 6072
rect 26234 6060 26240 6072
rect 26292 6060 26298 6112
rect 27430 6060 27436 6112
rect 27488 6100 27494 6112
rect 28353 6103 28411 6109
rect 28353 6100 28365 6103
rect 27488 6072 28365 6100
rect 27488 6060 27494 6072
rect 28353 6069 28365 6072
rect 28399 6069 28411 6103
rect 28966 6100 28994 6140
rect 29822 6128 29828 6180
rect 29880 6168 29886 6180
rect 31864 6177 31892 6276
rect 32309 6273 32321 6276
rect 32355 6273 32367 6307
rect 32309 6267 32367 6273
rect 32858 6264 32864 6316
rect 32916 6264 32922 6316
rect 33321 6307 33379 6313
rect 33321 6304 33333 6307
rect 32968 6276 33333 6304
rect 32585 6239 32643 6245
rect 32585 6205 32597 6239
rect 32631 6236 32643 6239
rect 32968 6236 32996 6276
rect 33321 6273 33333 6276
rect 33367 6304 33379 6307
rect 34422 6304 34428 6316
rect 33367 6276 34428 6304
rect 33367 6273 33379 6276
rect 33321 6267 33379 6273
rect 34422 6264 34428 6276
rect 34480 6264 34486 6316
rect 33042 6245 33048 6248
rect 32631 6208 32996 6236
rect 32631 6205 32643 6208
rect 32585 6199 32643 6205
rect 33041 6199 33048 6245
rect 33100 6236 33106 6248
rect 33100 6208 33141 6236
rect 33042 6196 33048 6199
rect 33100 6196 33106 6208
rect 31849 6171 31907 6177
rect 31849 6168 31861 6171
rect 29880 6140 31861 6168
rect 29880 6128 29886 6140
rect 31849 6137 31861 6140
rect 31895 6137 31907 6171
rect 31849 6131 31907 6137
rect 32508 6140 33088 6168
rect 32508 6112 32536 6140
rect 31294 6100 31300 6112
rect 28966 6072 31300 6100
rect 28353 6063 28411 6069
rect 31294 6060 31300 6072
rect 31352 6060 31358 6112
rect 32490 6060 32496 6112
rect 32548 6060 32554 6112
rect 33060 6100 33088 6140
rect 33134 6128 33140 6180
rect 33192 6128 33198 6180
rect 33226 6100 33232 6112
rect 33060 6072 33232 6100
rect 33226 6060 33232 6072
rect 33284 6060 33290 6112
rect 1104 6010 35328 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 35328 6010
rect 1104 5936 35328 5958
rect 22925 5899 22983 5905
rect 2746 5868 22876 5896
rect 1854 5720 1860 5772
rect 1912 5760 1918 5772
rect 2746 5760 2774 5868
rect 22848 5828 22876 5868
rect 22925 5865 22937 5899
rect 22971 5896 22983 5899
rect 23474 5896 23480 5908
rect 22971 5868 23480 5896
rect 22971 5865 22983 5868
rect 22925 5859 22983 5865
rect 23474 5856 23480 5868
rect 23532 5856 23538 5908
rect 24394 5856 24400 5908
rect 24452 5896 24458 5908
rect 25406 5896 25412 5908
rect 24452 5868 25412 5896
rect 24452 5856 24458 5868
rect 25406 5856 25412 5868
rect 25464 5896 25470 5908
rect 25464 5868 28488 5896
rect 25464 5856 25470 5868
rect 22848 5800 27016 5828
rect 1912 5732 2774 5760
rect 21177 5763 21235 5769
rect 1912 5720 1918 5732
rect 21177 5729 21189 5763
rect 21223 5760 21235 5763
rect 22186 5760 22192 5772
rect 21223 5732 22192 5760
rect 21223 5729 21235 5732
rect 21177 5723 21235 5729
rect 22186 5720 22192 5732
rect 22244 5720 22250 5772
rect 22462 5720 22468 5772
rect 22520 5760 22526 5772
rect 23382 5760 23388 5772
rect 22520 5732 23388 5760
rect 22520 5720 22526 5732
rect 22572 5678 22600 5732
rect 23382 5720 23388 5732
rect 23440 5720 23446 5772
rect 23477 5763 23535 5769
rect 23477 5729 23489 5763
rect 23523 5760 23535 5763
rect 23934 5760 23940 5772
rect 23523 5732 23940 5760
rect 23523 5729 23535 5732
rect 23477 5723 23535 5729
rect 23934 5720 23940 5732
rect 23992 5720 23998 5772
rect 24121 5763 24179 5769
rect 24121 5729 24133 5763
rect 24167 5760 24179 5763
rect 25038 5760 25044 5772
rect 24167 5732 25044 5760
rect 24167 5729 24179 5732
rect 24121 5723 24179 5729
rect 25038 5720 25044 5732
rect 25096 5720 25102 5772
rect 23569 5695 23627 5701
rect 23569 5692 23581 5695
rect 22848 5664 23581 5692
rect 21453 5627 21511 5633
rect 21453 5593 21465 5627
rect 21499 5593 21511 5627
rect 21453 5587 21511 5593
rect 21468 5556 21496 5587
rect 22848 5556 22876 5664
rect 23569 5661 23581 5664
rect 23615 5661 23627 5695
rect 23569 5655 23627 5661
rect 23750 5652 23756 5704
rect 23808 5652 23814 5704
rect 25222 5692 25228 5704
rect 23860 5664 25228 5692
rect 23106 5584 23112 5636
rect 23164 5584 23170 5636
rect 23198 5584 23204 5636
rect 23256 5624 23262 5636
rect 23293 5627 23351 5633
rect 23293 5624 23305 5627
rect 23256 5596 23305 5624
rect 23256 5584 23262 5596
rect 23293 5593 23305 5596
rect 23339 5593 23351 5627
rect 23293 5587 23351 5593
rect 21468 5528 22876 5556
rect 23309 5556 23337 5587
rect 23860 5556 23888 5664
rect 25222 5652 25228 5664
rect 25280 5652 25286 5704
rect 23309 5528 23888 5556
rect 26988 5556 27016 5800
rect 27065 5763 27123 5769
rect 27065 5729 27077 5763
rect 27111 5760 27123 5763
rect 27338 5760 27344 5772
rect 27111 5732 27344 5760
rect 27111 5729 27123 5732
rect 27065 5723 27123 5729
rect 27338 5720 27344 5732
rect 27396 5720 27402 5772
rect 28460 5678 28488 5868
rect 28810 5856 28816 5908
rect 28868 5856 28874 5908
rect 29086 5856 29092 5908
rect 29144 5856 29150 5908
rect 31205 5899 31263 5905
rect 31205 5865 31217 5899
rect 31251 5896 31263 5899
rect 31386 5896 31392 5908
rect 31251 5868 31392 5896
rect 31251 5865 31263 5868
rect 31205 5859 31263 5865
rect 31386 5856 31392 5868
rect 31444 5856 31450 5908
rect 32858 5856 32864 5908
rect 32916 5896 32922 5908
rect 33965 5899 34023 5905
rect 33965 5896 33977 5899
rect 32916 5868 33977 5896
rect 32916 5856 32922 5868
rect 33965 5865 33977 5868
rect 34011 5865 34023 5899
rect 33965 5859 34023 5865
rect 28828 5828 28856 5856
rect 28828 5800 29960 5828
rect 29932 5760 29960 5800
rect 30282 5788 30288 5840
rect 30340 5828 30346 5840
rect 30650 5828 30656 5840
rect 30340 5800 30656 5828
rect 30340 5788 30346 5800
rect 30650 5788 30656 5800
rect 30708 5788 30714 5840
rect 30837 5831 30895 5837
rect 30837 5797 30849 5831
rect 30883 5828 30895 5831
rect 32030 5828 32036 5840
rect 30883 5800 32036 5828
rect 30883 5797 30895 5800
rect 30837 5791 30895 5797
rect 32030 5788 32036 5800
rect 32088 5788 32094 5840
rect 33226 5788 33232 5840
rect 33284 5828 33290 5840
rect 33689 5831 33747 5837
rect 33689 5828 33701 5831
rect 33284 5800 33701 5828
rect 33284 5788 33290 5800
rect 33689 5797 33701 5800
rect 33735 5828 33747 5831
rect 34057 5831 34115 5837
rect 34057 5828 34069 5831
rect 33735 5800 34069 5828
rect 33735 5797 33747 5800
rect 33689 5791 33747 5797
rect 34057 5797 34069 5800
rect 34103 5828 34115 5831
rect 34146 5828 34152 5840
rect 34103 5800 34152 5828
rect 34103 5797 34115 5800
rect 34057 5791 34115 5797
rect 34146 5788 34152 5800
rect 34204 5788 34210 5840
rect 30742 5760 30748 5772
rect 29932 5732 30748 5760
rect 29638 5652 29644 5704
rect 29696 5692 29702 5704
rect 29932 5701 29960 5732
rect 30742 5720 30748 5732
rect 30800 5760 30806 5772
rect 30800 5732 30972 5760
rect 30800 5720 30806 5732
rect 29733 5695 29791 5701
rect 29733 5692 29745 5695
rect 29696 5664 29745 5692
rect 29696 5652 29702 5664
rect 29733 5661 29745 5664
rect 29779 5661 29791 5695
rect 29733 5655 29791 5661
rect 29917 5695 29975 5701
rect 29917 5661 29929 5695
rect 29963 5661 29975 5695
rect 29917 5655 29975 5661
rect 30190 5652 30196 5704
rect 30248 5652 30254 5704
rect 30374 5652 30380 5704
rect 30432 5652 30438 5704
rect 30469 5695 30527 5701
rect 30469 5661 30481 5695
rect 30515 5661 30527 5695
rect 30469 5655 30527 5661
rect 30561 5695 30619 5701
rect 30561 5661 30573 5695
rect 30607 5661 30619 5695
rect 30561 5655 30619 5661
rect 27341 5627 27399 5633
rect 27341 5593 27353 5627
rect 27387 5624 27399 5627
rect 27430 5624 27436 5636
rect 27387 5596 27436 5624
rect 27387 5593 27399 5596
rect 27341 5587 27399 5593
rect 27430 5584 27436 5596
rect 27488 5584 27494 5636
rect 28718 5584 28724 5636
rect 28776 5624 28782 5636
rect 29549 5627 29607 5633
rect 29549 5624 29561 5627
rect 28776 5596 29561 5624
rect 28776 5584 28782 5596
rect 29549 5593 29561 5596
rect 29595 5593 29607 5627
rect 29822 5624 29828 5636
rect 29549 5587 29607 5593
rect 29748 5596 29828 5624
rect 29273 5559 29331 5565
rect 29273 5556 29285 5559
rect 26988 5528 29285 5556
rect 29273 5525 29285 5528
rect 29319 5556 29331 5559
rect 29748 5556 29776 5596
rect 29822 5584 29828 5596
rect 29880 5584 29886 5636
rect 30006 5584 30012 5636
rect 30064 5633 30070 5636
rect 30064 5627 30093 5633
rect 30081 5624 30093 5627
rect 30484 5624 30512 5655
rect 30081 5596 30512 5624
rect 30081 5593 30093 5596
rect 30064 5587 30093 5593
rect 30064 5584 30070 5587
rect 29319 5528 29776 5556
rect 29319 5525 29331 5528
rect 29273 5519 29331 5525
rect 30190 5516 30196 5568
rect 30248 5556 30254 5568
rect 30576 5556 30604 5655
rect 30650 5652 30656 5704
rect 30708 5652 30714 5704
rect 30944 5701 30972 5732
rect 31018 5720 31024 5772
rect 31076 5720 31082 5772
rect 31662 5720 31668 5772
rect 31720 5760 31726 5772
rect 32582 5760 32588 5772
rect 31720 5732 32588 5760
rect 31720 5720 31726 5732
rect 32582 5720 32588 5732
rect 32640 5760 32646 5772
rect 33321 5763 33379 5769
rect 33321 5760 33333 5763
rect 32640 5732 33333 5760
rect 32640 5720 32646 5732
rect 33321 5729 33333 5732
rect 33367 5729 33379 5763
rect 33873 5763 33931 5769
rect 33873 5760 33885 5763
rect 33321 5723 33379 5729
rect 33520 5732 33885 5760
rect 30929 5695 30987 5701
rect 30929 5661 30941 5695
rect 30975 5661 30987 5695
rect 30929 5655 30987 5661
rect 31205 5695 31263 5701
rect 31205 5661 31217 5695
rect 31251 5692 31263 5695
rect 31478 5692 31484 5704
rect 31251 5664 31484 5692
rect 31251 5661 31263 5664
rect 31205 5655 31263 5661
rect 31478 5652 31484 5664
rect 31536 5652 31542 5704
rect 33520 5701 33548 5732
rect 33873 5729 33885 5732
rect 33919 5729 33931 5763
rect 33873 5723 33931 5729
rect 33505 5695 33563 5701
rect 33505 5692 33517 5695
rect 33152 5664 33517 5692
rect 33152 5636 33180 5664
rect 33505 5661 33517 5664
rect 33551 5661 33563 5695
rect 33505 5655 33563 5661
rect 33781 5695 33839 5701
rect 33781 5661 33793 5695
rect 33827 5661 33839 5695
rect 33781 5655 33839 5661
rect 34149 5695 34207 5701
rect 34149 5661 34161 5695
rect 34195 5692 34207 5695
rect 34333 5695 34391 5701
rect 34333 5692 34345 5695
rect 34195 5664 34345 5692
rect 34195 5661 34207 5664
rect 34149 5655 34207 5661
rect 34333 5661 34345 5664
rect 34379 5661 34391 5695
rect 34333 5655 34391 5661
rect 31294 5584 31300 5636
rect 31352 5624 31358 5636
rect 31352 5596 32628 5624
rect 31352 5584 31358 5596
rect 30248 5528 30604 5556
rect 31389 5559 31447 5565
rect 30248 5516 30254 5528
rect 31389 5525 31401 5559
rect 31435 5556 31447 5559
rect 32490 5556 32496 5568
rect 31435 5528 32496 5556
rect 31435 5525 31447 5528
rect 31389 5519 31447 5525
rect 32490 5516 32496 5528
rect 32548 5516 32554 5568
rect 32600 5556 32628 5596
rect 33134 5584 33140 5636
rect 33192 5584 33198 5636
rect 33796 5624 33824 5655
rect 33962 5624 33968 5636
rect 33796 5596 33968 5624
rect 33962 5584 33968 5596
rect 34020 5624 34026 5636
rect 34164 5624 34192 5655
rect 34422 5652 34428 5704
rect 34480 5652 34486 5704
rect 34020 5596 34192 5624
rect 34020 5584 34026 5596
rect 34606 5556 34612 5568
rect 32600 5528 34612 5556
rect 34606 5516 34612 5528
rect 34664 5516 34670 5568
rect 1104 5466 35328 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35328 5466
rect 1104 5392 35328 5414
rect 24026 5312 24032 5364
rect 24084 5352 24090 5364
rect 24762 5352 24768 5364
rect 24084 5324 24768 5352
rect 24084 5312 24090 5324
rect 24762 5312 24768 5324
rect 24820 5352 24826 5364
rect 26237 5355 26295 5361
rect 26237 5352 26249 5355
rect 24820 5324 26249 5352
rect 24820 5312 24826 5324
rect 26237 5321 26249 5324
rect 26283 5321 26295 5355
rect 26237 5315 26295 5321
rect 30374 5312 30380 5364
rect 30432 5352 30438 5364
rect 30469 5355 30527 5361
rect 30469 5352 30481 5355
rect 30432 5324 30481 5352
rect 30432 5312 30438 5324
rect 30469 5321 30481 5324
rect 30515 5321 30527 5355
rect 30469 5315 30527 5321
rect 33134 5312 33140 5364
rect 33192 5352 33198 5364
rect 33689 5355 33747 5361
rect 33689 5352 33701 5355
rect 33192 5324 33701 5352
rect 33192 5312 33198 5324
rect 33689 5321 33701 5324
rect 33735 5321 33747 5355
rect 33689 5315 33747 5321
rect 22278 5244 22284 5296
rect 22336 5284 22342 5296
rect 24854 5284 24860 5296
rect 22336 5256 24860 5284
rect 22336 5244 22342 5256
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1489 5219 1547 5225
rect 1489 5216 1501 5219
rect 1360 5188 1501 5216
rect 1360 5176 1366 5188
rect 1489 5185 1501 5188
rect 1535 5216 1547 5219
rect 1949 5219 2007 5225
rect 1949 5216 1961 5219
rect 1535 5188 1961 5216
rect 1535 5185 1547 5188
rect 1489 5179 1547 5185
rect 1949 5185 1961 5188
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 23566 5176 23572 5228
rect 23624 5176 23630 5228
rect 24026 5176 24032 5228
rect 24084 5176 24090 5228
rect 24504 5225 24532 5256
rect 24854 5244 24860 5256
rect 24912 5244 24918 5296
rect 26050 5284 26056 5296
rect 25990 5256 26056 5284
rect 26050 5244 26056 5256
rect 26108 5244 26114 5296
rect 24489 5219 24547 5225
rect 24489 5185 24501 5219
rect 24535 5185 24547 5219
rect 24489 5179 24547 5185
rect 30466 5176 30472 5228
rect 30524 5216 30530 5228
rect 30653 5219 30711 5225
rect 30653 5216 30665 5219
rect 30524 5188 30665 5216
rect 30524 5176 30530 5188
rect 30653 5185 30665 5188
rect 30699 5185 30711 5219
rect 30653 5179 30711 5185
rect 33962 5176 33968 5228
rect 34020 5176 34026 5228
rect 34146 5176 34152 5228
rect 34204 5216 34210 5228
rect 34241 5219 34299 5225
rect 34241 5216 34253 5219
rect 34204 5188 34253 5216
rect 34204 5176 34210 5188
rect 34241 5185 34253 5188
rect 34287 5185 34299 5219
rect 34241 5179 34299 5185
rect 34422 5176 34428 5228
rect 34480 5176 34486 5228
rect 34517 5219 34575 5225
rect 34517 5185 34529 5219
rect 34563 5185 34575 5219
rect 34517 5179 34575 5185
rect 23290 5108 23296 5160
rect 23348 5148 23354 5160
rect 23842 5148 23848 5160
rect 23348 5120 23848 5148
rect 23348 5108 23354 5120
rect 23842 5108 23848 5120
rect 23900 5108 23906 5160
rect 23934 5108 23940 5160
rect 23992 5108 23998 5160
rect 24765 5151 24823 5157
rect 24765 5148 24777 5151
rect 24412 5120 24777 5148
rect 24412 5089 24440 5120
rect 24765 5117 24777 5120
rect 24811 5117 24823 5151
rect 24765 5111 24823 5117
rect 30834 5108 30840 5160
rect 30892 5148 30898 5160
rect 30929 5151 30987 5157
rect 30929 5148 30941 5151
rect 30892 5120 30941 5148
rect 30892 5108 30898 5120
rect 30929 5117 30941 5120
rect 30975 5148 30987 5151
rect 31018 5148 31024 5160
rect 30975 5120 31024 5148
rect 30975 5117 30987 5120
rect 30929 5111 30987 5117
rect 31018 5108 31024 5120
rect 31076 5108 31082 5160
rect 34333 5151 34391 5157
rect 34333 5117 34345 5151
rect 34379 5148 34391 5151
rect 34532 5148 34560 5179
rect 34379 5120 34560 5148
rect 34793 5151 34851 5157
rect 34379 5117 34391 5120
rect 34333 5111 34391 5117
rect 34793 5117 34805 5151
rect 34839 5148 34851 5151
rect 35342 5148 35348 5160
rect 34839 5120 35348 5148
rect 34839 5117 34851 5120
rect 34793 5111 34851 5117
rect 35342 5108 35348 5120
rect 35400 5108 35406 5160
rect 24397 5083 24455 5089
rect 24397 5049 24409 5083
rect 24443 5049 24455 5083
rect 24397 5043 24455 5049
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 1854 5012 1860 5024
rect 1627 4984 1860 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 1854 4972 1860 4984
rect 1912 4972 1918 5024
rect 30742 4972 30748 5024
rect 30800 5012 30806 5024
rect 30837 5015 30895 5021
rect 30837 5012 30849 5015
rect 30800 4984 30849 5012
rect 30800 4972 30806 4984
rect 30837 4981 30849 4984
rect 30883 4981 30895 5015
rect 30837 4975 30895 4981
rect 34054 4972 34060 5024
rect 34112 5012 34118 5024
rect 34149 5015 34207 5021
rect 34149 5012 34161 5015
rect 34112 4984 34161 5012
rect 34112 4972 34118 4984
rect 34149 4981 34161 4984
rect 34195 4981 34207 5015
rect 34149 4975 34207 4981
rect 1104 4922 35328 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 35328 4922
rect 1104 4848 35328 4870
rect 1854 4768 1860 4820
rect 1912 4808 1918 4820
rect 33134 4808 33140 4820
rect 1912 4780 33140 4808
rect 1912 4768 1918 4780
rect 33134 4768 33140 4780
rect 33192 4768 33198 4820
rect 31757 4743 31815 4749
rect 31757 4709 31769 4743
rect 31803 4709 31815 4743
rect 31757 4703 31815 4709
rect 22278 4632 22284 4684
rect 22336 4672 22342 4684
rect 22465 4675 22523 4681
rect 22465 4672 22477 4675
rect 22336 4644 22477 4672
rect 22336 4632 22342 4644
rect 22465 4641 22477 4644
rect 22511 4641 22523 4675
rect 22465 4635 22523 4641
rect 23474 4632 23480 4684
rect 23532 4672 23538 4684
rect 23532 4644 23980 4672
rect 23532 4632 23538 4644
rect 22738 4496 22744 4548
rect 22796 4496 22802 4548
rect 23952 4536 23980 4644
rect 28994 4632 29000 4684
rect 29052 4672 29058 4684
rect 30282 4672 30288 4684
rect 29052 4644 30288 4672
rect 29052 4632 29058 4644
rect 30282 4632 30288 4644
rect 30340 4632 30346 4684
rect 30466 4632 30472 4684
rect 30524 4672 30530 4684
rect 30561 4675 30619 4681
rect 30561 4672 30573 4675
rect 30524 4644 30573 4672
rect 30524 4632 30530 4644
rect 30561 4641 30573 4644
rect 30607 4672 30619 4675
rect 31297 4675 31355 4681
rect 31297 4672 31309 4675
rect 30607 4644 31309 4672
rect 30607 4641 30619 4644
rect 30561 4635 30619 4641
rect 31297 4641 31309 4644
rect 31343 4641 31355 4675
rect 31772 4672 31800 4703
rect 32398 4700 32404 4752
rect 32456 4700 32462 4752
rect 31941 4675 31999 4681
rect 31941 4672 31953 4675
rect 31772 4644 31953 4672
rect 31297 4635 31355 4641
rect 31941 4641 31953 4644
rect 31987 4641 31999 4675
rect 31941 4635 31999 4641
rect 30653 4607 30711 4613
rect 30653 4573 30665 4607
rect 30699 4604 30711 4607
rect 30834 4604 30840 4616
rect 30699 4576 30840 4604
rect 30699 4573 30711 4576
rect 30653 4567 30711 4573
rect 30834 4564 30840 4576
rect 30892 4564 30898 4616
rect 31386 4564 31392 4616
rect 31444 4564 31450 4616
rect 32030 4564 32036 4616
rect 32088 4564 32094 4616
rect 32677 4607 32735 4613
rect 32677 4573 32689 4607
rect 32723 4573 32735 4607
rect 32677 4567 32735 4573
rect 24394 4536 24400 4548
rect 23952 4522 24400 4536
rect 23966 4508 24400 4522
rect 24394 4496 24400 4508
rect 24452 4496 24458 4548
rect 29086 4496 29092 4548
rect 29144 4536 29150 4548
rect 29914 4536 29920 4548
rect 29144 4508 29920 4536
rect 29144 4496 29150 4508
rect 29914 4496 29920 4508
rect 29972 4536 29978 4548
rect 32692 4536 32720 4567
rect 29972 4508 32720 4536
rect 32953 4539 33011 4545
rect 29972 4496 29978 4508
rect 32953 4505 32965 4539
rect 32999 4536 33011 4539
rect 33226 4536 33232 4548
rect 32999 4508 33232 4536
rect 32999 4505 33011 4508
rect 32953 4499 33011 4505
rect 33226 4496 33232 4508
rect 33284 4496 33290 4548
rect 33336 4508 33442 4536
rect 23566 4428 23572 4480
rect 23624 4468 23630 4480
rect 24213 4471 24271 4477
rect 24213 4468 24225 4471
rect 23624 4440 24225 4468
rect 23624 4428 23630 4440
rect 24213 4437 24225 4440
rect 24259 4437 24271 4471
rect 24213 4431 24271 4437
rect 31110 4428 31116 4480
rect 31168 4468 31174 4480
rect 33336 4468 33364 4508
rect 31168 4440 33364 4468
rect 31168 4428 31174 4440
rect 34422 4428 34428 4480
rect 34480 4428 34486 4480
rect 1104 4378 35328 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35328 4378
rect 1104 4304 35328 4326
rect 22465 4267 22523 4273
rect 22465 4233 22477 4267
rect 22511 4264 22523 4267
rect 22738 4264 22744 4276
rect 22511 4236 22744 4264
rect 22511 4233 22523 4236
rect 22465 4227 22523 4233
rect 22738 4224 22744 4236
rect 22796 4224 22802 4276
rect 31110 4224 31116 4276
rect 31168 4224 31174 4276
rect 32398 4224 32404 4276
rect 32456 4264 32462 4276
rect 32769 4267 32827 4273
rect 32769 4264 32781 4267
rect 32456 4236 32781 4264
rect 32456 4224 32462 4236
rect 32769 4233 32781 4236
rect 32815 4233 32827 4267
rect 32769 4227 32827 4233
rect 33226 4224 33232 4276
rect 33284 4224 33290 4276
rect 31128 4196 31156 4224
rect 31294 4196 31300 4208
rect 30590 4168 31156 4196
rect 31220 4168 31300 4196
rect 22833 4131 22891 4137
rect 22833 4097 22845 4131
rect 22879 4128 22891 4131
rect 23290 4128 23296 4140
rect 22879 4100 23296 4128
rect 22879 4097 22891 4100
rect 22833 4091 22891 4097
rect 23290 4088 23296 4100
rect 23348 4088 23354 4140
rect 28629 4131 28687 4137
rect 28629 4097 28641 4131
rect 28675 4128 28687 4131
rect 28994 4128 29000 4140
rect 28675 4100 29000 4128
rect 28675 4097 28687 4100
rect 28629 4091 28687 4097
rect 28994 4088 29000 4100
rect 29052 4088 29058 4140
rect 29086 4088 29092 4140
rect 29144 4088 29150 4140
rect 30944 4137 30972 4168
rect 30929 4131 30987 4137
rect 30929 4097 30941 4131
rect 30975 4128 30987 4131
rect 31113 4131 31171 4137
rect 30975 4100 31009 4128
rect 30975 4097 30987 4100
rect 30929 4091 30987 4097
rect 31113 4097 31125 4131
rect 31159 4128 31171 4131
rect 31220 4128 31248 4168
rect 31294 4156 31300 4168
rect 31352 4156 31358 4208
rect 31386 4156 31392 4208
rect 31444 4196 31450 4208
rect 32861 4199 32919 4205
rect 32861 4196 32873 4199
rect 31444 4168 32873 4196
rect 31444 4156 31450 4168
rect 32861 4165 32873 4168
rect 32907 4196 32919 4199
rect 34422 4196 34428 4208
rect 32907 4168 34428 4196
rect 32907 4165 32919 4168
rect 32861 4159 32919 4165
rect 34422 4156 34428 4168
rect 34480 4156 34486 4208
rect 31159 4100 31248 4128
rect 31159 4097 31171 4100
rect 31113 4091 31171 4097
rect 22925 4063 22983 4069
rect 22925 4029 22937 4063
rect 22971 4060 22983 4063
rect 23198 4060 23204 4072
rect 22971 4032 23204 4060
rect 22971 4029 22983 4032
rect 22925 4023 22983 4029
rect 23198 4020 23204 4032
rect 23256 4020 23262 4072
rect 28718 4020 28724 4072
rect 28776 4020 28782 4072
rect 29365 4063 29423 4069
rect 29365 4029 29377 4063
rect 29411 4060 29423 4063
rect 29822 4060 29828 4072
rect 29411 4032 29828 4060
rect 29411 4029 29423 4032
rect 29365 4023 29423 4029
rect 29822 4020 29828 4032
rect 29880 4020 29886 4072
rect 30098 4020 30104 4072
rect 30156 4060 30162 4072
rect 32585 4063 32643 4069
rect 32585 4060 32597 4063
rect 30156 4032 32597 4060
rect 30156 4020 30162 4032
rect 32585 4029 32597 4032
rect 32631 4029 32643 4063
rect 32585 4023 32643 4029
rect 28994 3884 29000 3936
rect 29052 3884 29058 3936
rect 30834 3884 30840 3936
rect 30892 3884 30898 3936
rect 1104 3834 35328 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 35328 3834
rect 1104 3760 35328 3782
rect 29822 3680 29828 3732
rect 29880 3680 29886 3732
rect 30098 3612 30104 3664
rect 30156 3652 30162 3664
rect 30156 3624 30420 3652
rect 30156 3612 30162 3624
rect 28994 3544 29000 3596
rect 29052 3584 29058 3596
rect 30392 3593 30420 3624
rect 30285 3587 30343 3593
rect 30285 3584 30297 3587
rect 29052 3556 30297 3584
rect 29052 3544 29058 3556
rect 30285 3553 30297 3556
rect 30331 3553 30343 3587
rect 30285 3547 30343 3553
rect 30377 3587 30435 3593
rect 30377 3553 30389 3587
rect 30423 3553 30435 3587
rect 30377 3547 30435 3553
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 1360 3488 1409 3516
rect 1360 3476 1366 3488
rect 1397 3485 1409 3488
rect 1443 3516 1455 3519
rect 1857 3519 1915 3525
rect 1857 3516 1869 3519
rect 1443 3488 1869 3516
rect 1443 3485 1455 3488
rect 1397 3479 1455 3485
rect 1857 3485 1869 3488
rect 1903 3485 1915 3519
rect 1857 3479 1915 3485
rect 30193 3519 30251 3525
rect 30193 3485 30205 3519
rect 30239 3516 30251 3519
rect 30834 3516 30840 3528
rect 30239 3488 30840 3516
rect 30239 3485 30251 3488
rect 30193 3479 30251 3485
rect 30834 3476 30840 3488
rect 30892 3476 30898 3528
rect 34054 3476 34060 3528
rect 34112 3476 34118 3528
rect 1765 3451 1823 3457
rect 1765 3448 1777 3451
rect 1596 3420 1777 3448
rect 1596 3389 1624 3420
rect 1765 3417 1777 3420
rect 1811 3448 1823 3451
rect 1811 3420 2774 3448
rect 1811 3417 1823 3420
rect 1765 3411 1823 3417
rect 1581 3383 1639 3389
rect 1581 3349 1593 3383
rect 1627 3349 1639 3383
rect 2746 3380 2774 3420
rect 34330 3408 34336 3460
rect 34388 3408 34394 3460
rect 21542 3380 21548 3392
rect 2746 3352 21548 3380
rect 1581 3343 1639 3349
rect 21542 3340 21548 3352
rect 21600 3340 21606 3392
rect 1104 3290 35328 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35328 3290
rect 1104 3216 35328 3238
rect 1104 2746 35328 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 35328 2746
rect 1104 2672 35328 2694
rect 1104 2202 35328 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35328 2202
rect 1104 2128 35328 2150
<< via1 >>
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 1216 35708 1268 35760
rect 1308 35640 1360 35692
rect 19708 35708 19760 35760
rect 10968 35640 11020 35692
rect 12072 35572 12124 35624
rect 3608 35504 3660 35556
rect 11336 35436 11388 35488
rect 14004 35436 14056 35488
rect 18880 35436 18932 35488
rect 25688 35683 25740 35692
rect 25688 35649 25697 35683
rect 25697 35649 25731 35683
rect 25731 35649 25740 35683
rect 25688 35640 25740 35649
rect 28724 35640 28776 35692
rect 34520 35683 34572 35692
rect 34520 35649 34529 35683
rect 34529 35649 34563 35683
rect 34563 35649 34572 35683
rect 34520 35640 34572 35649
rect 19064 35572 19116 35624
rect 25596 35615 25648 35624
rect 25596 35581 25605 35615
rect 25605 35581 25639 35615
rect 25639 35581 25648 35615
rect 25596 35572 25648 35581
rect 27988 35615 28040 35624
rect 27988 35581 27997 35615
rect 27997 35581 28031 35615
rect 28031 35581 28040 35615
rect 27988 35572 28040 35581
rect 34336 35615 34388 35624
rect 34336 35581 34345 35615
rect 34345 35581 34379 35615
rect 34379 35581 34388 35615
rect 34336 35572 34388 35581
rect 19156 35436 19208 35488
rect 19248 35479 19300 35488
rect 19248 35445 19257 35479
rect 19257 35445 19291 35479
rect 19291 35445 19300 35479
rect 19248 35436 19300 35445
rect 26056 35479 26108 35488
rect 26056 35445 26065 35479
rect 26065 35445 26099 35479
rect 26099 35445 26108 35479
rect 26056 35436 26108 35445
rect 26240 35479 26292 35488
rect 26240 35445 26249 35479
rect 26249 35445 26283 35479
rect 26283 35445 26292 35479
rect 26240 35436 26292 35445
rect 27436 35479 27488 35488
rect 27436 35445 27445 35479
rect 27445 35445 27479 35479
rect 27479 35445 27488 35479
rect 27436 35436 27488 35445
rect 27620 35436 27672 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 1308 35232 1360 35284
rect 9036 35232 9088 35284
rect 17224 35232 17276 35284
rect 19064 35275 19116 35284
rect 19064 35241 19073 35275
rect 19073 35241 19107 35275
rect 19107 35241 19116 35275
rect 19064 35232 19116 35241
rect 19156 35232 19208 35284
rect 25596 35232 25648 35284
rect 27988 35232 28040 35284
rect 28448 35232 28500 35284
rect 28724 35275 28776 35284
rect 28724 35241 28733 35275
rect 28733 35241 28767 35275
rect 28767 35241 28776 35275
rect 28724 35232 28776 35241
rect 14004 35096 14056 35148
rect 7104 35028 7156 35080
rect 11888 35028 11940 35080
rect 15108 35071 15160 35080
rect 15108 35037 15117 35071
rect 15117 35037 15151 35071
rect 15151 35037 15160 35071
rect 15108 35028 15160 35037
rect 17408 35028 17460 35080
rect 19248 35028 19300 35080
rect 22192 35071 22244 35080
rect 22192 35037 22201 35071
rect 22201 35037 22235 35071
rect 22235 35037 22244 35071
rect 22192 35028 22244 35037
rect 26056 35028 26108 35080
rect 27252 35071 27304 35080
rect 27252 35037 27261 35071
rect 27261 35037 27295 35071
rect 27295 35037 27304 35071
rect 27252 35028 27304 35037
rect 27620 35071 27672 35080
rect 27620 35037 27654 35071
rect 27654 35037 27672 35071
rect 27620 35028 27672 35037
rect 8116 34960 8168 35012
rect 9588 34960 9640 35012
rect 11336 35003 11388 35012
rect 11336 34969 11370 35003
rect 11370 34969 11388 35003
rect 11336 34960 11388 34969
rect 11520 34960 11572 35012
rect 15568 34960 15620 35012
rect 20168 34960 20220 35012
rect 23296 34960 23348 35012
rect 24676 35003 24728 35012
rect 24676 34969 24710 35003
rect 24710 34969 24728 35003
rect 24676 34960 24728 34969
rect 8760 34935 8812 34944
rect 8760 34901 8769 34935
rect 8769 34901 8803 34935
rect 8803 34901 8812 34935
rect 8760 34892 8812 34901
rect 10876 34935 10928 34944
rect 10876 34901 10885 34935
rect 10885 34901 10919 34935
rect 10919 34901 10928 34935
rect 10876 34892 10928 34901
rect 10968 34892 11020 34944
rect 13636 34935 13688 34944
rect 13636 34901 13645 34935
rect 13645 34901 13679 34935
rect 13679 34901 13688 34935
rect 13636 34892 13688 34901
rect 13728 34892 13780 34944
rect 14464 34935 14516 34944
rect 14464 34901 14473 34935
rect 14473 34901 14507 34935
rect 14507 34901 14516 34935
rect 14464 34892 14516 34901
rect 16028 34892 16080 34944
rect 20996 34935 21048 34944
rect 20996 34901 21005 34935
rect 21005 34901 21039 34935
rect 21039 34901 21048 34935
rect 20996 34892 21048 34901
rect 23572 34935 23624 34944
rect 23572 34901 23581 34935
rect 23581 34901 23615 34935
rect 23615 34901 23624 34935
rect 23572 34892 23624 34901
rect 25780 34935 25832 34944
rect 25780 34901 25789 34935
rect 25789 34901 25823 34935
rect 25823 34901 25832 34935
rect 25780 34892 25832 34901
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 8116 34731 8168 34740
rect 8116 34697 8125 34731
rect 8125 34697 8159 34731
rect 8159 34697 8168 34731
rect 8116 34688 8168 34697
rect 9036 34731 9088 34740
rect 9036 34697 9045 34731
rect 9045 34697 9079 34731
rect 9079 34697 9088 34731
rect 9036 34688 9088 34697
rect 9588 34731 9640 34740
rect 9588 34697 9597 34731
rect 9597 34697 9631 34731
rect 9631 34697 9640 34731
rect 9588 34688 9640 34697
rect 10600 34688 10652 34740
rect 10876 34688 10928 34740
rect 14464 34688 14516 34740
rect 15568 34731 15620 34740
rect 15568 34697 15577 34731
rect 15577 34697 15611 34731
rect 15611 34697 15620 34731
rect 15568 34688 15620 34697
rect 16028 34731 16080 34740
rect 16028 34697 16037 34731
rect 16037 34697 16071 34731
rect 16071 34697 16080 34731
rect 16028 34688 16080 34697
rect 20168 34731 20220 34740
rect 20168 34697 20177 34731
rect 20177 34697 20211 34731
rect 20211 34697 20220 34731
rect 20168 34688 20220 34697
rect 20720 34688 20772 34740
rect 20996 34688 21048 34740
rect 10416 34620 10468 34672
rect 8760 34552 8812 34604
rect 9680 34552 9732 34604
rect 12072 34552 12124 34604
rect 13176 34552 13228 34604
rect 14096 34620 14148 34672
rect 15108 34620 15160 34672
rect 17224 34620 17276 34672
rect 13728 34595 13780 34604
rect 13728 34561 13762 34595
rect 13762 34561 13780 34595
rect 13728 34552 13780 34561
rect 9036 34484 9088 34536
rect 9404 34484 9456 34536
rect 10416 34527 10468 34536
rect 10416 34493 10425 34527
rect 10425 34493 10459 34527
rect 10459 34493 10468 34527
rect 10416 34484 10468 34493
rect 11520 34484 11572 34536
rect 10324 34416 10376 34468
rect 11612 34459 11664 34468
rect 11612 34425 11621 34459
rect 11621 34425 11655 34459
rect 11655 34425 11664 34459
rect 11612 34416 11664 34425
rect 13360 34391 13412 34400
rect 13360 34357 13369 34391
rect 13369 34357 13403 34391
rect 13403 34357 13412 34391
rect 13360 34348 13412 34357
rect 13636 34348 13688 34400
rect 18328 34595 18380 34604
rect 18328 34561 18337 34595
rect 18337 34561 18371 34595
rect 18371 34561 18380 34595
rect 18328 34552 18380 34561
rect 22192 34620 22244 34672
rect 22560 34620 22612 34672
rect 23296 34731 23348 34740
rect 23296 34697 23305 34731
rect 23305 34697 23339 34731
rect 23339 34697 23348 34731
rect 23296 34688 23348 34697
rect 23572 34688 23624 34740
rect 24676 34688 24728 34740
rect 25320 34688 25372 34740
rect 25780 34688 25832 34740
rect 27988 34688 28040 34740
rect 22100 34595 22152 34604
rect 22100 34561 22134 34595
rect 22134 34561 22152 34595
rect 22100 34552 22152 34561
rect 23756 34595 23808 34604
rect 23756 34561 23765 34595
rect 23765 34561 23799 34595
rect 23799 34561 23808 34595
rect 23756 34552 23808 34561
rect 16212 34527 16264 34536
rect 16212 34493 16221 34527
rect 16221 34493 16255 34527
rect 16255 34493 16264 34527
rect 16212 34484 16264 34493
rect 18420 34527 18472 34536
rect 18420 34493 18429 34527
rect 18429 34493 18463 34527
rect 18463 34493 18472 34527
rect 18420 34484 18472 34493
rect 18880 34484 18932 34536
rect 19708 34484 19760 34536
rect 20812 34527 20864 34536
rect 20812 34493 20821 34527
rect 20821 34493 20855 34527
rect 20855 34493 20864 34527
rect 20812 34484 20864 34493
rect 16120 34348 16172 34400
rect 17684 34348 17736 34400
rect 22468 34348 22520 34400
rect 28080 34595 28132 34604
rect 28080 34561 28089 34595
rect 28089 34561 28123 34595
rect 28123 34561 28132 34595
rect 28080 34552 28132 34561
rect 27804 34416 27856 34468
rect 23204 34391 23256 34400
rect 23204 34357 23213 34391
rect 23213 34357 23247 34391
rect 23247 34357 23256 34391
rect 23204 34348 23256 34357
rect 27620 34348 27672 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 13176 34187 13228 34196
rect 13176 34153 13185 34187
rect 13185 34153 13219 34187
rect 13219 34153 13228 34187
rect 13176 34144 13228 34153
rect 13452 34144 13504 34196
rect 14740 34144 14792 34196
rect 18328 34144 18380 34196
rect 18788 34187 18840 34196
rect 18788 34153 18797 34187
rect 18797 34153 18831 34187
rect 18831 34153 18840 34187
rect 18788 34144 18840 34153
rect 22100 34187 22152 34196
rect 22100 34153 22109 34187
rect 22109 34153 22143 34187
rect 22143 34153 22152 34187
rect 22100 34144 22152 34153
rect 25780 34144 25832 34196
rect 26332 34144 26384 34196
rect 28080 34144 28132 34196
rect 28632 34144 28684 34196
rect 4804 34008 4856 34060
rect 1308 33940 1360 33992
rect 3608 33940 3660 33992
rect 5908 33940 5960 33992
rect 7104 33940 7156 33992
rect 10232 33940 10284 33992
rect 10600 33983 10652 33992
rect 10600 33949 10610 33983
rect 10610 33949 10644 33983
rect 10644 33949 10652 33983
rect 16304 34076 16356 34128
rect 18420 34076 18472 34128
rect 19248 34076 19300 34128
rect 13728 34051 13780 34060
rect 13728 34017 13737 34051
rect 13737 34017 13771 34051
rect 13771 34017 13780 34051
rect 13728 34008 13780 34017
rect 17224 34008 17276 34060
rect 23756 34076 23808 34128
rect 23296 34008 23348 34060
rect 10600 33940 10652 33949
rect 7380 33872 7432 33924
rect 4068 33804 4120 33856
rect 6368 33804 6420 33856
rect 9036 33872 9088 33924
rect 9220 33915 9272 33924
rect 9220 33881 9254 33915
rect 9254 33881 9272 33915
rect 9220 33872 9272 33881
rect 10876 33915 10928 33924
rect 10876 33881 10885 33915
rect 10885 33881 10919 33915
rect 10919 33881 10928 33915
rect 10876 33872 10928 33881
rect 13360 33940 13412 33992
rect 14464 33940 14516 33992
rect 14740 33983 14792 33992
rect 14740 33949 14749 33983
rect 14749 33949 14783 33983
rect 14783 33949 14792 33983
rect 14740 33940 14792 33949
rect 15292 33940 15344 33992
rect 16488 33940 16540 33992
rect 16672 33940 16724 33992
rect 17408 33983 17460 33992
rect 17408 33949 17417 33983
rect 17417 33949 17451 33983
rect 17451 33949 17460 33983
rect 17408 33940 17460 33949
rect 17684 33983 17736 33992
rect 17684 33949 17718 33983
rect 17718 33949 17736 33983
rect 17684 33940 17736 33949
rect 18880 33983 18932 33992
rect 18880 33949 18889 33983
rect 18889 33949 18923 33983
rect 18923 33949 18932 33983
rect 18880 33940 18932 33949
rect 20904 33940 20956 33992
rect 23204 33983 23256 33992
rect 23204 33949 23213 33983
rect 23213 33949 23247 33983
rect 23247 33949 23256 33983
rect 23204 33940 23256 33949
rect 13452 33872 13504 33924
rect 14556 33915 14608 33924
rect 14556 33881 14565 33915
rect 14565 33881 14599 33915
rect 14599 33881 14608 33915
rect 14556 33872 14608 33881
rect 15660 33872 15712 33924
rect 16304 33872 16356 33924
rect 7656 33847 7708 33856
rect 7656 33813 7665 33847
rect 7665 33813 7699 33847
rect 7699 33813 7708 33847
rect 7656 33804 7708 33813
rect 9956 33804 10008 33856
rect 11152 33847 11204 33856
rect 11152 33813 11161 33847
rect 11161 33813 11195 33847
rect 11195 33813 11204 33847
rect 11152 33804 11204 33813
rect 13636 33847 13688 33856
rect 13636 33813 13645 33847
rect 13645 33813 13679 33847
rect 13679 33813 13688 33847
rect 13636 33804 13688 33813
rect 14924 33847 14976 33856
rect 14924 33813 14933 33847
rect 14933 33813 14967 33847
rect 14967 33813 14976 33847
rect 14924 33804 14976 33813
rect 15384 33804 15436 33856
rect 16580 33804 16632 33856
rect 17316 33804 17368 33856
rect 17592 33872 17644 33924
rect 23480 33983 23532 33992
rect 23480 33949 23489 33983
rect 23489 33949 23523 33983
rect 23523 33949 23532 33983
rect 23480 33940 23532 33949
rect 23848 33940 23900 33992
rect 25320 33983 25372 33992
rect 25320 33949 25329 33983
rect 25329 33949 25363 33983
rect 25363 33949 25372 33983
rect 25320 33940 25372 33949
rect 25596 33983 25648 33992
rect 25596 33949 25605 33983
rect 25605 33949 25639 33983
rect 25639 33949 25648 33983
rect 25596 33940 25648 33949
rect 25780 33940 25832 33992
rect 23664 33872 23716 33924
rect 20812 33804 20864 33856
rect 22928 33804 22980 33856
rect 23296 33804 23348 33856
rect 26424 33872 26476 33924
rect 26792 33940 26844 33992
rect 27252 33940 27304 33992
rect 27620 33983 27672 33992
rect 27620 33949 27654 33983
rect 27654 33949 27672 33983
rect 27620 33940 27672 33949
rect 23848 33847 23900 33856
rect 23848 33813 23857 33847
rect 23857 33813 23891 33847
rect 23891 33813 23900 33847
rect 23848 33804 23900 33813
rect 24124 33847 24176 33856
rect 24124 33813 24133 33847
rect 24133 33813 24167 33847
rect 24167 33813 24176 33847
rect 24124 33804 24176 33813
rect 25872 33847 25924 33856
rect 25872 33813 25881 33847
rect 25881 33813 25915 33847
rect 25915 33813 25924 33847
rect 25872 33804 25924 33813
rect 34060 33983 34112 33992
rect 34060 33949 34069 33983
rect 34069 33949 34103 33983
rect 34103 33949 34112 33983
rect 34060 33940 34112 33949
rect 34336 33915 34388 33924
rect 34336 33881 34345 33915
rect 34345 33881 34379 33915
rect 34379 33881 34388 33915
rect 34336 33872 34388 33881
rect 29184 33804 29236 33856
rect 32864 33847 32916 33856
rect 32864 33813 32873 33847
rect 32873 33813 32907 33847
rect 32907 33813 32916 33847
rect 32864 33804 32916 33813
rect 34428 33804 34480 33856
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 7380 33643 7432 33652
rect 7380 33609 7389 33643
rect 7389 33609 7423 33643
rect 7423 33609 7432 33643
rect 7380 33600 7432 33609
rect 7656 33600 7708 33652
rect 9220 33600 9272 33652
rect 10232 33643 10284 33652
rect 10232 33609 10241 33643
rect 10241 33609 10275 33643
rect 10275 33609 10284 33643
rect 10232 33600 10284 33609
rect 10508 33600 10560 33652
rect 7104 33575 7156 33584
rect 7104 33541 7113 33575
rect 7113 33541 7147 33575
rect 7147 33541 7156 33575
rect 7104 33532 7156 33541
rect 5448 33464 5500 33516
rect 6368 33507 6420 33516
rect 6368 33473 6377 33507
rect 6377 33473 6411 33507
rect 6411 33473 6420 33507
rect 6368 33464 6420 33473
rect 9680 33507 9732 33516
rect 9680 33473 9689 33507
rect 9689 33473 9723 33507
rect 9723 33473 9732 33507
rect 9680 33464 9732 33473
rect 9864 33575 9916 33584
rect 9864 33541 9873 33575
rect 9873 33541 9907 33575
rect 9907 33541 9916 33575
rect 9864 33532 9916 33541
rect 9956 33575 10008 33584
rect 9956 33541 9965 33575
rect 9965 33541 9999 33575
rect 9999 33541 10008 33575
rect 9956 33532 10008 33541
rect 14556 33600 14608 33652
rect 16304 33600 16356 33652
rect 4804 33439 4856 33448
rect 4804 33405 4813 33439
rect 4813 33405 4847 33439
rect 4847 33405 4856 33439
rect 4804 33396 4856 33405
rect 7840 33439 7892 33448
rect 7840 33405 7849 33439
rect 7849 33405 7883 33439
rect 7883 33405 7892 33439
rect 7840 33396 7892 33405
rect 6184 33303 6236 33312
rect 6184 33269 6193 33303
rect 6193 33269 6227 33303
rect 6227 33269 6236 33303
rect 6184 33260 6236 33269
rect 9772 33396 9824 33448
rect 9220 33328 9272 33380
rect 10048 33507 10100 33516
rect 10048 33473 10057 33507
rect 10057 33473 10091 33507
rect 10091 33473 10100 33507
rect 10048 33464 10100 33473
rect 9956 33328 10008 33380
rect 10048 33328 10100 33380
rect 11796 33507 11848 33516
rect 11796 33473 11830 33507
rect 11830 33473 11848 33507
rect 11796 33464 11848 33473
rect 11520 33439 11572 33448
rect 11520 33405 11529 33439
rect 11529 33405 11563 33439
rect 11563 33405 11572 33439
rect 11520 33396 11572 33405
rect 16028 33532 16080 33584
rect 16120 33575 16172 33584
rect 16120 33541 16129 33575
rect 16129 33541 16163 33575
rect 16163 33541 16172 33575
rect 16120 33532 16172 33541
rect 17040 33532 17092 33584
rect 19064 33575 19116 33584
rect 19064 33541 19073 33575
rect 19073 33541 19107 33575
rect 19107 33541 19116 33575
rect 19064 33532 19116 33541
rect 14924 33464 14976 33516
rect 15108 33507 15160 33516
rect 15108 33473 15118 33507
rect 15118 33473 15152 33507
rect 15152 33473 15160 33507
rect 15108 33464 15160 33473
rect 15660 33464 15712 33516
rect 15384 33396 15436 33448
rect 15844 33328 15896 33380
rect 16672 33439 16724 33448
rect 16672 33405 16681 33439
rect 16681 33405 16715 33439
rect 16715 33405 16724 33439
rect 16672 33396 16724 33405
rect 16580 33328 16632 33380
rect 18696 33507 18748 33516
rect 18696 33473 18705 33507
rect 18705 33473 18739 33507
rect 18739 33473 18748 33507
rect 18696 33464 18748 33473
rect 18788 33507 18840 33516
rect 18788 33473 18798 33507
rect 18798 33473 18832 33507
rect 18832 33473 18840 33507
rect 18788 33464 18840 33473
rect 25780 33600 25832 33652
rect 19616 33532 19668 33584
rect 22008 33532 22060 33584
rect 20444 33507 20496 33516
rect 20444 33473 20453 33507
rect 20453 33473 20487 33507
rect 20487 33473 20496 33507
rect 20444 33464 20496 33473
rect 20720 33507 20772 33516
rect 20720 33473 20729 33507
rect 20729 33473 20763 33507
rect 20763 33473 20772 33507
rect 20720 33464 20772 33473
rect 20812 33507 20864 33516
rect 20812 33473 20821 33507
rect 20821 33473 20855 33507
rect 20855 33473 20864 33507
rect 20812 33464 20864 33473
rect 20996 33464 21048 33516
rect 17776 33328 17828 33380
rect 23112 33464 23164 33516
rect 27528 33532 27580 33584
rect 28632 33575 28684 33584
rect 28632 33541 28641 33575
rect 28641 33541 28675 33575
rect 28675 33541 28684 33575
rect 28632 33532 28684 33541
rect 22560 33396 22612 33448
rect 26792 33439 26844 33448
rect 26792 33405 26801 33439
rect 26801 33405 26835 33439
rect 26835 33405 26844 33439
rect 26792 33396 26844 33405
rect 12164 33260 12216 33312
rect 17408 33260 17460 33312
rect 21088 33303 21140 33312
rect 21088 33269 21097 33303
rect 21097 33269 21131 33303
rect 21131 33269 21140 33303
rect 21088 33260 21140 33269
rect 23112 33303 23164 33312
rect 23112 33269 23121 33303
rect 23121 33269 23155 33303
rect 23155 33269 23164 33303
rect 23112 33260 23164 33269
rect 26608 33260 26660 33312
rect 28264 33507 28316 33516
rect 28264 33473 28273 33507
rect 28273 33473 28307 33507
rect 28307 33473 28316 33507
rect 28264 33464 28316 33473
rect 28448 33507 28500 33516
rect 28448 33473 28455 33507
rect 28455 33473 28500 33507
rect 28448 33464 28500 33473
rect 27712 33396 27764 33448
rect 28724 33507 28776 33516
rect 28724 33473 28738 33507
rect 28738 33473 28772 33507
rect 28772 33473 28776 33507
rect 28724 33464 28776 33473
rect 29276 33507 29328 33516
rect 29276 33473 29285 33507
rect 29285 33473 29319 33507
rect 29319 33473 29328 33507
rect 29276 33464 29328 33473
rect 34520 33600 34572 33652
rect 29828 33507 29880 33516
rect 29828 33473 29837 33507
rect 29837 33473 29871 33507
rect 29871 33473 29880 33507
rect 29828 33464 29880 33473
rect 33508 33464 33560 33516
rect 34152 33507 34204 33516
rect 34152 33473 34161 33507
rect 34161 33473 34195 33507
rect 34195 33473 34204 33507
rect 34152 33464 34204 33473
rect 34428 33507 34480 33516
rect 34428 33473 34437 33507
rect 34437 33473 34471 33507
rect 34471 33473 34480 33507
rect 34428 33464 34480 33473
rect 29552 33328 29604 33380
rect 32128 33439 32180 33448
rect 32128 33405 32137 33439
rect 32137 33405 32171 33439
rect 32171 33405 32180 33439
rect 32128 33396 32180 33405
rect 32404 33439 32456 33448
rect 32404 33405 32413 33439
rect 32413 33405 32447 33439
rect 32447 33405 32456 33439
rect 32404 33396 32456 33405
rect 31024 33328 31076 33380
rect 33416 33328 33468 33380
rect 29184 33260 29236 33312
rect 33140 33260 33192 33312
rect 34060 33260 34112 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 5448 33099 5500 33108
rect 5448 33065 5457 33099
rect 5457 33065 5491 33099
rect 5491 33065 5500 33099
rect 5448 33056 5500 33065
rect 9588 33056 9640 33108
rect 11796 33056 11848 33108
rect 14096 33056 14148 33108
rect 7012 32920 7064 32972
rect 7656 32920 7708 32972
rect 7748 32920 7800 32972
rect 9772 32963 9824 32972
rect 9772 32929 9781 32963
rect 9781 32929 9815 32963
rect 9815 32929 9824 32963
rect 9772 32920 9824 32929
rect 9956 32920 10008 32972
rect 4804 32852 4856 32904
rect 7380 32895 7432 32904
rect 7380 32861 7389 32895
rect 7389 32861 7423 32895
rect 7423 32861 7432 32895
rect 7380 32852 7432 32861
rect 6184 32784 6236 32836
rect 5908 32759 5960 32768
rect 5908 32725 5917 32759
rect 5917 32725 5951 32759
rect 5951 32725 5960 32759
rect 5908 32716 5960 32725
rect 7012 32759 7064 32768
rect 7012 32725 7021 32759
rect 7021 32725 7055 32759
rect 7055 32725 7064 32759
rect 7012 32716 7064 32725
rect 7656 32827 7708 32836
rect 7656 32793 7665 32827
rect 7665 32793 7699 32827
rect 7699 32793 7708 32827
rect 7656 32784 7708 32793
rect 9772 32784 9824 32836
rect 10508 32895 10560 32904
rect 10508 32861 10517 32895
rect 10517 32861 10551 32895
rect 10551 32861 10560 32895
rect 10508 32852 10560 32861
rect 11796 32852 11848 32904
rect 12164 32895 12216 32904
rect 12164 32861 12173 32895
rect 12173 32861 12207 32895
rect 12207 32861 12216 32895
rect 12164 32852 12216 32861
rect 7840 32716 7892 32768
rect 11888 32716 11940 32768
rect 12072 32759 12124 32768
rect 12072 32725 12081 32759
rect 12081 32725 12115 32759
rect 12115 32725 12124 32759
rect 12072 32716 12124 32725
rect 13912 32920 13964 32972
rect 12992 32895 13044 32904
rect 12992 32861 13001 32895
rect 13001 32861 13035 32895
rect 13035 32861 13044 32895
rect 12992 32852 13044 32861
rect 13176 32895 13228 32904
rect 13176 32861 13185 32895
rect 13185 32861 13219 32895
rect 13219 32861 13228 32895
rect 13176 32852 13228 32861
rect 13360 32716 13412 32768
rect 13544 32759 13596 32768
rect 13544 32725 13553 32759
rect 13553 32725 13587 32759
rect 13587 32725 13596 32759
rect 13544 32716 13596 32725
rect 14096 32963 14148 32972
rect 14096 32929 14105 32963
rect 14105 32929 14139 32963
rect 14139 32929 14148 32963
rect 14096 32920 14148 32929
rect 14188 32852 14240 32904
rect 28356 33056 28408 33108
rect 29828 33056 29880 33108
rect 32404 33056 32456 33108
rect 34520 33099 34572 33108
rect 34520 33065 34529 33099
rect 34529 33065 34563 33099
rect 34563 33065 34572 33099
rect 34520 33056 34572 33065
rect 23756 33031 23808 33040
rect 23756 32997 23765 33031
rect 23765 32997 23799 33031
rect 23799 32997 23808 33031
rect 23756 32988 23808 32997
rect 14464 32784 14516 32836
rect 16672 32852 16724 32904
rect 22100 32920 22152 32972
rect 32772 32963 32824 32972
rect 14832 32716 14884 32768
rect 15108 32716 15160 32768
rect 16764 32784 16816 32836
rect 17408 32895 17460 32904
rect 17408 32861 17417 32895
rect 17417 32861 17451 32895
rect 17451 32861 17460 32895
rect 17408 32852 17460 32861
rect 17776 32895 17828 32904
rect 17776 32861 17785 32895
rect 17785 32861 17819 32895
rect 17819 32861 17828 32895
rect 17776 32852 17828 32861
rect 18604 32852 18656 32904
rect 19616 32784 19668 32836
rect 17684 32716 17736 32768
rect 21180 32784 21232 32836
rect 21456 32784 21508 32836
rect 23572 32895 23624 32904
rect 23572 32861 23581 32895
rect 23581 32861 23615 32895
rect 23615 32861 23624 32895
rect 23572 32852 23624 32861
rect 24400 32895 24452 32904
rect 24400 32861 24409 32895
rect 24409 32861 24443 32895
rect 24443 32861 24452 32895
rect 24400 32852 24452 32861
rect 25872 32895 25924 32904
rect 25872 32861 25881 32895
rect 25881 32861 25915 32895
rect 25915 32861 25924 32895
rect 25872 32852 25924 32861
rect 32772 32929 32781 32963
rect 32781 32929 32815 32963
rect 32815 32929 32824 32963
rect 32772 32920 32824 32929
rect 33416 32920 33468 32972
rect 22560 32827 22612 32836
rect 22560 32793 22569 32827
rect 22569 32793 22603 32827
rect 22603 32793 22612 32827
rect 22560 32784 22612 32793
rect 24492 32784 24544 32836
rect 28724 32852 28776 32904
rect 29644 32852 29696 32904
rect 32128 32852 32180 32904
rect 26608 32784 26660 32836
rect 28172 32784 28224 32836
rect 29828 32827 29880 32836
rect 29828 32793 29862 32827
rect 29862 32793 29880 32827
rect 29828 32784 29880 32793
rect 31024 32784 31076 32836
rect 19984 32716 20036 32768
rect 20444 32716 20496 32768
rect 21272 32716 21324 32768
rect 25780 32759 25832 32768
rect 25780 32725 25789 32759
rect 25789 32725 25823 32759
rect 25823 32725 25832 32759
rect 25780 32716 25832 32725
rect 26056 32716 26108 32768
rect 26976 32759 27028 32768
rect 26976 32725 26985 32759
rect 26985 32725 27019 32759
rect 27019 32725 27028 32759
rect 26976 32716 27028 32725
rect 28632 32759 28684 32768
rect 28632 32725 28641 32759
rect 28641 32725 28675 32759
rect 28675 32725 28684 32759
rect 28632 32716 28684 32725
rect 33140 32784 33192 32836
rect 33508 32784 33560 32836
rect 34428 32716 34480 32768
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 4804 32444 4856 32496
rect 3976 32376 4028 32428
rect 5908 32376 5960 32428
rect 7840 32512 7892 32564
rect 9128 32555 9180 32564
rect 9128 32521 9137 32555
rect 9137 32521 9171 32555
rect 9171 32521 9180 32555
rect 9128 32512 9180 32521
rect 9772 32512 9824 32564
rect 10784 32512 10836 32564
rect 12992 32512 13044 32564
rect 13912 32512 13964 32564
rect 14372 32512 14424 32564
rect 14464 32555 14516 32564
rect 14464 32521 14473 32555
rect 14473 32521 14507 32555
rect 14507 32521 14516 32555
rect 14464 32512 14516 32521
rect 14832 32555 14884 32564
rect 14832 32521 14841 32555
rect 14841 32521 14875 32555
rect 14875 32521 14884 32555
rect 14832 32512 14884 32521
rect 8208 32444 8260 32496
rect 9036 32444 9088 32496
rect 12716 32444 12768 32496
rect 12900 32444 12952 32496
rect 14188 32444 14240 32496
rect 16212 32512 16264 32564
rect 16580 32512 16632 32564
rect 19524 32512 19576 32564
rect 19616 32555 19668 32564
rect 19616 32521 19625 32555
rect 19625 32521 19659 32555
rect 19659 32521 19668 32555
rect 19616 32512 19668 32521
rect 19984 32555 20036 32564
rect 19984 32521 19993 32555
rect 19993 32521 20027 32555
rect 20027 32521 20036 32555
rect 19984 32512 20036 32521
rect 20996 32555 21048 32564
rect 20996 32521 21005 32555
rect 21005 32521 21039 32555
rect 21039 32521 21048 32555
rect 20996 32512 21048 32521
rect 21180 32512 21232 32564
rect 3424 32351 3476 32360
rect 3424 32317 3433 32351
rect 3433 32317 3467 32351
rect 3467 32317 3476 32351
rect 3424 32308 3476 32317
rect 9404 32376 9456 32428
rect 9496 32308 9548 32360
rect 10508 32376 10560 32428
rect 12624 32419 12676 32428
rect 12624 32385 12658 32419
rect 12658 32385 12676 32419
rect 12624 32376 12676 32385
rect 15108 32444 15160 32496
rect 18236 32444 18288 32496
rect 19248 32444 19300 32496
rect 25780 32512 25832 32564
rect 28264 32512 28316 32564
rect 28356 32512 28408 32564
rect 34152 32512 34204 32564
rect 11060 32308 11112 32360
rect 11520 32308 11572 32360
rect 13360 32308 13412 32360
rect 17040 32419 17092 32428
rect 17040 32385 17049 32419
rect 17049 32385 17083 32419
rect 17083 32385 17092 32419
rect 17040 32376 17092 32385
rect 4804 32215 4856 32224
rect 4804 32181 4813 32215
rect 4813 32181 4847 32215
rect 4847 32181 4856 32215
rect 4804 32172 4856 32181
rect 6736 32172 6788 32224
rect 7196 32172 7248 32224
rect 13084 32172 13136 32224
rect 13636 32172 13688 32224
rect 15108 32351 15160 32360
rect 15108 32317 15117 32351
rect 15117 32317 15151 32351
rect 15151 32317 15160 32351
rect 15108 32308 15160 32317
rect 14556 32240 14608 32292
rect 14464 32172 14516 32224
rect 16580 32308 16632 32360
rect 17132 32351 17184 32360
rect 17132 32317 17141 32351
rect 17141 32317 17175 32351
rect 17175 32317 17184 32351
rect 17132 32308 17184 32317
rect 17316 32351 17368 32360
rect 17316 32317 17325 32351
rect 17325 32317 17359 32351
rect 17359 32317 17368 32351
rect 17316 32308 17368 32317
rect 21272 32419 21324 32428
rect 21272 32385 21281 32419
rect 21281 32385 21315 32419
rect 21315 32385 21324 32419
rect 21272 32376 21324 32385
rect 21364 32376 21416 32428
rect 16120 32240 16172 32292
rect 21732 32308 21784 32360
rect 15568 32172 15620 32224
rect 17316 32172 17368 32224
rect 20444 32172 20496 32224
rect 22560 32419 22612 32428
rect 22560 32385 22569 32419
rect 22569 32385 22603 32419
rect 22603 32385 22612 32419
rect 22560 32376 22612 32385
rect 22836 32419 22888 32428
rect 22836 32385 22870 32419
rect 22870 32385 22888 32419
rect 22836 32376 22888 32385
rect 23756 32376 23808 32428
rect 26148 32308 26200 32360
rect 23940 32215 23992 32224
rect 23940 32181 23949 32215
rect 23949 32181 23983 32215
rect 23983 32181 23992 32215
rect 23940 32172 23992 32181
rect 24492 32240 24544 32292
rect 27804 32444 27856 32496
rect 28632 32444 28684 32496
rect 29644 32487 29696 32496
rect 29644 32453 29653 32487
rect 29653 32453 29687 32487
rect 29687 32453 29696 32487
rect 29644 32444 29696 32453
rect 27620 32376 27672 32428
rect 28172 32419 28224 32428
rect 28172 32385 28181 32419
rect 28181 32385 28215 32419
rect 28215 32385 28224 32419
rect 28172 32376 28224 32385
rect 28264 32419 28316 32428
rect 28264 32385 28273 32419
rect 28273 32385 28307 32419
rect 28307 32385 28316 32419
rect 28264 32376 28316 32385
rect 28540 32419 28592 32428
rect 28540 32385 28549 32419
rect 28549 32385 28583 32419
rect 28583 32385 28592 32419
rect 28540 32376 28592 32385
rect 28448 32308 28500 32360
rect 29552 32240 29604 32292
rect 30288 32240 30340 32292
rect 26700 32172 26752 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 7104 31968 7156 32020
rect 7380 31968 7432 32020
rect 8852 31968 8904 32020
rect 9312 31968 9364 32020
rect 9588 32011 9640 32020
rect 9588 31977 9597 32011
rect 9597 31977 9631 32011
rect 9631 31977 9640 32011
rect 9588 31968 9640 31977
rect 9864 31968 9916 32020
rect 4712 31832 4764 31884
rect 1400 31807 1452 31816
rect 1400 31773 1409 31807
rect 1409 31773 1443 31807
rect 1443 31773 1452 31807
rect 1400 31764 1452 31773
rect 4620 31807 4672 31816
rect 4620 31773 4629 31807
rect 4629 31773 4663 31807
rect 4663 31773 4672 31807
rect 4620 31764 4672 31773
rect 5264 31807 5316 31816
rect 5264 31773 5273 31807
rect 5273 31773 5307 31807
rect 5307 31773 5316 31807
rect 5264 31764 5316 31773
rect 7288 31875 7340 31884
rect 7288 31841 7297 31875
rect 7297 31841 7331 31875
rect 7331 31841 7340 31875
rect 7288 31832 7340 31841
rect 9496 31900 9548 31952
rect 7196 31807 7248 31816
rect 7196 31773 7205 31807
rect 7205 31773 7239 31807
rect 7239 31773 7248 31807
rect 8208 31832 8260 31884
rect 11060 31968 11112 32020
rect 12624 31968 12676 32020
rect 17132 31968 17184 32020
rect 21456 32011 21508 32020
rect 21456 31977 21465 32011
rect 21465 31977 21499 32011
rect 21499 31977 21508 32011
rect 21456 31968 21508 31977
rect 22100 31968 22152 32020
rect 7196 31764 7248 31773
rect 7472 31764 7524 31816
rect 8116 31807 8168 31816
rect 8116 31773 8125 31807
rect 8125 31773 8159 31807
rect 8159 31773 8168 31807
rect 8116 31764 8168 31773
rect 8760 31764 8812 31816
rect 9128 31807 9180 31816
rect 9128 31773 9135 31807
rect 9135 31773 9180 31807
rect 9128 31764 9180 31773
rect 9312 31807 9364 31816
rect 9312 31773 9321 31807
rect 9321 31773 9355 31807
rect 9355 31773 9364 31807
rect 9312 31764 9364 31773
rect 9404 31807 9456 31816
rect 9404 31773 9418 31807
rect 9418 31773 9452 31807
rect 9452 31773 9456 31807
rect 9404 31764 9456 31773
rect 7104 31739 7156 31748
rect 7104 31705 7113 31739
rect 7113 31705 7147 31739
rect 7147 31705 7156 31739
rect 7104 31696 7156 31705
rect 9864 31764 9916 31816
rect 18236 31900 18288 31952
rect 22836 31968 22888 32020
rect 26056 32011 26108 32020
rect 26056 31977 26065 32011
rect 26065 31977 26099 32011
rect 26099 31977 26108 32011
rect 26056 31968 26108 31977
rect 27988 31968 28040 32020
rect 28540 31968 28592 32020
rect 29828 31968 29880 32020
rect 12716 31832 12768 31884
rect 12072 31764 12124 31816
rect 12992 31764 13044 31816
rect 7564 31628 7616 31680
rect 11888 31696 11940 31748
rect 20904 31832 20956 31884
rect 21180 31832 21232 31884
rect 22100 31875 22152 31884
rect 22100 31841 22109 31875
rect 22109 31841 22143 31875
rect 22143 31841 22152 31875
rect 22100 31832 22152 31841
rect 16672 31764 16724 31816
rect 21272 31764 21324 31816
rect 22928 31900 22980 31952
rect 27896 31900 27948 31952
rect 23756 31764 23808 31816
rect 25872 31807 25924 31816
rect 25872 31773 25881 31807
rect 25881 31773 25915 31807
rect 25915 31773 25924 31807
rect 25872 31764 25924 31773
rect 25964 31807 26016 31816
rect 25964 31773 25973 31807
rect 25973 31773 26007 31807
rect 26007 31773 26016 31807
rect 25964 31764 26016 31773
rect 26792 31764 26844 31816
rect 28540 31807 28592 31816
rect 28540 31773 28549 31807
rect 28549 31773 28583 31807
rect 28583 31773 28592 31807
rect 28540 31764 28592 31773
rect 29920 31832 29972 31884
rect 30104 31832 30156 31884
rect 32772 31875 32824 31884
rect 32772 31841 32781 31875
rect 32781 31841 32815 31875
rect 32815 31841 32824 31875
rect 32772 31832 32824 31841
rect 33784 31832 33836 31884
rect 29460 31764 29512 31816
rect 10692 31628 10744 31680
rect 12072 31671 12124 31680
rect 12072 31637 12081 31671
rect 12081 31637 12115 31671
rect 12115 31637 12124 31671
rect 12072 31628 12124 31637
rect 15568 31739 15620 31748
rect 15568 31705 15602 31739
rect 15602 31705 15620 31739
rect 15568 31696 15620 31705
rect 17776 31696 17828 31748
rect 16120 31628 16172 31680
rect 17408 31628 17460 31680
rect 23020 31696 23072 31748
rect 23112 31696 23164 31748
rect 18144 31628 18196 31680
rect 22744 31628 22796 31680
rect 23296 31628 23348 31680
rect 23480 31671 23532 31680
rect 23480 31637 23489 31671
rect 23489 31637 23523 31671
rect 23523 31637 23532 31671
rect 23480 31628 23532 31637
rect 27068 31696 27120 31748
rect 27436 31696 27488 31748
rect 27528 31696 27580 31748
rect 27804 31628 27856 31680
rect 28172 31696 28224 31748
rect 28908 31696 28960 31748
rect 33508 31696 33560 31748
rect 30380 31671 30432 31680
rect 30380 31637 30389 31671
rect 30389 31637 30423 31671
rect 30423 31637 30432 31671
rect 30380 31628 30432 31637
rect 30840 31671 30892 31680
rect 30840 31637 30849 31671
rect 30849 31637 30883 31671
rect 30883 31637 30892 31671
rect 30840 31628 30892 31637
rect 34520 31671 34572 31680
rect 34520 31637 34529 31671
rect 34529 31637 34563 31671
rect 34563 31637 34572 31671
rect 34520 31628 34572 31637
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 1400 31467 1452 31476
rect 1400 31433 1409 31467
rect 1409 31433 1443 31467
rect 1443 31433 1452 31467
rect 1400 31424 1452 31433
rect 5172 31424 5224 31476
rect 6920 31424 6972 31476
rect 8116 31424 8168 31476
rect 9312 31424 9364 31476
rect 3424 31356 3476 31408
rect 4068 31331 4120 31340
rect 4068 31297 4077 31331
rect 4077 31297 4111 31331
rect 4111 31297 4120 31331
rect 4068 31288 4120 31297
rect 4620 31288 4672 31340
rect 4712 31220 4764 31272
rect 5356 31220 5408 31272
rect 7288 31356 7340 31408
rect 9680 31424 9732 31476
rect 6276 31288 6328 31340
rect 8208 31288 8260 31340
rect 9312 31288 9364 31340
rect 10876 31331 10928 31340
rect 10876 31297 10885 31331
rect 10885 31297 10919 31331
rect 10919 31297 10928 31331
rect 10876 31288 10928 31297
rect 11060 31331 11112 31340
rect 11060 31297 11069 31331
rect 11069 31297 11103 31331
rect 11103 31297 11112 31331
rect 11060 31288 11112 31297
rect 11244 31288 11296 31340
rect 12348 31424 12400 31476
rect 15660 31424 15712 31476
rect 16488 31424 16540 31476
rect 17408 31467 17460 31476
rect 17408 31433 17417 31467
rect 17417 31433 17451 31467
rect 17451 31433 17460 31467
rect 17408 31424 17460 31433
rect 17776 31467 17828 31476
rect 17776 31433 17785 31467
rect 17785 31433 17819 31467
rect 17819 31433 17828 31467
rect 17776 31424 17828 31433
rect 21088 31467 21140 31476
rect 21088 31433 21097 31467
rect 21097 31433 21131 31467
rect 21131 31433 21140 31467
rect 21088 31424 21140 31433
rect 11796 31399 11848 31408
rect 11796 31365 11805 31399
rect 11805 31365 11839 31399
rect 11839 31365 11848 31399
rect 11796 31356 11848 31365
rect 12716 31356 12768 31408
rect 12072 31331 12124 31340
rect 12072 31297 12080 31331
rect 12080 31297 12114 31331
rect 12114 31297 12124 31331
rect 12072 31288 12124 31297
rect 12532 31288 12584 31340
rect 13544 31288 13596 31340
rect 16764 31356 16816 31408
rect 17592 31356 17644 31408
rect 19708 31356 19760 31408
rect 21272 31356 21324 31408
rect 16856 31331 16908 31340
rect 16856 31297 16865 31331
rect 16865 31297 16899 31331
rect 16899 31297 16908 31331
rect 16856 31288 16908 31297
rect 17132 31288 17184 31340
rect 17316 31288 17368 31340
rect 9680 31152 9732 31204
rect 4620 31084 4672 31136
rect 10416 31084 10468 31136
rect 17684 31220 17736 31272
rect 18144 31331 18196 31340
rect 18144 31297 18153 31331
rect 18153 31297 18187 31331
rect 18187 31297 18196 31331
rect 18144 31288 18196 31297
rect 18604 31331 18656 31340
rect 18604 31297 18613 31331
rect 18613 31297 18647 31331
rect 18647 31297 18656 31331
rect 18604 31288 18656 31297
rect 19248 31288 19300 31340
rect 18328 31263 18380 31272
rect 18328 31229 18337 31263
rect 18337 31229 18371 31263
rect 18371 31229 18380 31263
rect 18328 31220 18380 31229
rect 12348 31127 12400 31136
rect 12348 31093 12357 31127
rect 12357 31093 12391 31127
rect 12391 31093 12400 31127
rect 12348 31084 12400 31093
rect 12532 31127 12584 31136
rect 12532 31093 12541 31127
rect 12541 31093 12575 31127
rect 12575 31093 12584 31127
rect 12532 31084 12584 31093
rect 12716 31127 12768 31136
rect 12716 31093 12725 31127
rect 12725 31093 12759 31127
rect 12759 31093 12768 31127
rect 12716 31084 12768 31093
rect 25596 31424 25648 31476
rect 25872 31424 25924 31476
rect 24676 31356 24728 31408
rect 25136 31288 25188 31340
rect 27620 31424 27672 31476
rect 28264 31424 28316 31476
rect 28816 31424 28868 31476
rect 30840 31424 30892 31476
rect 33784 31424 33836 31476
rect 27436 31356 27488 31408
rect 23388 31220 23440 31272
rect 23572 31263 23624 31272
rect 23572 31229 23581 31263
rect 23581 31229 23615 31263
rect 23615 31229 23624 31263
rect 23572 31220 23624 31229
rect 24400 31220 24452 31272
rect 26516 31331 26568 31340
rect 26516 31297 26525 31331
rect 26525 31297 26559 31331
rect 26559 31297 26568 31331
rect 26516 31288 26568 31297
rect 26792 31288 26844 31340
rect 30380 31356 30432 31408
rect 34796 31399 34848 31408
rect 34796 31365 34805 31399
rect 34805 31365 34839 31399
rect 34839 31365 34848 31399
rect 34796 31356 34848 31365
rect 28356 31331 28408 31340
rect 28356 31297 28390 31331
rect 28390 31297 28408 31331
rect 28356 31288 28408 31297
rect 29644 31288 29696 31340
rect 17868 31084 17920 31136
rect 19984 31127 20036 31136
rect 19984 31093 19993 31127
rect 19993 31093 20027 31127
rect 20027 31093 20036 31127
rect 19984 31084 20036 31093
rect 23296 31084 23348 31136
rect 25228 31084 25280 31136
rect 25964 31127 26016 31136
rect 25964 31093 25973 31127
rect 25973 31093 26007 31127
rect 26007 31093 26016 31127
rect 25964 31084 26016 31093
rect 26792 31084 26844 31136
rect 27068 31084 27120 31136
rect 34428 31331 34480 31340
rect 34428 31297 34437 31331
rect 34437 31297 34471 31331
rect 34471 31297 34480 31331
rect 34428 31288 34480 31297
rect 34520 31331 34572 31340
rect 34520 31297 34529 31331
rect 34529 31297 34563 31331
rect 34563 31297 34572 31331
rect 34520 31288 34572 31297
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 3976 30923 4028 30932
rect 3976 30889 3985 30923
rect 3985 30889 4019 30923
rect 4019 30889 4028 30923
rect 3976 30880 4028 30889
rect 6276 30923 6328 30932
rect 6276 30889 6285 30923
rect 6285 30889 6319 30923
rect 6319 30889 6328 30923
rect 6276 30880 6328 30889
rect 7564 30880 7616 30932
rect 23388 30880 23440 30932
rect 23480 30880 23532 30932
rect 23940 30880 23992 30932
rect 10876 30812 10928 30864
rect 15660 30812 15712 30864
rect 16120 30812 16172 30864
rect 18328 30812 18380 30864
rect 4620 30787 4672 30796
rect 4620 30753 4629 30787
rect 4629 30753 4663 30787
rect 4663 30753 4672 30787
rect 4620 30744 4672 30753
rect 6736 30787 6788 30796
rect 6736 30753 6745 30787
rect 6745 30753 6779 30787
rect 6779 30753 6788 30787
rect 6736 30744 6788 30753
rect 19248 30855 19300 30864
rect 19248 30821 19257 30855
rect 19257 30821 19291 30855
rect 19291 30821 19300 30855
rect 19248 30812 19300 30821
rect 4712 30676 4764 30728
rect 4804 30719 4856 30728
rect 4804 30685 4813 30719
rect 4813 30685 4847 30719
rect 4847 30685 4856 30719
rect 4804 30676 4856 30685
rect 4896 30719 4948 30728
rect 4896 30685 4906 30719
rect 4906 30685 4940 30719
rect 4940 30685 4948 30719
rect 4896 30676 4948 30685
rect 5172 30719 5224 30728
rect 5172 30685 5181 30719
rect 5181 30685 5215 30719
rect 5215 30685 5224 30719
rect 5172 30676 5224 30685
rect 5816 30540 5868 30592
rect 6920 30676 6972 30728
rect 7472 30608 7524 30660
rect 19800 30744 19852 30796
rect 11336 30676 11388 30728
rect 12900 30676 12952 30728
rect 13268 30676 13320 30728
rect 15108 30676 15160 30728
rect 15292 30676 15344 30728
rect 15476 30676 15528 30728
rect 12808 30608 12860 30660
rect 10324 30540 10376 30592
rect 10416 30540 10468 30592
rect 13636 30583 13688 30592
rect 13636 30549 13645 30583
rect 13645 30549 13679 30583
rect 13679 30549 13688 30583
rect 13636 30540 13688 30549
rect 14556 30608 14608 30660
rect 19984 30676 20036 30728
rect 15568 30540 15620 30592
rect 15752 30583 15804 30592
rect 15752 30549 15761 30583
rect 15761 30549 15795 30583
rect 15795 30549 15804 30583
rect 15752 30540 15804 30549
rect 17592 30583 17644 30592
rect 17592 30549 17601 30583
rect 17601 30549 17635 30583
rect 17635 30549 17644 30583
rect 17592 30540 17644 30549
rect 19708 30583 19760 30592
rect 19708 30549 19717 30583
rect 19717 30549 19751 30583
rect 19751 30549 19760 30583
rect 19708 30540 19760 30549
rect 21824 30676 21876 30728
rect 23664 30676 23716 30728
rect 25136 30923 25188 30932
rect 25136 30889 25145 30923
rect 25145 30889 25179 30923
rect 25179 30889 25188 30923
rect 25136 30880 25188 30889
rect 25228 30880 25280 30932
rect 27528 30880 27580 30932
rect 28356 30880 28408 30932
rect 25872 30812 25924 30864
rect 25320 30744 25372 30796
rect 28908 30787 28960 30796
rect 28908 30753 28917 30787
rect 28917 30753 28951 30787
rect 28951 30753 28960 30787
rect 28908 30744 28960 30753
rect 30288 30744 30340 30796
rect 20536 30540 20588 30592
rect 22836 30608 22888 30660
rect 20812 30540 20864 30592
rect 21272 30540 21324 30592
rect 23204 30540 23256 30592
rect 24860 30719 24912 30728
rect 24860 30685 24874 30719
rect 24874 30685 24908 30719
rect 24908 30685 24912 30719
rect 24860 30676 24912 30685
rect 25964 30676 26016 30728
rect 28816 30719 28868 30728
rect 28816 30685 28825 30719
rect 28825 30685 28859 30719
rect 28859 30685 28868 30719
rect 28816 30676 28868 30685
rect 29276 30676 29328 30728
rect 24676 30651 24728 30660
rect 24676 30617 24685 30651
rect 24685 30617 24719 30651
rect 24719 30617 24728 30651
rect 24676 30608 24728 30617
rect 25688 30608 25740 30660
rect 25780 30608 25832 30660
rect 27988 30608 28040 30660
rect 24860 30540 24912 30592
rect 25964 30583 26016 30592
rect 25964 30549 25973 30583
rect 25973 30549 26007 30583
rect 26007 30549 26016 30583
rect 25964 30540 26016 30549
rect 27620 30540 27672 30592
rect 27896 30540 27948 30592
rect 29000 30608 29052 30660
rect 30840 30676 30892 30728
rect 31208 30719 31260 30728
rect 31208 30685 31217 30719
rect 31217 30685 31251 30719
rect 31251 30685 31260 30719
rect 31208 30676 31260 30685
rect 34152 30676 34204 30728
rect 33048 30608 33100 30660
rect 34520 30608 34572 30660
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 4620 30336 4672 30388
rect 4804 30379 4856 30388
rect 4804 30345 4813 30379
rect 4813 30345 4847 30379
rect 4847 30345 4856 30379
rect 4804 30336 4856 30345
rect 4896 30268 4948 30320
rect 5356 30268 5408 30320
rect 9220 30268 9272 30320
rect 11060 30311 11112 30320
rect 1308 30200 1360 30252
rect 3608 30200 3660 30252
rect 2872 29996 2924 30048
rect 5448 30200 5500 30252
rect 9772 30200 9824 30252
rect 9312 30132 9364 30184
rect 9588 30175 9640 30184
rect 9588 30141 9597 30175
rect 9597 30141 9631 30175
rect 9631 30141 9640 30175
rect 9588 30132 9640 30141
rect 10232 30132 10284 30184
rect 11060 30277 11069 30311
rect 11069 30277 11103 30311
rect 11103 30277 11112 30311
rect 11060 30268 11112 30277
rect 12808 30379 12860 30388
rect 12808 30345 12817 30379
rect 12817 30345 12851 30379
rect 12851 30345 12860 30379
rect 12808 30336 12860 30345
rect 14464 30336 14516 30388
rect 14556 30379 14608 30388
rect 14556 30345 14565 30379
rect 14565 30345 14599 30379
rect 14599 30345 14608 30379
rect 14556 30336 14608 30345
rect 15292 30336 15344 30388
rect 15752 30336 15804 30388
rect 16304 30336 16356 30388
rect 13084 30268 13136 30320
rect 13636 30268 13688 30320
rect 14280 30268 14332 30320
rect 18144 30268 18196 30320
rect 19708 30336 19760 30388
rect 20812 30379 20864 30388
rect 20812 30345 20821 30379
rect 20821 30345 20855 30379
rect 20855 30345 20864 30379
rect 20812 30336 20864 30345
rect 21272 30379 21324 30388
rect 21272 30345 21281 30379
rect 21281 30345 21315 30379
rect 21315 30345 21324 30379
rect 21272 30336 21324 30345
rect 22836 30379 22888 30388
rect 22836 30345 22845 30379
rect 22845 30345 22879 30379
rect 22879 30345 22888 30379
rect 22836 30336 22888 30345
rect 23204 30379 23256 30388
rect 23204 30345 23213 30379
rect 23213 30345 23247 30379
rect 23247 30345 23256 30379
rect 23204 30336 23256 30345
rect 24676 30336 24728 30388
rect 25780 30336 25832 30388
rect 18512 30268 18564 30320
rect 20904 30268 20956 30320
rect 21180 30311 21232 30320
rect 21180 30277 21189 30311
rect 21189 30277 21223 30311
rect 21223 30277 21232 30311
rect 21180 30268 21232 30277
rect 10600 30243 10652 30252
rect 10600 30209 10609 30243
rect 10609 30209 10643 30243
rect 10643 30209 10652 30243
rect 10600 30200 10652 30209
rect 10692 30243 10744 30252
rect 10692 30209 10701 30243
rect 10701 30209 10735 30243
rect 10735 30209 10744 30243
rect 10692 30200 10744 30209
rect 11888 30200 11940 30252
rect 12716 30200 12768 30252
rect 4620 30064 4672 30116
rect 9036 30064 9088 30116
rect 11244 30064 11296 30116
rect 4804 29996 4856 30048
rect 8944 30039 8996 30048
rect 8944 30005 8953 30039
rect 8953 30005 8987 30039
rect 8987 30005 8996 30039
rect 8944 29996 8996 30005
rect 9588 29996 9640 30048
rect 11060 29996 11112 30048
rect 13268 30132 13320 30184
rect 14096 30200 14148 30252
rect 15200 30200 15252 30252
rect 15568 30243 15620 30252
rect 15568 30209 15578 30243
rect 15578 30209 15612 30243
rect 15612 30209 15620 30243
rect 15568 30200 15620 30209
rect 13176 30064 13228 30116
rect 14280 29996 14332 30048
rect 15660 30132 15712 30184
rect 15844 30243 15896 30252
rect 15844 30209 15853 30243
rect 15853 30209 15887 30243
rect 15887 30209 15896 30243
rect 15844 30200 15896 30209
rect 16212 30200 16264 30252
rect 16580 30132 16632 30184
rect 17040 30132 17092 30184
rect 16856 30064 16908 30116
rect 18420 30243 18472 30252
rect 18420 30209 18429 30243
rect 18429 30209 18463 30243
rect 18463 30209 18472 30243
rect 18420 30200 18472 30209
rect 24492 30268 24544 30320
rect 18328 30064 18380 30116
rect 18696 30064 18748 30116
rect 20628 30132 20680 30184
rect 23020 30200 23072 30252
rect 21640 30132 21692 30184
rect 21916 30064 21968 30116
rect 23296 30175 23348 30184
rect 23296 30141 23305 30175
rect 23305 30141 23339 30175
rect 23339 30141 23348 30175
rect 23296 30132 23348 30141
rect 27068 30243 27120 30252
rect 27068 30209 27078 30243
rect 27078 30209 27112 30243
rect 27112 30209 27120 30243
rect 27068 30200 27120 30209
rect 14556 29996 14608 30048
rect 16304 29996 16356 30048
rect 19340 29996 19392 30048
rect 20720 29996 20772 30048
rect 27160 30132 27212 30184
rect 24492 30064 24544 30116
rect 27344 30243 27396 30252
rect 27344 30209 27353 30243
rect 27353 30209 27387 30243
rect 27387 30209 27396 30243
rect 27344 30200 27396 30209
rect 34152 30268 34204 30320
rect 24032 29996 24084 30048
rect 25320 29996 25372 30048
rect 25596 29996 25648 30048
rect 26056 29996 26108 30048
rect 29000 30064 29052 30116
rect 27528 29996 27580 30048
rect 29092 30039 29144 30048
rect 29092 30005 29101 30039
rect 29101 30005 29135 30039
rect 29135 30005 29144 30039
rect 33048 30200 33100 30252
rect 34244 30200 34296 30252
rect 33508 30064 33560 30116
rect 29092 29996 29144 30005
rect 30196 29996 30248 30048
rect 33416 30039 33468 30048
rect 33416 30005 33425 30039
rect 33425 30005 33459 30039
rect 33459 30005 33468 30039
rect 33416 29996 33468 30005
rect 33600 30039 33652 30048
rect 33600 30005 33609 30039
rect 33609 30005 33643 30039
rect 33643 30005 33652 30039
rect 33600 29996 33652 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 3608 29835 3660 29844
rect 3608 29801 3617 29835
rect 3617 29801 3651 29835
rect 3651 29801 3660 29835
rect 3608 29792 3660 29801
rect 8760 29835 8812 29844
rect 8760 29801 8769 29835
rect 8769 29801 8803 29835
rect 8803 29801 8812 29835
rect 8760 29792 8812 29801
rect 10600 29792 10652 29844
rect 11060 29792 11112 29844
rect 5264 29699 5316 29708
rect 5264 29665 5273 29699
rect 5273 29665 5307 29699
rect 5307 29665 5316 29699
rect 5264 29656 5316 29665
rect 2228 29631 2280 29640
rect 2228 29597 2237 29631
rect 2237 29597 2271 29631
rect 2271 29597 2280 29631
rect 2228 29588 2280 29597
rect 3056 29520 3108 29572
rect 4252 29520 4304 29572
rect 4528 29520 4580 29572
rect 4896 29520 4948 29572
rect 6276 29520 6328 29572
rect 4620 29452 4672 29504
rect 6736 29452 6788 29504
rect 8576 29631 8628 29640
rect 8576 29597 8585 29631
rect 8585 29597 8619 29631
rect 8619 29597 8628 29631
rect 9036 29631 9088 29640
rect 8576 29588 8628 29597
rect 9036 29597 9045 29631
rect 9045 29597 9079 29631
rect 9079 29597 9088 29631
rect 9036 29588 9088 29597
rect 7380 29520 7432 29572
rect 7748 29452 7800 29504
rect 11336 29699 11388 29708
rect 11336 29665 11345 29699
rect 11345 29665 11379 29699
rect 11379 29665 11388 29699
rect 11336 29656 11388 29665
rect 14372 29835 14424 29844
rect 14372 29801 14381 29835
rect 14381 29801 14415 29835
rect 14415 29801 14424 29835
rect 14372 29792 14424 29801
rect 15200 29792 15252 29844
rect 18420 29792 18472 29844
rect 20536 29792 20588 29844
rect 20628 29835 20680 29844
rect 20628 29801 20637 29835
rect 20637 29801 20671 29835
rect 20671 29801 20680 29835
rect 20628 29792 20680 29801
rect 9588 29631 9640 29640
rect 9588 29597 9597 29631
rect 9597 29597 9631 29631
rect 9631 29597 9640 29631
rect 9588 29588 9640 29597
rect 13084 29588 13136 29640
rect 14280 29656 14332 29708
rect 14096 29588 14148 29640
rect 14648 29631 14700 29640
rect 14648 29597 14657 29631
rect 14657 29597 14691 29631
rect 14691 29597 14700 29631
rect 14648 29588 14700 29597
rect 15108 29588 15160 29640
rect 16672 29656 16724 29708
rect 10140 29520 10192 29572
rect 10508 29452 10560 29504
rect 15752 29520 15804 29572
rect 17408 29520 17460 29572
rect 19248 29631 19300 29640
rect 19248 29597 19257 29631
rect 19257 29597 19291 29631
rect 19291 29597 19300 29631
rect 19248 29588 19300 29597
rect 19340 29588 19392 29640
rect 21088 29724 21140 29776
rect 21364 29792 21416 29844
rect 23664 29835 23716 29844
rect 23664 29801 23673 29835
rect 23673 29801 23707 29835
rect 23707 29801 23716 29835
rect 23664 29792 23716 29801
rect 25044 29792 25096 29844
rect 27068 29792 27120 29844
rect 27160 29792 27212 29844
rect 27344 29792 27396 29844
rect 29920 29792 29972 29844
rect 34152 29792 34204 29844
rect 22008 29656 22060 29708
rect 23204 29588 23256 29640
rect 23572 29588 23624 29640
rect 29368 29767 29420 29776
rect 29368 29733 29377 29767
rect 29377 29733 29411 29767
rect 29411 29733 29420 29767
rect 29368 29724 29420 29733
rect 24400 29699 24452 29708
rect 24400 29665 24409 29699
rect 24409 29665 24443 29699
rect 24443 29665 24452 29699
rect 24400 29656 24452 29665
rect 27252 29656 27304 29708
rect 25504 29588 25556 29640
rect 29552 29588 29604 29640
rect 33600 29656 33652 29708
rect 15844 29452 15896 29504
rect 18328 29495 18380 29504
rect 18328 29461 18337 29495
rect 18337 29461 18371 29495
rect 18371 29461 18380 29495
rect 18328 29452 18380 29461
rect 19892 29452 19944 29504
rect 23664 29520 23716 29572
rect 24676 29563 24728 29572
rect 24676 29529 24710 29563
rect 24710 29529 24728 29563
rect 24676 29520 24728 29529
rect 26976 29520 27028 29572
rect 28540 29520 28592 29572
rect 29828 29563 29880 29572
rect 29828 29529 29837 29563
rect 29837 29529 29871 29563
rect 29871 29529 29880 29563
rect 29828 29520 29880 29529
rect 29920 29563 29972 29572
rect 29920 29529 29929 29563
rect 29929 29529 29963 29563
rect 29963 29529 29972 29563
rect 29920 29520 29972 29529
rect 32772 29631 32824 29640
rect 32772 29597 32781 29631
rect 32781 29597 32815 29631
rect 32815 29597 32824 29631
rect 32772 29588 32824 29597
rect 33508 29520 33560 29572
rect 22100 29452 22152 29504
rect 22376 29495 22428 29504
rect 22376 29461 22385 29495
rect 22385 29461 22419 29495
rect 22419 29461 22428 29495
rect 22376 29452 22428 29461
rect 23020 29452 23072 29504
rect 26424 29452 26476 29504
rect 27528 29452 27580 29504
rect 29092 29452 29144 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 3056 29291 3108 29300
rect 3056 29257 3065 29291
rect 3065 29257 3099 29291
rect 3099 29257 3108 29291
rect 3056 29248 3108 29257
rect 3608 29248 3660 29300
rect 4252 29291 4304 29300
rect 4252 29257 4261 29291
rect 4261 29257 4295 29291
rect 4295 29257 4304 29291
rect 4252 29248 4304 29257
rect 4620 29291 4672 29300
rect 4620 29257 4629 29291
rect 4629 29257 4663 29291
rect 4663 29257 4672 29291
rect 4620 29248 4672 29257
rect 4712 29291 4764 29300
rect 4712 29257 4721 29291
rect 4721 29257 4755 29291
rect 4755 29257 4764 29291
rect 4712 29248 4764 29257
rect 6736 29291 6788 29300
rect 6736 29257 6745 29291
rect 6745 29257 6779 29291
rect 6779 29257 6788 29291
rect 6736 29248 6788 29257
rect 6828 29291 6880 29300
rect 6828 29257 6837 29291
rect 6837 29257 6871 29291
rect 6871 29257 6880 29291
rect 6828 29248 6880 29257
rect 7380 29291 7432 29300
rect 7380 29257 7389 29291
rect 7389 29257 7423 29291
rect 7423 29257 7432 29291
rect 7380 29248 7432 29257
rect 7748 29291 7800 29300
rect 7748 29257 7757 29291
rect 7757 29257 7791 29291
rect 7791 29257 7800 29291
rect 7748 29248 7800 29257
rect 6368 29180 6420 29232
rect 3700 29087 3752 29096
rect 3700 29053 3709 29087
rect 3709 29053 3743 29087
rect 3743 29053 3752 29087
rect 3700 29044 3752 29053
rect 5632 29112 5684 29164
rect 9680 29248 9732 29300
rect 9772 29291 9824 29300
rect 9772 29257 9781 29291
rect 9781 29257 9815 29291
rect 9815 29257 9824 29291
rect 9772 29248 9824 29257
rect 10140 29291 10192 29300
rect 10140 29257 10149 29291
rect 10149 29257 10183 29291
rect 10183 29257 10192 29291
rect 10140 29248 10192 29257
rect 10600 29248 10652 29300
rect 8208 29180 8260 29232
rect 9588 29180 9640 29232
rect 15292 29248 15344 29300
rect 15752 29291 15804 29300
rect 15752 29257 15761 29291
rect 15761 29257 15795 29291
rect 15795 29257 15804 29291
rect 15752 29248 15804 29257
rect 15844 29248 15896 29300
rect 17408 29291 17460 29300
rect 17408 29257 17417 29291
rect 17417 29257 17451 29291
rect 17451 29257 17460 29291
rect 17408 29248 17460 29257
rect 18328 29248 18380 29300
rect 8944 29112 8996 29164
rect 11980 29112 12032 29164
rect 5264 29044 5316 29096
rect 5540 29044 5592 29096
rect 6184 29044 6236 29096
rect 3792 28976 3844 29028
rect 6276 28976 6328 29028
rect 10416 29044 10468 29096
rect 12992 29087 13044 29096
rect 12992 29053 13001 29087
rect 13001 29053 13035 29087
rect 13035 29053 13044 29087
rect 12992 29044 13044 29053
rect 8668 28908 8720 28960
rect 14648 29112 14700 29164
rect 16028 29044 16080 29096
rect 19248 29180 19300 29232
rect 22100 29223 22152 29232
rect 22100 29189 22134 29223
rect 22134 29189 22152 29223
rect 22100 29180 22152 29189
rect 20260 29112 20312 29164
rect 21824 29155 21876 29164
rect 21824 29121 21833 29155
rect 21833 29121 21867 29155
rect 21867 29121 21876 29155
rect 21824 29112 21876 29121
rect 23204 29291 23256 29300
rect 23204 29257 23213 29291
rect 23213 29257 23247 29291
rect 23247 29257 23256 29291
rect 23204 29248 23256 29257
rect 24676 29291 24728 29300
rect 24676 29257 24685 29291
rect 24685 29257 24719 29291
rect 24719 29257 24728 29291
rect 24676 29248 24728 29257
rect 25044 29291 25096 29300
rect 25044 29257 25053 29291
rect 25053 29257 25087 29291
rect 25087 29257 25096 29291
rect 25044 29248 25096 29257
rect 22376 29180 22428 29232
rect 23296 29180 23348 29232
rect 25688 29248 25740 29300
rect 26976 29291 27028 29300
rect 26976 29257 26985 29291
rect 26985 29257 27019 29291
rect 27019 29257 27028 29291
rect 26976 29248 27028 29257
rect 27344 29248 27396 29300
rect 28540 29291 28592 29300
rect 28540 29257 28549 29291
rect 28549 29257 28583 29291
rect 28583 29257 28592 29291
rect 28540 29248 28592 29257
rect 29368 29248 29420 29300
rect 29828 29248 29880 29300
rect 19708 28976 19760 29028
rect 21640 29044 21692 29096
rect 19156 28908 19208 28960
rect 21088 29019 21140 29028
rect 21088 28985 21097 29019
rect 21097 28985 21131 29019
rect 21131 28985 21140 29019
rect 21088 28976 21140 28985
rect 23664 29155 23716 29164
rect 23664 29121 23673 29155
rect 23673 29121 23707 29155
rect 23707 29121 23716 29155
rect 23664 29112 23716 29121
rect 27436 29112 27488 29164
rect 32772 29180 32824 29232
rect 29736 29155 29788 29164
rect 29736 29121 29770 29155
rect 29770 29121 29788 29155
rect 29736 29112 29788 29121
rect 23480 29044 23532 29096
rect 25872 29044 25924 29096
rect 27528 29087 27580 29096
rect 27528 29053 27537 29087
rect 27537 29053 27571 29087
rect 27571 29053 27580 29087
rect 27528 29044 27580 29053
rect 29092 29087 29144 29096
rect 29092 29053 29101 29087
rect 29101 29053 29135 29087
rect 29135 29053 29144 29087
rect 29092 29044 29144 29053
rect 20720 28908 20772 28960
rect 23020 28908 23072 28960
rect 23296 28951 23348 28960
rect 23296 28917 23305 28951
rect 23305 28917 23339 28951
rect 23339 28917 23348 28951
rect 23296 28908 23348 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 6368 28747 6420 28756
rect 6368 28713 6377 28747
rect 6377 28713 6411 28747
rect 6411 28713 6420 28747
rect 6368 28704 6420 28713
rect 20260 28747 20312 28756
rect 20260 28713 20269 28747
rect 20269 28713 20303 28747
rect 20303 28713 20312 28747
rect 20260 28704 20312 28713
rect 6184 28636 6236 28688
rect 20352 28636 20404 28688
rect 19708 28568 19760 28620
rect 23480 28704 23532 28756
rect 23664 28704 23716 28756
rect 29736 28747 29788 28756
rect 29736 28713 29745 28747
rect 29745 28713 29779 28747
rect 29779 28713 29788 28747
rect 29736 28704 29788 28713
rect 27160 28611 27212 28620
rect 27160 28577 27169 28611
rect 27169 28577 27203 28611
rect 27203 28577 27212 28611
rect 27160 28568 27212 28577
rect 29368 28568 29420 28620
rect 5540 28543 5592 28552
rect 5540 28509 5549 28543
rect 5549 28509 5583 28543
rect 5583 28509 5592 28543
rect 5540 28500 5592 28509
rect 8208 28500 8260 28552
rect 15016 28500 15068 28552
rect 21088 28500 21140 28552
rect 21824 28500 21876 28552
rect 22284 28500 22336 28552
rect 23296 28500 23348 28552
rect 23388 28500 23440 28552
rect 27620 28432 27672 28484
rect 3424 28407 3476 28416
rect 3424 28373 3433 28407
rect 3433 28373 3467 28407
rect 3467 28373 3476 28407
rect 3424 28364 3476 28373
rect 5264 28364 5316 28416
rect 10232 28364 10284 28416
rect 17224 28407 17276 28416
rect 17224 28373 17233 28407
rect 17233 28373 17267 28407
rect 17267 28373 17276 28407
rect 17224 28364 17276 28373
rect 22744 28364 22796 28416
rect 28172 28432 28224 28484
rect 29828 28500 29880 28552
rect 27988 28364 28040 28416
rect 29368 28407 29420 28416
rect 29368 28373 29377 28407
rect 29377 28373 29411 28407
rect 29411 28373 29420 28407
rect 29368 28364 29420 28373
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 2872 28092 2924 28144
rect 4712 28092 4764 28144
rect 1308 28024 1360 28076
rect 3424 28024 3476 28076
rect 4160 28067 4212 28076
rect 4160 28033 4169 28067
rect 4169 28033 4203 28067
rect 4203 28033 4212 28067
rect 4160 28024 4212 28033
rect 4252 28067 4304 28076
rect 4252 28033 4261 28067
rect 4261 28033 4295 28067
rect 4295 28033 4304 28067
rect 4252 28024 4304 28033
rect 3792 27956 3844 28008
rect 4896 28024 4948 28076
rect 5264 28092 5316 28144
rect 10048 28160 10100 28212
rect 14188 28203 14240 28212
rect 14188 28169 14197 28203
rect 14197 28169 14231 28203
rect 14231 28169 14240 28203
rect 14188 28160 14240 28169
rect 15476 28092 15528 28144
rect 16212 28160 16264 28212
rect 23112 28203 23164 28212
rect 23112 28169 23121 28203
rect 23121 28169 23155 28203
rect 23155 28169 23164 28203
rect 23112 28160 23164 28169
rect 24768 28160 24820 28212
rect 26884 28160 26936 28212
rect 27068 28160 27120 28212
rect 27620 28203 27672 28212
rect 27620 28169 27629 28203
rect 27629 28169 27663 28203
rect 27663 28169 27672 28203
rect 27620 28160 27672 28169
rect 27988 28203 28040 28212
rect 27988 28169 27997 28203
rect 27997 28169 28031 28203
rect 28031 28169 28040 28203
rect 27988 28160 28040 28169
rect 6092 28024 6144 28076
rect 7472 28067 7524 28076
rect 7472 28033 7481 28067
rect 7481 28033 7515 28067
rect 7515 28033 7524 28067
rect 7472 28024 7524 28033
rect 7564 28067 7616 28076
rect 7564 28033 7573 28067
rect 7573 28033 7607 28067
rect 7607 28033 7616 28067
rect 7564 28024 7616 28033
rect 12164 28024 12216 28076
rect 16672 28067 16724 28076
rect 16672 28033 16681 28067
rect 16681 28033 16715 28067
rect 16715 28033 16724 28067
rect 16672 28024 16724 28033
rect 16764 28024 16816 28076
rect 20076 28067 20128 28076
rect 20076 28033 20085 28067
rect 20085 28033 20119 28067
rect 20119 28033 20128 28067
rect 20076 28024 20128 28033
rect 4804 27956 4856 28008
rect 4804 27863 4856 27872
rect 4804 27829 4813 27863
rect 4813 27829 4847 27863
rect 4847 27829 4856 27863
rect 4804 27820 4856 27829
rect 9956 27956 10008 28008
rect 12992 27956 13044 28008
rect 14556 27956 14608 28008
rect 15108 27999 15160 28008
rect 15108 27965 15117 27999
rect 15117 27965 15151 27999
rect 15151 27965 15160 27999
rect 15108 27956 15160 27965
rect 20168 27999 20220 28008
rect 20168 27965 20177 27999
rect 20177 27965 20211 27999
rect 20211 27965 20220 27999
rect 20168 27956 20220 27965
rect 20444 27956 20496 28008
rect 7196 27888 7248 27940
rect 9036 27888 9088 27940
rect 22652 28024 22704 28076
rect 25596 28024 25648 28076
rect 26424 28024 26476 28076
rect 29000 28024 29052 28076
rect 34520 28067 34572 28076
rect 34520 28033 34529 28067
rect 34529 28033 34563 28067
rect 34563 28033 34572 28067
rect 34520 28024 34572 28033
rect 22284 27956 22336 28008
rect 24124 27956 24176 28008
rect 23296 27888 23348 27940
rect 23848 27888 23900 27940
rect 28172 27999 28224 28008
rect 28172 27965 28181 27999
rect 28181 27965 28215 27999
rect 28215 27965 28224 27999
rect 28172 27956 28224 27965
rect 35348 27956 35400 28008
rect 29920 27888 29972 27940
rect 5356 27820 5408 27872
rect 6276 27820 6328 27872
rect 8300 27820 8352 27872
rect 8852 27863 8904 27872
rect 8852 27829 8861 27863
rect 8861 27829 8895 27863
rect 8895 27829 8904 27863
rect 8852 27820 8904 27829
rect 11796 27820 11848 27872
rect 12532 27820 12584 27872
rect 13084 27820 13136 27872
rect 18052 27863 18104 27872
rect 18052 27829 18061 27863
rect 18061 27829 18095 27863
rect 18095 27829 18104 27863
rect 18052 27820 18104 27829
rect 18144 27863 18196 27872
rect 18144 27829 18153 27863
rect 18153 27829 18187 27863
rect 18187 27829 18196 27863
rect 18144 27820 18196 27829
rect 19708 27863 19760 27872
rect 19708 27829 19717 27863
rect 19717 27829 19751 27863
rect 19751 27829 19760 27863
rect 19708 27820 19760 27829
rect 20628 27863 20680 27872
rect 20628 27829 20637 27863
rect 20637 27829 20671 27863
rect 20671 27829 20680 27863
rect 20628 27820 20680 27829
rect 21640 27820 21692 27872
rect 22100 27820 22152 27872
rect 26424 27863 26476 27872
rect 26424 27829 26433 27863
rect 26433 27829 26467 27863
rect 26467 27829 26476 27863
rect 26424 27820 26476 27829
rect 26516 27863 26568 27872
rect 26516 27829 26525 27863
rect 26525 27829 26559 27863
rect 26559 27829 26568 27863
rect 26516 27820 26568 27829
rect 27436 27820 27488 27872
rect 29000 27820 29052 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 6092 27659 6144 27668
rect 6092 27625 6101 27659
rect 6101 27625 6135 27659
rect 6135 27625 6144 27659
rect 6092 27616 6144 27625
rect 7472 27616 7524 27668
rect 15844 27616 15896 27668
rect 16764 27659 16816 27668
rect 16764 27625 16773 27659
rect 16773 27625 16807 27659
rect 16807 27625 16816 27659
rect 16764 27616 16816 27625
rect 4068 27548 4120 27600
rect 12164 27591 12216 27600
rect 12164 27557 12173 27591
rect 12173 27557 12207 27591
rect 12207 27557 12216 27591
rect 12164 27548 12216 27557
rect 2228 27523 2280 27532
rect 2228 27489 2237 27523
rect 2237 27489 2271 27523
rect 2271 27489 2280 27523
rect 2228 27480 2280 27489
rect 4252 27480 4304 27532
rect 7196 27480 7248 27532
rect 8208 27480 8260 27532
rect 6184 27455 6236 27464
rect 6184 27421 6193 27455
rect 6193 27421 6227 27455
rect 6227 27421 6236 27455
rect 6184 27412 6236 27421
rect 8300 27412 8352 27464
rect 9128 27480 9180 27532
rect 10692 27480 10744 27532
rect 9036 27455 9088 27464
rect 9036 27421 9045 27455
rect 9045 27421 9079 27455
rect 9079 27421 9088 27455
rect 9036 27412 9088 27421
rect 9220 27455 9272 27464
rect 2596 27344 2648 27396
rect 3056 27344 3108 27396
rect 6276 27344 6328 27396
rect 6828 27344 6880 27396
rect 9220 27421 9229 27455
rect 9229 27421 9263 27455
rect 9263 27421 9272 27455
rect 9220 27412 9272 27421
rect 9588 27455 9640 27464
rect 9588 27421 9597 27455
rect 9597 27421 9631 27455
rect 9631 27421 9640 27455
rect 9588 27412 9640 27421
rect 11796 27455 11848 27464
rect 11796 27421 11805 27455
rect 11805 27421 11839 27455
rect 11839 27421 11848 27455
rect 11796 27412 11848 27421
rect 11980 27480 12032 27532
rect 13544 27548 13596 27600
rect 15660 27548 15712 27600
rect 17960 27548 18012 27600
rect 14096 27480 14148 27532
rect 16948 27480 17000 27532
rect 18144 27616 18196 27668
rect 20168 27616 20220 27668
rect 20536 27616 20588 27668
rect 20904 27616 20956 27668
rect 22376 27616 22428 27668
rect 25596 27659 25648 27668
rect 25596 27625 25605 27659
rect 25605 27625 25639 27659
rect 25639 27625 25648 27659
rect 25596 27616 25648 27625
rect 34520 27659 34572 27668
rect 34520 27625 34529 27659
rect 34529 27625 34563 27659
rect 34563 27625 34572 27659
rect 34520 27616 34572 27625
rect 22468 27480 22520 27532
rect 24216 27548 24268 27600
rect 31852 27548 31904 27600
rect 14280 27412 14332 27464
rect 14556 27455 14608 27464
rect 14556 27421 14565 27455
rect 14565 27421 14599 27455
rect 14599 27421 14608 27455
rect 14556 27412 14608 27421
rect 16028 27455 16080 27464
rect 10140 27344 10192 27396
rect 12900 27344 12952 27396
rect 16028 27421 16037 27455
rect 16037 27421 16071 27455
rect 16071 27421 16080 27455
rect 16028 27412 16080 27421
rect 16212 27455 16264 27464
rect 16212 27421 16221 27455
rect 16221 27421 16255 27455
rect 16255 27421 16264 27455
rect 16212 27412 16264 27421
rect 16396 27455 16448 27464
rect 16396 27421 16405 27455
rect 16405 27421 16439 27455
rect 16439 27421 16448 27455
rect 16396 27412 16448 27421
rect 18052 27412 18104 27464
rect 15108 27344 15160 27396
rect 3884 27319 3936 27328
rect 3884 27285 3893 27319
rect 3893 27285 3927 27319
rect 3927 27285 3936 27319
rect 3884 27276 3936 27285
rect 4344 27319 4396 27328
rect 4344 27285 4353 27319
rect 4353 27285 4387 27319
rect 4387 27285 4396 27319
rect 4344 27276 4396 27285
rect 4620 27276 4672 27328
rect 4896 27276 4948 27328
rect 8024 27319 8076 27328
rect 8024 27285 8033 27319
rect 8033 27285 8067 27319
rect 8067 27285 8076 27319
rect 8024 27276 8076 27285
rect 9772 27276 9824 27328
rect 10968 27319 11020 27328
rect 10968 27285 10977 27319
rect 10977 27285 11011 27319
rect 11011 27285 11020 27319
rect 10968 27276 11020 27285
rect 11612 27276 11664 27328
rect 12624 27276 12676 27328
rect 13912 27319 13964 27328
rect 13912 27285 13921 27319
rect 13921 27285 13955 27319
rect 13955 27285 13964 27319
rect 13912 27276 13964 27285
rect 14096 27319 14148 27328
rect 14096 27285 14105 27319
rect 14105 27285 14139 27319
rect 14139 27285 14148 27319
rect 14096 27276 14148 27285
rect 14280 27276 14332 27328
rect 15016 27276 15068 27328
rect 15936 27319 15988 27328
rect 15936 27285 15945 27319
rect 15945 27285 15979 27319
rect 15979 27285 15988 27319
rect 17316 27344 17368 27396
rect 18972 27344 19024 27396
rect 19708 27344 19760 27396
rect 21456 27344 21508 27396
rect 22100 27412 22152 27464
rect 22652 27455 22704 27464
rect 22652 27421 22661 27455
rect 22661 27421 22695 27455
rect 22695 27421 22704 27455
rect 22652 27412 22704 27421
rect 23204 27412 23256 27464
rect 23756 27480 23808 27532
rect 26148 27523 26200 27532
rect 26148 27489 26157 27523
rect 26157 27489 26191 27523
rect 26191 27489 26200 27523
rect 26148 27480 26200 27489
rect 27528 27480 27580 27532
rect 28724 27480 28776 27532
rect 29276 27480 29328 27532
rect 30104 27523 30156 27532
rect 30104 27489 30113 27523
rect 30113 27489 30147 27523
rect 30147 27489 30156 27523
rect 30104 27480 30156 27489
rect 23664 27455 23716 27464
rect 23664 27421 23673 27455
rect 23673 27421 23707 27455
rect 23707 27421 23716 27455
rect 23664 27412 23716 27421
rect 26424 27412 26476 27464
rect 27160 27455 27212 27464
rect 27160 27421 27169 27455
rect 27169 27421 27203 27455
rect 27203 27421 27212 27455
rect 27160 27412 27212 27421
rect 27436 27455 27488 27464
rect 27436 27421 27445 27455
rect 27445 27421 27479 27455
rect 27479 27421 27488 27455
rect 27436 27412 27488 27421
rect 22284 27344 22336 27396
rect 15936 27276 15988 27285
rect 16580 27319 16632 27328
rect 16580 27285 16589 27319
rect 16589 27285 16623 27319
rect 16623 27285 16632 27319
rect 16580 27276 16632 27285
rect 16764 27276 16816 27328
rect 17224 27319 17276 27328
rect 17224 27285 17233 27319
rect 17233 27285 17267 27319
rect 17267 27285 17276 27319
rect 17224 27276 17276 27285
rect 17500 27276 17552 27328
rect 17776 27276 17828 27328
rect 26516 27344 26568 27396
rect 23848 27319 23900 27328
rect 23848 27285 23857 27319
rect 23857 27285 23891 27319
rect 23891 27285 23900 27319
rect 23848 27276 23900 27285
rect 26976 27276 27028 27328
rect 27620 27319 27672 27328
rect 27620 27285 27629 27319
rect 27629 27285 27663 27319
rect 27663 27285 27672 27319
rect 27620 27276 27672 27285
rect 29092 27412 29144 27464
rect 31484 27412 31536 27464
rect 31760 27480 31812 27532
rect 32772 27523 32824 27532
rect 32772 27489 32781 27523
rect 32781 27489 32815 27523
rect 32815 27489 32824 27523
rect 32772 27480 32824 27489
rect 27988 27319 28040 27328
rect 27988 27285 27997 27319
rect 27997 27285 28031 27319
rect 28031 27285 28040 27319
rect 27988 27276 28040 27285
rect 28724 27319 28776 27328
rect 28724 27285 28733 27319
rect 28733 27285 28767 27319
rect 28767 27285 28776 27319
rect 28724 27276 28776 27285
rect 30104 27344 30156 27396
rect 33324 27344 33376 27396
rect 34060 27344 34112 27396
rect 29644 27276 29696 27328
rect 29920 27319 29972 27328
rect 29920 27285 29929 27319
rect 29929 27285 29963 27319
rect 29963 27285 29972 27319
rect 29920 27276 29972 27285
rect 30012 27319 30064 27328
rect 30012 27285 30021 27319
rect 30021 27285 30055 27319
rect 30055 27285 30064 27319
rect 30012 27276 30064 27285
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 2596 27115 2648 27124
rect 2596 27081 2605 27115
rect 2605 27081 2639 27115
rect 2639 27081 2648 27115
rect 2596 27072 2648 27081
rect 4160 27072 4212 27124
rect 4344 27072 4396 27124
rect 4712 27072 4764 27124
rect 6828 27115 6880 27124
rect 6828 27081 6837 27115
rect 6837 27081 6871 27115
rect 6871 27081 6880 27115
rect 6828 27072 6880 27081
rect 7472 27072 7524 27124
rect 9220 27072 9272 27124
rect 10140 27115 10192 27124
rect 10140 27081 10149 27115
rect 10149 27081 10183 27115
rect 10183 27081 10192 27115
rect 10140 27072 10192 27081
rect 10968 27072 11020 27124
rect 3884 27004 3936 27056
rect 4252 27004 4304 27056
rect 4988 27004 5040 27056
rect 6184 27004 6236 27056
rect 7196 26936 7248 26988
rect 7380 26936 7432 26988
rect 9588 27004 9640 27056
rect 3056 26911 3108 26920
rect 3056 26877 3065 26911
rect 3065 26877 3099 26911
rect 3099 26877 3108 26911
rect 3056 26868 3108 26877
rect 3424 26911 3476 26920
rect 3424 26877 3433 26911
rect 3433 26877 3467 26911
rect 3467 26877 3476 26911
rect 3424 26868 3476 26877
rect 8024 26936 8076 26988
rect 9036 26936 9088 26988
rect 11612 27004 11664 27056
rect 10600 26979 10652 26988
rect 8944 26868 8996 26920
rect 10600 26945 10609 26979
rect 10609 26945 10643 26979
rect 10643 26945 10652 26979
rect 10600 26936 10652 26945
rect 11796 27047 11848 27056
rect 11796 27013 11805 27047
rect 11805 27013 11839 27047
rect 11839 27013 11848 27047
rect 11796 27004 11848 27013
rect 11980 27004 12032 27056
rect 12348 27115 12400 27124
rect 12348 27081 12357 27115
rect 12357 27081 12391 27115
rect 12391 27081 12400 27115
rect 12348 27072 12400 27081
rect 12624 27072 12676 27124
rect 12808 27047 12860 27056
rect 12808 27013 12817 27047
rect 12817 27013 12851 27047
rect 12851 27013 12860 27047
rect 12808 27004 12860 27013
rect 13452 27004 13504 27056
rect 13912 27004 13964 27056
rect 16028 27072 16080 27124
rect 17040 27115 17092 27124
rect 17040 27081 17049 27115
rect 17049 27081 17083 27115
rect 17083 27081 17092 27115
rect 17040 27072 17092 27081
rect 18972 27115 19024 27124
rect 18972 27081 18981 27115
rect 18981 27081 19015 27115
rect 19015 27081 19024 27115
rect 18972 27072 19024 27081
rect 23480 27072 23532 27124
rect 26700 27072 26752 27124
rect 26976 27115 27028 27124
rect 26976 27081 26985 27115
rect 26985 27081 27019 27115
rect 27019 27081 27028 27115
rect 26976 27072 27028 27081
rect 29184 27072 29236 27124
rect 30012 27072 30064 27124
rect 33324 27072 33376 27124
rect 34520 27072 34572 27124
rect 16212 27004 16264 27056
rect 17500 27047 17552 27056
rect 17500 27013 17509 27047
rect 17509 27013 17543 27047
rect 17543 27013 17552 27047
rect 17500 27004 17552 27013
rect 12716 26979 12768 26988
rect 12716 26945 12725 26979
rect 12725 26945 12759 26979
rect 12759 26945 12768 26979
rect 12716 26936 12768 26945
rect 12992 26979 13044 26988
rect 12992 26945 13000 26979
rect 13000 26945 13034 26979
rect 13034 26945 13044 26979
rect 12992 26936 13044 26945
rect 13084 26979 13136 26988
rect 13084 26945 13093 26979
rect 13093 26945 13127 26979
rect 13127 26945 13136 26979
rect 13084 26936 13136 26945
rect 14556 26936 14608 26988
rect 14832 26979 14884 26988
rect 14832 26945 14841 26979
rect 14841 26945 14875 26979
rect 14875 26945 14884 26979
rect 14832 26936 14884 26945
rect 16580 26936 16632 26988
rect 17316 26979 17368 26988
rect 17316 26945 17323 26979
rect 17323 26945 17368 26979
rect 17316 26936 17368 26945
rect 17408 26979 17460 26988
rect 17408 26945 17417 26979
rect 17417 26945 17451 26979
rect 17451 26945 17460 26979
rect 17408 26936 17460 26945
rect 10416 26868 10468 26920
rect 9128 26800 9180 26852
rect 3700 26732 3752 26784
rect 4528 26732 4580 26784
rect 4712 26732 4764 26784
rect 4988 26775 5040 26784
rect 4988 26741 4997 26775
rect 4997 26741 5031 26775
rect 5031 26741 5040 26775
rect 4988 26732 5040 26741
rect 9772 26732 9824 26784
rect 10508 26732 10560 26784
rect 13360 26911 13412 26920
rect 13360 26877 13369 26911
rect 13369 26877 13403 26911
rect 13403 26877 13412 26911
rect 13360 26868 13412 26877
rect 17040 26868 17092 26920
rect 18052 26936 18104 26988
rect 19800 26936 19852 26988
rect 19984 26979 20036 26988
rect 19984 26945 19993 26979
rect 19993 26945 20027 26979
rect 20027 26945 20036 26979
rect 19984 26936 20036 26945
rect 20168 26979 20220 26988
rect 20168 26945 20177 26979
rect 20177 26945 20211 26979
rect 20211 26945 20220 26979
rect 20168 26936 20220 26945
rect 20536 26979 20588 26988
rect 20536 26945 20545 26979
rect 20545 26945 20579 26979
rect 20579 26945 20588 26979
rect 20536 26936 20588 26945
rect 17960 26911 18012 26920
rect 17960 26877 17969 26911
rect 17969 26877 18003 26911
rect 18003 26877 18012 26911
rect 17960 26868 18012 26877
rect 14740 26800 14792 26852
rect 16396 26800 16448 26852
rect 20260 26911 20312 26920
rect 20260 26877 20269 26911
rect 20269 26877 20303 26911
rect 20303 26877 20312 26911
rect 20260 26868 20312 26877
rect 21824 27047 21876 27056
rect 21824 27013 21833 27047
rect 21833 27013 21867 27047
rect 21867 27013 21876 27047
rect 21824 27004 21876 27013
rect 20996 26868 21048 26920
rect 11152 26732 11204 26784
rect 11520 26775 11572 26784
rect 11520 26741 11529 26775
rect 11529 26741 11563 26775
rect 11563 26741 11572 26775
rect 11520 26732 11572 26741
rect 12348 26732 12400 26784
rect 16764 26732 16816 26784
rect 17776 26775 17828 26784
rect 17776 26741 17785 26775
rect 17785 26741 17819 26775
rect 17819 26741 17828 26775
rect 17776 26732 17828 26741
rect 17868 26732 17920 26784
rect 21824 26800 21876 26852
rect 22284 26911 22336 26920
rect 22284 26877 22293 26911
rect 22293 26877 22327 26911
rect 22327 26877 22336 26911
rect 22836 26936 22888 26988
rect 25504 27047 25556 27056
rect 25504 27013 25513 27047
rect 25513 27013 25547 27047
rect 25547 27013 25556 27047
rect 25504 27004 25556 27013
rect 24124 26936 24176 26988
rect 24584 26936 24636 26988
rect 26332 26936 26384 26988
rect 27344 26936 27396 26988
rect 29644 26979 29696 26988
rect 30104 27004 30156 27056
rect 31760 27047 31812 27056
rect 31760 27013 31769 27047
rect 31769 27013 31803 27047
rect 31803 27013 31812 27047
rect 31760 27004 31812 27013
rect 29644 26945 29662 26979
rect 29662 26945 29696 26979
rect 29644 26936 29696 26945
rect 30380 26936 30432 26988
rect 33968 26979 34020 26988
rect 33968 26945 33977 26979
rect 33977 26945 34011 26979
rect 34011 26945 34020 26979
rect 33968 26936 34020 26945
rect 34244 26979 34296 26988
rect 34244 26945 34253 26979
rect 34253 26945 34287 26979
rect 34287 26945 34296 26979
rect 34244 26936 34296 26945
rect 34520 26979 34572 26988
rect 34520 26945 34529 26979
rect 34529 26945 34563 26979
rect 34563 26945 34572 26979
rect 34520 26936 34572 26945
rect 22284 26868 22336 26877
rect 34796 26911 34848 26920
rect 34796 26877 34805 26911
rect 34805 26877 34839 26911
rect 34839 26877 34848 26911
rect 34796 26868 34848 26877
rect 23664 26775 23716 26784
rect 23664 26741 23673 26775
rect 23673 26741 23707 26775
rect 23707 26741 23716 26775
rect 23664 26732 23716 26741
rect 24216 26732 24268 26784
rect 25412 26775 25464 26784
rect 25412 26741 25421 26775
rect 25421 26741 25455 26775
rect 25455 26741 25464 26775
rect 25412 26732 25464 26741
rect 26332 26775 26384 26784
rect 26332 26741 26341 26775
rect 26341 26741 26375 26775
rect 26375 26741 26384 26775
rect 26332 26732 26384 26741
rect 26608 26732 26660 26784
rect 30288 26732 30340 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 5448 26528 5500 26580
rect 5724 26571 5776 26580
rect 5724 26537 5733 26571
rect 5733 26537 5767 26571
rect 5767 26537 5776 26571
rect 5724 26528 5776 26537
rect 9772 26571 9824 26580
rect 9772 26537 9781 26571
rect 9781 26537 9815 26571
rect 9815 26537 9824 26571
rect 9772 26528 9824 26537
rect 9956 26528 10008 26580
rect 12348 26528 12400 26580
rect 4988 26460 5040 26512
rect 5264 26460 5316 26512
rect 9496 26460 9548 26512
rect 11704 26503 11756 26512
rect 11704 26469 11713 26503
rect 11713 26469 11747 26503
rect 11747 26469 11756 26503
rect 11704 26460 11756 26469
rect 12716 26528 12768 26580
rect 15108 26571 15160 26580
rect 15108 26537 15117 26571
rect 15117 26537 15151 26571
rect 15151 26537 15160 26571
rect 15108 26528 15160 26537
rect 15384 26528 15436 26580
rect 16488 26528 16540 26580
rect 11336 26435 11388 26444
rect 11336 26401 11345 26435
rect 11345 26401 11379 26435
rect 11379 26401 11388 26435
rect 11336 26392 11388 26401
rect 1308 26324 1360 26376
rect 3884 26324 3936 26376
rect 5724 26324 5776 26376
rect 11520 26367 11572 26376
rect 11520 26333 11529 26367
rect 11529 26333 11563 26367
rect 11563 26333 11572 26367
rect 11520 26324 11572 26333
rect 13360 26324 13412 26376
rect 13728 26324 13780 26376
rect 1860 26299 1912 26308
rect 1860 26265 1869 26299
rect 1869 26265 1903 26299
rect 1903 26265 1912 26299
rect 1860 26256 1912 26265
rect 3700 26256 3752 26308
rect 3056 26188 3108 26240
rect 4252 26188 4304 26240
rect 6552 26188 6604 26240
rect 7748 26188 7800 26240
rect 8576 26188 8628 26240
rect 9404 26188 9456 26240
rect 10600 26256 10652 26308
rect 12532 26256 12584 26308
rect 14464 26256 14516 26308
rect 15936 26324 15988 26376
rect 16028 26324 16080 26376
rect 16856 26367 16908 26376
rect 16856 26333 16866 26367
rect 16866 26333 16900 26367
rect 16900 26333 16908 26367
rect 16856 26324 16908 26333
rect 17132 26460 17184 26512
rect 17132 26367 17184 26376
rect 17132 26333 17141 26367
rect 17141 26333 17175 26367
rect 17175 26333 17184 26367
rect 17132 26324 17184 26333
rect 17408 26503 17460 26512
rect 17408 26469 17417 26503
rect 17417 26469 17451 26503
rect 17451 26469 17460 26503
rect 17408 26460 17460 26469
rect 17684 26571 17736 26580
rect 17684 26537 17693 26571
rect 17693 26537 17727 26571
rect 17727 26537 17736 26571
rect 17684 26528 17736 26537
rect 20260 26528 20312 26580
rect 21456 26571 21508 26580
rect 21456 26537 21465 26571
rect 21465 26537 21499 26571
rect 21499 26537 21508 26571
rect 21456 26528 21508 26537
rect 17776 26460 17828 26512
rect 19984 26460 20036 26512
rect 21824 26528 21876 26580
rect 22836 26571 22888 26580
rect 22836 26537 22845 26571
rect 22845 26537 22879 26571
rect 22879 26537 22888 26571
rect 22836 26528 22888 26537
rect 22928 26528 22980 26580
rect 20260 26392 20312 26444
rect 22376 26460 22428 26512
rect 24584 26571 24636 26580
rect 24584 26537 24593 26571
rect 24593 26537 24627 26571
rect 24627 26537 24636 26571
rect 24584 26528 24636 26537
rect 26240 26528 26292 26580
rect 27344 26571 27396 26580
rect 27344 26537 27353 26571
rect 27353 26537 27387 26571
rect 27387 26537 27396 26571
rect 27344 26528 27396 26537
rect 33968 26528 34020 26580
rect 22008 26435 22060 26444
rect 22008 26401 22017 26435
rect 22017 26401 22051 26435
rect 22051 26401 22060 26435
rect 22008 26392 22060 26401
rect 22744 26435 22796 26444
rect 22744 26401 22753 26435
rect 22753 26401 22787 26435
rect 22787 26401 22796 26435
rect 25412 26460 25464 26512
rect 25504 26460 25556 26512
rect 22744 26392 22796 26401
rect 17592 26367 17644 26376
rect 17592 26333 17601 26367
rect 17601 26333 17635 26367
rect 17635 26333 17644 26367
rect 17592 26324 17644 26333
rect 18052 26367 18104 26376
rect 18052 26333 18061 26367
rect 18061 26333 18095 26367
rect 18095 26333 18104 26367
rect 18052 26324 18104 26333
rect 18236 26367 18288 26376
rect 18236 26333 18245 26367
rect 18245 26333 18279 26367
rect 18279 26333 18288 26367
rect 18236 26324 18288 26333
rect 21640 26324 21692 26376
rect 15016 26256 15068 26308
rect 15844 26256 15896 26308
rect 10416 26188 10468 26240
rect 13084 26188 13136 26240
rect 13636 26231 13688 26240
rect 13636 26197 13645 26231
rect 13645 26197 13679 26231
rect 13679 26197 13688 26231
rect 13636 26188 13688 26197
rect 14096 26188 14148 26240
rect 15108 26188 15160 26240
rect 16396 26188 16448 26240
rect 18144 26256 18196 26308
rect 23664 26324 23716 26376
rect 21548 26188 21600 26240
rect 21732 26188 21784 26240
rect 22100 26188 22152 26240
rect 23480 26256 23532 26308
rect 23848 26256 23900 26308
rect 25596 26324 25648 26376
rect 25964 26460 26016 26512
rect 27436 26460 27488 26512
rect 26700 26435 26752 26444
rect 26700 26401 26709 26435
rect 26709 26401 26743 26435
rect 26743 26401 26752 26435
rect 26700 26392 26752 26401
rect 27620 26392 27672 26444
rect 26240 26367 26292 26376
rect 26240 26333 26249 26367
rect 26249 26333 26283 26367
rect 26283 26333 26292 26367
rect 26240 26324 26292 26333
rect 26516 26324 26568 26376
rect 26976 26367 27028 26376
rect 26976 26333 26985 26367
rect 26985 26333 27019 26367
rect 27019 26333 27028 26367
rect 26976 26324 27028 26333
rect 28724 26324 28776 26376
rect 28908 26435 28960 26444
rect 28908 26401 28917 26435
rect 28917 26401 28951 26435
rect 28951 26401 28960 26435
rect 28908 26392 28960 26401
rect 29184 26367 29236 26376
rect 29184 26333 29193 26367
rect 29193 26333 29227 26367
rect 29227 26333 29236 26367
rect 29184 26324 29236 26333
rect 30104 26435 30156 26444
rect 30104 26401 30113 26435
rect 30113 26401 30147 26435
rect 30147 26401 30156 26435
rect 30104 26392 30156 26401
rect 31116 26324 31168 26376
rect 31852 26324 31904 26376
rect 34244 26367 34296 26376
rect 34244 26333 34253 26367
rect 34253 26333 34287 26367
rect 34287 26333 34296 26367
rect 34244 26324 34296 26333
rect 25964 26256 26016 26308
rect 30472 26256 30524 26308
rect 34520 26256 34572 26308
rect 34980 26256 35032 26308
rect 23756 26188 23808 26240
rect 25320 26188 25372 26240
rect 26056 26231 26108 26240
rect 26056 26197 26065 26231
rect 26065 26197 26099 26231
rect 26099 26197 26108 26231
rect 26056 26188 26108 26197
rect 31484 26231 31536 26240
rect 31484 26197 31493 26231
rect 31493 26197 31527 26231
rect 31527 26197 31536 26231
rect 31484 26188 31536 26197
rect 33784 26231 33836 26240
rect 33784 26197 33793 26231
rect 33793 26197 33827 26231
rect 33827 26197 33836 26231
rect 33784 26188 33836 26197
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 4712 25984 4764 26036
rect 4068 25916 4120 25968
rect 4804 25891 4856 25900
rect 4804 25857 4813 25891
rect 4813 25857 4847 25891
rect 4847 25857 4856 25891
rect 4804 25848 4856 25857
rect 5540 25916 5592 25968
rect 4712 25780 4764 25832
rect 5172 25891 5224 25900
rect 5172 25857 5181 25891
rect 5181 25857 5215 25891
rect 5215 25857 5224 25891
rect 5172 25848 5224 25857
rect 5448 25848 5500 25900
rect 4252 25712 4304 25764
rect 5448 25712 5500 25764
rect 3608 25687 3660 25696
rect 3608 25653 3617 25687
rect 3617 25653 3651 25687
rect 3651 25653 3660 25687
rect 3608 25644 3660 25653
rect 5632 25644 5684 25696
rect 5816 25780 5868 25832
rect 7288 25848 7340 25900
rect 8208 25848 8260 25900
rect 8576 25891 8628 25900
rect 8576 25857 8585 25891
rect 8585 25857 8619 25891
rect 8619 25857 8628 25891
rect 8576 25848 8628 25857
rect 9680 25916 9732 25968
rect 10600 26027 10652 26036
rect 10600 25993 10609 26027
rect 10609 25993 10643 26027
rect 10643 25993 10652 26027
rect 10600 25984 10652 25993
rect 12532 26027 12584 26036
rect 12532 25993 12541 26027
rect 12541 25993 12575 26027
rect 12575 25993 12584 26027
rect 12532 25984 12584 25993
rect 12716 25984 12768 26036
rect 13268 25984 13320 26036
rect 15384 25984 15436 26036
rect 15660 26027 15712 26036
rect 15660 25993 15669 26027
rect 15669 25993 15703 26027
rect 15703 25993 15712 26027
rect 15660 25984 15712 25993
rect 16396 26027 16448 26036
rect 16396 25993 16405 26027
rect 16405 25993 16439 26027
rect 16439 25993 16448 26027
rect 16396 25984 16448 25993
rect 16856 25984 16908 26036
rect 20076 25984 20128 26036
rect 20168 25984 20220 26036
rect 20444 25984 20496 26036
rect 22744 25984 22796 26036
rect 23204 25984 23256 26036
rect 9496 25848 9548 25900
rect 11336 25916 11388 25968
rect 12900 25959 12952 25968
rect 12900 25925 12909 25959
rect 12909 25925 12943 25959
rect 12943 25925 12952 25959
rect 12900 25916 12952 25925
rect 10140 25848 10192 25900
rect 6552 25823 6604 25832
rect 6552 25789 6561 25823
rect 6561 25789 6595 25823
rect 6595 25789 6604 25823
rect 6552 25780 6604 25789
rect 8300 25780 8352 25832
rect 9772 25780 9824 25832
rect 10324 25891 10376 25900
rect 10324 25857 10333 25891
rect 10333 25857 10367 25891
rect 10367 25857 10376 25891
rect 10324 25848 10376 25857
rect 10416 25848 10468 25900
rect 13728 25848 13780 25900
rect 14832 25916 14884 25968
rect 16488 25916 16540 25968
rect 14648 25848 14700 25900
rect 16396 25848 16448 25900
rect 10968 25823 11020 25832
rect 10968 25789 10977 25823
rect 10977 25789 11011 25823
rect 11011 25789 11020 25823
rect 10968 25780 11020 25789
rect 13268 25780 13320 25832
rect 15108 25780 15160 25832
rect 17224 25848 17276 25900
rect 18052 25823 18104 25832
rect 18052 25789 18061 25823
rect 18061 25789 18095 25823
rect 18095 25789 18104 25823
rect 18052 25780 18104 25789
rect 11704 25712 11756 25764
rect 6184 25644 6236 25696
rect 7564 25687 7616 25696
rect 7564 25653 7573 25687
rect 7573 25653 7607 25687
rect 7607 25653 7616 25687
rect 7564 25644 7616 25653
rect 7656 25644 7708 25696
rect 8760 25687 8812 25696
rect 8760 25653 8769 25687
rect 8769 25653 8803 25687
rect 8803 25653 8812 25687
rect 8760 25644 8812 25653
rect 8852 25687 8904 25696
rect 8852 25653 8861 25687
rect 8861 25653 8895 25687
rect 8895 25653 8904 25687
rect 8852 25644 8904 25653
rect 9128 25644 9180 25696
rect 9864 25644 9916 25696
rect 10508 25644 10560 25696
rect 15568 25644 15620 25696
rect 16120 25644 16172 25696
rect 18328 25687 18380 25696
rect 18328 25653 18337 25687
rect 18337 25653 18371 25687
rect 18371 25653 18380 25687
rect 18328 25644 18380 25653
rect 19064 25848 19116 25900
rect 19616 25891 19668 25900
rect 19616 25857 19625 25891
rect 19625 25857 19659 25891
rect 19659 25857 19668 25891
rect 19616 25848 19668 25857
rect 20628 25916 20680 25968
rect 19984 25891 20036 25900
rect 19984 25857 19993 25891
rect 19993 25857 20027 25891
rect 20027 25857 20036 25891
rect 19984 25848 20036 25857
rect 21916 25891 21968 25900
rect 21916 25857 21925 25891
rect 21925 25857 21959 25891
rect 21959 25857 21968 25891
rect 21916 25848 21968 25857
rect 23020 25916 23072 25968
rect 23572 25848 23624 25900
rect 24124 25848 24176 25900
rect 24860 25848 24912 25900
rect 18880 25823 18932 25832
rect 18880 25789 18889 25823
rect 18889 25789 18923 25823
rect 18923 25789 18932 25823
rect 18880 25780 18932 25789
rect 21732 25780 21784 25832
rect 26516 26027 26568 26036
rect 26516 25993 26525 26027
rect 26525 25993 26559 26027
rect 26559 25993 26568 26027
rect 26516 25984 26568 25993
rect 28172 25984 28224 26036
rect 27252 25848 27304 25900
rect 30472 25984 30524 26036
rect 30748 25984 30800 26036
rect 31484 25984 31536 26036
rect 33600 25984 33652 26036
rect 33784 25916 33836 25968
rect 34980 26027 35032 26036
rect 34980 25993 34989 26027
rect 34989 25993 35023 26027
rect 35023 25993 35032 26027
rect 34980 25984 35032 25993
rect 33968 25916 34020 25968
rect 30104 25780 30156 25832
rect 30656 25780 30708 25832
rect 32772 25780 32824 25832
rect 25320 25712 25372 25764
rect 29000 25712 29052 25764
rect 20628 25644 20680 25696
rect 22100 25687 22152 25696
rect 22100 25653 22109 25687
rect 22109 25653 22143 25687
rect 22143 25653 22152 25687
rect 22100 25644 22152 25653
rect 22468 25687 22520 25696
rect 22468 25653 22477 25687
rect 22477 25653 22511 25687
rect 22511 25653 22520 25687
rect 22468 25644 22520 25653
rect 25228 25644 25280 25696
rect 25596 25644 25648 25696
rect 31024 25644 31076 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 5172 25440 5224 25492
rect 8208 25483 8260 25492
rect 8208 25449 8217 25483
rect 8217 25449 8251 25483
rect 8251 25449 8260 25483
rect 8208 25440 8260 25449
rect 9496 25483 9548 25492
rect 9496 25449 9505 25483
rect 9505 25449 9539 25483
rect 9539 25449 9548 25483
rect 9496 25440 9548 25449
rect 3424 25304 3476 25356
rect 7564 25236 7616 25288
rect 9404 25372 9456 25424
rect 12716 25440 12768 25492
rect 12992 25483 13044 25492
rect 12992 25449 13001 25483
rect 13001 25449 13035 25483
rect 13035 25449 13044 25483
rect 12992 25440 13044 25449
rect 14648 25483 14700 25492
rect 14648 25449 14657 25483
rect 14657 25449 14691 25483
rect 14691 25449 14700 25483
rect 14648 25440 14700 25449
rect 16028 25483 16080 25492
rect 16028 25449 16037 25483
rect 16037 25449 16071 25483
rect 16071 25449 16080 25483
rect 16028 25440 16080 25449
rect 16304 25483 16356 25492
rect 16304 25449 16313 25483
rect 16313 25449 16347 25483
rect 16347 25449 16356 25483
rect 16304 25440 16356 25449
rect 17224 25440 17276 25492
rect 8760 25304 8812 25356
rect 4528 25168 4580 25220
rect 6368 25168 6420 25220
rect 9772 25236 9824 25288
rect 11704 25236 11756 25288
rect 14004 25236 14056 25288
rect 15200 25304 15252 25356
rect 16028 25304 16080 25356
rect 15108 25236 15160 25288
rect 15568 25236 15620 25288
rect 9128 25211 9180 25220
rect 9128 25177 9137 25211
rect 9137 25177 9171 25211
rect 9171 25177 9180 25211
rect 9128 25168 9180 25177
rect 10140 25168 10192 25220
rect 6736 25143 6788 25152
rect 6736 25109 6745 25143
rect 6745 25109 6779 25143
rect 6779 25109 6788 25143
rect 6736 25100 6788 25109
rect 8300 25100 8352 25152
rect 10968 25168 11020 25220
rect 12164 25168 12216 25220
rect 15660 25211 15712 25220
rect 15660 25177 15669 25211
rect 15669 25177 15703 25211
rect 15703 25177 15712 25211
rect 15660 25168 15712 25177
rect 10324 25100 10376 25152
rect 14924 25100 14976 25152
rect 16488 25372 16540 25424
rect 18052 25440 18104 25492
rect 19064 25483 19116 25492
rect 19064 25449 19073 25483
rect 19073 25449 19107 25483
rect 19107 25449 19116 25483
rect 19064 25440 19116 25449
rect 19156 25440 19208 25492
rect 16580 25347 16632 25356
rect 16580 25313 16589 25347
rect 16589 25313 16623 25347
rect 16623 25313 16632 25347
rect 16580 25304 16632 25313
rect 16856 25304 16908 25356
rect 22100 25372 22152 25424
rect 24860 25483 24912 25492
rect 24860 25449 24869 25483
rect 24869 25449 24903 25483
rect 24903 25449 24912 25483
rect 24860 25440 24912 25449
rect 25780 25440 25832 25492
rect 27252 25440 27304 25492
rect 22192 25304 22244 25356
rect 22468 25304 22520 25356
rect 16764 25279 16816 25288
rect 16764 25245 16773 25279
rect 16773 25245 16807 25279
rect 16807 25245 16816 25279
rect 16764 25236 16816 25245
rect 18328 25236 18380 25288
rect 18972 25236 19024 25288
rect 20444 25236 20496 25288
rect 22284 25236 22336 25288
rect 22560 25279 22612 25288
rect 22560 25245 22569 25279
rect 22569 25245 22603 25279
rect 22603 25245 22612 25279
rect 22560 25236 22612 25245
rect 19708 25168 19760 25220
rect 21824 25168 21876 25220
rect 23112 25168 23164 25220
rect 23756 25168 23808 25220
rect 16304 25100 16356 25152
rect 16580 25100 16632 25152
rect 17500 25100 17552 25152
rect 19984 25100 20036 25152
rect 22284 25143 22336 25152
rect 22284 25109 22293 25143
rect 22293 25109 22327 25143
rect 22327 25109 22336 25143
rect 22284 25100 22336 25109
rect 23940 25143 23992 25152
rect 23940 25109 23949 25143
rect 23949 25109 23983 25143
rect 23983 25109 23992 25143
rect 23940 25100 23992 25109
rect 24584 25100 24636 25152
rect 24952 25236 25004 25288
rect 25228 25211 25280 25220
rect 25228 25177 25237 25211
rect 25237 25177 25271 25211
rect 25271 25177 25280 25211
rect 25228 25168 25280 25177
rect 26976 25168 27028 25220
rect 27988 25279 28040 25288
rect 27988 25245 27997 25279
rect 27997 25245 28031 25279
rect 28031 25245 28040 25279
rect 27988 25236 28040 25245
rect 30656 25440 30708 25492
rect 30932 25440 30984 25492
rect 30196 25347 30248 25356
rect 30196 25313 30205 25347
rect 30205 25313 30239 25347
rect 30239 25313 30248 25347
rect 31300 25372 31352 25424
rect 30196 25304 30248 25313
rect 30564 25304 30616 25356
rect 28080 25168 28132 25220
rect 30748 25279 30800 25288
rect 30748 25245 30757 25279
rect 30757 25245 30791 25279
rect 30791 25245 30800 25279
rect 30748 25236 30800 25245
rect 31024 25236 31076 25288
rect 25320 25143 25372 25152
rect 25320 25109 25329 25143
rect 25329 25109 25363 25143
rect 25363 25109 25372 25143
rect 25320 25100 25372 25109
rect 25688 25143 25740 25152
rect 25688 25109 25697 25143
rect 25697 25109 25731 25143
rect 25731 25109 25740 25143
rect 25688 25100 25740 25109
rect 26240 25143 26292 25152
rect 26240 25109 26249 25143
rect 26249 25109 26283 25143
rect 26283 25109 26292 25143
rect 26240 25100 26292 25109
rect 27344 25100 27396 25152
rect 30104 25100 30156 25152
rect 30840 25100 30892 25152
rect 31300 25143 31352 25152
rect 31300 25109 31309 25143
rect 31309 25109 31343 25143
rect 31343 25109 31352 25143
rect 31300 25100 31352 25109
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 4160 24896 4212 24948
rect 4528 24939 4580 24948
rect 4528 24905 4537 24939
rect 4537 24905 4571 24939
rect 4571 24905 4580 24939
rect 4528 24896 4580 24905
rect 5264 24896 5316 24948
rect 6368 24939 6420 24948
rect 6368 24905 6377 24939
rect 6377 24905 6411 24939
rect 6411 24905 6420 24939
rect 6368 24896 6420 24905
rect 6736 24939 6788 24948
rect 6736 24905 6745 24939
rect 6745 24905 6779 24939
rect 6779 24905 6788 24939
rect 6736 24896 6788 24905
rect 9680 24939 9732 24948
rect 9680 24905 9689 24939
rect 9689 24905 9723 24939
rect 9723 24905 9732 24939
rect 9680 24896 9732 24905
rect 10140 24939 10192 24948
rect 10140 24905 10149 24939
rect 10149 24905 10183 24939
rect 10183 24905 10192 24939
rect 10140 24896 10192 24905
rect 10324 24896 10376 24948
rect 11060 24939 11112 24948
rect 11060 24905 11069 24939
rect 11069 24905 11103 24939
rect 11103 24905 11112 24939
rect 11060 24896 11112 24905
rect 14924 24896 14976 24948
rect 15108 24939 15160 24948
rect 15108 24905 15117 24939
rect 15117 24905 15151 24939
rect 15151 24905 15160 24939
rect 15108 24896 15160 24905
rect 16120 24896 16172 24948
rect 19524 24896 19576 24948
rect 19708 24939 19760 24948
rect 19708 24905 19717 24939
rect 19717 24905 19751 24939
rect 19751 24905 19760 24939
rect 19708 24896 19760 24905
rect 19984 24896 20036 24948
rect 21824 24939 21876 24948
rect 21824 24905 21833 24939
rect 21833 24905 21867 24939
rect 21867 24905 21876 24939
rect 21824 24896 21876 24905
rect 22284 24896 22336 24948
rect 23112 24939 23164 24948
rect 23112 24905 23121 24939
rect 23121 24905 23155 24939
rect 23155 24905 23164 24939
rect 23112 24896 23164 24905
rect 3424 24828 3476 24880
rect 8852 24828 8904 24880
rect 3608 24760 3660 24812
rect 5448 24760 5500 24812
rect 5632 24692 5684 24744
rect 3884 24624 3936 24676
rect 7288 24692 7340 24744
rect 10968 24828 11020 24880
rect 13268 24828 13320 24880
rect 15016 24828 15068 24880
rect 12532 24760 12584 24812
rect 12900 24760 12952 24812
rect 13636 24803 13688 24812
rect 13636 24769 13645 24803
rect 13645 24769 13679 24803
rect 13679 24769 13688 24803
rect 13636 24760 13688 24769
rect 13728 24803 13780 24812
rect 13728 24769 13737 24803
rect 13737 24769 13771 24803
rect 13771 24769 13780 24803
rect 13728 24760 13780 24769
rect 11060 24692 11112 24744
rect 10048 24624 10100 24676
rect 9772 24556 9824 24608
rect 10232 24556 10284 24608
rect 11704 24556 11756 24608
rect 14096 24556 14148 24608
rect 14372 24556 14424 24608
rect 15476 24556 15528 24608
rect 16672 24599 16724 24608
rect 16672 24565 16681 24599
rect 16681 24565 16715 24599
rect 16715 24565 16724 24599
rect 16672 24556 16724 24565
rect 17132 24803 17184 24812
rect 17132 24769 17141 24803
rect 17141 24769 17175 24803
rect 17175 24769 17184 24803
rect 17132 24760 17184 24769
rect 19800 24828 19852 24880
rect 23664 24896 23716 24948
rect 25780 24896 25832 24948
rect 26976 24939 27028 24948
rect 26976 24905 26985 24939
rect 26985 24905 27019 24939
rect 27019 24905 27028 24939
rect 26976 24896 27028 24905
rect 27344 24939 27396 24948
rect 27344 24905 27353 24939
rect 27353 24905 27387 24939
rect 27387 24905 27396 24939
rect 27344 24896 27396 24905
rect 20076 24760 20128 24812
rect 21640 24760 21692 24812
rect 22928 24803 22980 24812
rect 22928 24769 22937 24803
rect 22937 24769 22971 24803
rect 22971 24769 22980 24803
rect 22928 24760 22980 24769
rect 23020 24760 23072 24812
rect 24032 24803 24084 24812
rect 24032 24769 24042 24803
rect 24042 24769 24076 24803
rect 24076 24769 24084 24803
rect 24032 24760 24084 24769
rect 24308 24803 24360 24812
rect 24308 24769 24317 24803
rect 24317 24769 24351 24803
rect 24351 24769 24360 24803
rect 24308 24760 24360 24769
rect 25596 24828 25648 24880
rect 26240 24828 26292 24880
rect 28080 24896 28132 24948
rect 28448 24896 28500 24948
rect 29184 24896 29236 24948
rect 30104 24939 30156 24948
rect 30104 24905 30113 24939
rect 30113 24905 30147 24939
rect 30147 24905 30156 24939
rect 30104 24896 30156 24905
rect 17224 24735 17276 24744
rect 17224 24701 17233 24735
rect 17233 24701 17267 24735
rect 17267 24701 17276 24735
rect 17224 24692 17276 24701
rect 17316 24692 17368 24744
rect 18328 24624 18380 24676
rect 20076 24624 20128 24676
rect 20352 24735 20404 24744
rect 20352 24701 20361 24735
rect 20361 24701 20395 24735
rect 20395 24701 20404 24735
rect 20352 24692 20404 24701
rect 22100 24692 22152 24744
rect 22468 24692 22520 24744
rect 17592 24556 17644 24608
rect 19984 24556 20036 24608
rect 20168 24556 20220 24608
rect 22376 24556 22428 24608
rect 22928 24624 22980 24676
rect 23572 24735 23624 24744
rect 23572 24701 23581 24735
rect 23581 24701 23615 24735
rect 23615 24701 23624 24735
rect 23572 24692 23624 24701
rect 23756 24735 23808 24744
rect 23756 24701 23765 24735
rect 23765 24701 23799 24735
rect 23799 24701 23808 24735
rect 23756 24692 23808 24701
rect 24768 24760 24820 24812
rect 25780 24760 25832 24812
rect 27252 24760 27304 24812
rect 26884 24692 26936 24744
rect 26976 24692 27028 24744
rect 27620 24828 27672 24880
rect 28540 24760 28592 24812
rect 29736 24760 29788 24812
rect 30012 24760 30064 24812
rect 30288 24760 30340 24812
rect 30840 24803 30892 24812
rect 30840 24769 30849 24803
rect 30849 24769 30883 24803
rect 30883 24769 30892 24803
rect 30840 24760 30892 24769
rect 31760 24760 31812 24812
rect 27620 24692 27672 24744
rect 28724 24692 28776 24744
rect 28908 24692 28960 24744
rect 22652 24556 22704 24608
rect 23204 24556 23256 24608
rect 24032 24556 24084 24608
rect 26056 24624 26108 24676
rect 26148 24556 26200 24608
rect 26240 24599 26292 24608
rect 26240 24565 26249 24599
rect 26249 24565 26283 24599
rect 26283 24565 26292 24599
rect 26240 24556 26292 24565
rect 31116 24692 31168 24744
rect 27068 24556 27120 24608
rect 28080 24556 28132 24608
rect 28172 24599 28224 24608
rect 28172 24565 28181 24599
rect 28181 24565 28215 24599
rect 28215 24565 28224 24599
rect 28172 24556 28224 24565
rect 28356 24599 28408 24608
rect 28356 24565 28365 24599
rect 28365 24565 28399 24599
rect 28399 24565 28408 24599
rect 28356 24556 28408 24565
rect 28816 24599 28868 24608
rect 28816 24565 28825 24599
rect 28825 24565 28859 24599
rect 28859 24565 28868 24599
rect 28816 24556 28868 24565
rect 29736 24599 29788 24608
rect 29736 24565 29745 24599
rect 29745 24565 29779 24599
rect 29779 24565 29788 24599
rect 29736 24556 29788 24565
rect 31392 24599 31444 24608
rect 31392 24565 31401 24599
rect 31401 24565 31435 24599
rect 31435 24565 31444 24599
rect 31392 24556 31444 24565
rect 31484 24599 31536 24608
rect 31484 24565 31493 24599
rect 31493 24565 31527 24599
rect 31527 24565 31536 24599
rect 31484 24556 31536 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 10048 24395 10100 24404
rect 10048 24361 10057 24395
rect 10057 24361 10091 24395
rect 10091 24361 10100 24395
rect 10048 24352 10100 24361
rect 12164 24395 12216 24404
rect 12164 24361 12173 24395
rect 12173 24361 12207 24395
rect 12207 24361 12216 24395
rect 12164 24352 12216 24361
rect 14188 24395 14240 24404
rect 14188 24361 14197 24395
rect 14197 24361 14231 24395
rect 14231 24361 14240 24395
rect 14188 24352 14240 24361
rect 5448 24284 5500 24336
rect 11152 24284 11204 24336
rect 12256 24284 12308 24336
rect 1216 24148 1268 24200
rect 9680 24216 9732 24268
rect 11060 24216 11112 24268
rect 12716 24216 12768 24268
rect 13176 24284 13228 24336
rect 16580 24352 16632 24404
rect 17132 24352 17184 24404
rect 19616 24352 19668 24404
rect 19892 24395 19944 24404
rect 19892 24361 19901 24395
rect 19901 24361 19935 24395
rect 19935 24361 19944 24395
rect 19892 24352 19944 24361
rect 19984 24352 20036 24404
rect 19524 24284 19576 24336
rect 21732 24327 21784 24336
rect 21732 24293 21741 24327
rect 21741 24293 21775 24327
rect 21775 24293 21784 24327
rect 21732 24284 21784 24293
rect 12900 24216 12952 24268
rect 13544 24216 13596 24268
rect 3424 24080 3476 24132
rect 3884 24080 3936 24132
rect 9772 24148 9824 24200
rect 8300 24080 8352 24132
rect 12532 24191 12584 24200
rect 12532 24157 12541 24191
rect 12541 24157 12575 24191
rect 12575 24157 12584 24191
rect 12532 24148 12584 24157
rect 12992 24148 13044 24200
rect 15936 24191 15988 24200
rect 15936 24157 15945 24191
rect 15945 24157 15979 24191
rect 15979 24157 15988 24191
rect 15936 24148 15988 24157
rect 17500 24216 17552 24268
rect 22008 24216 22060 24268
rect 22284 24216 22336 24268
rect 22468 24352 22520 24404
rect 23756 24352 23808 24404
rect 24492 24352 24544 24404
rect 25688 24352 25740 24404
rect 23020 24284 23072 24336
rect 23204 24327 23256 24336
rect 23204 24293 23213 24327
rect 23213 24293 23247 24327
rect 23247 24293 23256 24327
rect 23204 24284 23256 24293
rect 25688 24216 25740 24268
rect 6092 24055 6144 24064
rect 6092 24021 6101 24055
rect 6101 24021 6135 24055
rect 6135 24021 6144 24055
rect 6092 24012 6144 24021
rect 6460 24055 6512 24064
rect 6460 24021 6469 24055
rect 6469 24021 6503 24055
rect 6503 24021 6512 24055
rect 6460 24012 6512 24021
rect 6644 24012 6696 24064
rect 13452 24080 13504 24132
rect 16672 24080 16724 24132
rect 19248 24191 19300 24200
rect 19248 24157 19257 24191
rect 19257 24157 19291 24191
rect 19291 24157 19300 24191
rect 19248 24148 19300 24157
rect 12440 24012 12492 24064
rect 13636 24012 13688 24064
rect 19524 24123 19576 24132
rect 19524 24089 19533 24123
rect 19533 24089 19567 24123
rect 19567 24089 19576 24123
rect 19524 24080 19576 24089
rect 20076 24191 20128 24200
rect 20076 24157 20085 24191
rect 20085 24157 20119 24191
rect 20119 24157 20128 24191
rect 20076 24148 20128 24157
rect 20168 24123 20220 24132
rect 20168 24089 20177 24123
rect 20177 24089 20211 24123
rect 20211 24089 20220 24123
rect 20168 24080 20220 24089
rect 19892 24012 19944 24064
rect 22100 24191 22152 24200
rect 22100 24157 22109 24191
rect 22109 24157 22143 24191
rect 22143 24157 22152 24191
rect 22100 24148 22152 24157
rect 22928 24148 22980 24200
rect 23112 24148 23164 24200
rect 23296 24191 23348 24200
rect 23296 24157 23305 24191
rect 23305 24157 23339 24191
rect 23339 24157 23348 24191
rect 23296 24148 23348 24157
rect 23480 24191 23532 24200
rect 23480 24157 23489 24191
rect 23489 24157 23523 24191
rect 23523 24157 23532 24191
rect 23480 24148 23532 24157
rect 23756 24148 23808 24200
rect 23848 24148 23900 24200
rect 22652 24080 22704 24132
rect 23204 24012 23256 24064
rect 23572 24012 23624 24064
rect 25320 24148 25372 24200
rect 26240 24284 26292 24336
rect 26884 24395 26936 24404
rect 26884 24361 26893 24395
rect 26893 24361 26927 24395
rect 26927 24361 26936 24395
rect 26884 24352 26936 24361
rect 27252 24352 27304 24404
rect 28080 24352 28132 24404
rect 28448 24352 28500 24404
rect 28540 24395 28592 24404
rect 28540 24361 28549 24395
rect 28549 24361 28583 24395
rect 28583 24361 28592 24395
rect 28540 24352 28592 24361
rect 28724 24395 28776 24404
rect 28724 24361 28733 24395
rect 28733 24361 28767 24395
rect 28767 24361 28776 24395
rect 28724 24352 28776 24361
rect 29276 24352 29328 24404
rect 30564 24352 30616 24404
rect 31760 24395 31812 24404
rect 31760 24361 31769 24395
rect 31769 24361 31803 24395
rect 31803 24361 31812 24395
rect 31760 24352 31812 24361
rect 25964 24191 26016 24200
rect 25964 24157 25971 24191
rect 25971 24157 26016 24191
rect 25964 24148 26016 24157
rect 26148 24216 26200 24268
rect 29000 24284 29052 24336
rect 26240 24191 26292 24200
rect 26240 24157 26254 24191
rect 26254 24157 26288 24191
rect 26288 24157 26292 24191
rect 26240 24148 26292 24157
rect 26516 24191 26568 24200
rect 26516 24157 26525 24191
rect 26525 24157 26559 24191
rect 26559 24157 26568 24191
rect 26516 24148 26568 24157
rect 27068 24191 27120 24200
rect 27068 24157 27072 24191
rect 27072 24157 27106 24191
rect 27106 24157 27120 24191
rect 27068 24148 27120 24157
rect 27252 24191 27304 24200
rect 27252 24157 27261 24191
rect 27261 24157 27295 24191
rect 27295 24157 27304 24191
rect 27252 24148 27304 24157
rect 27344 24191 27396 24200
rect 28172 24216 28224 24268
rect 27344 24157 27389 24191
rect 27389 24157 27396 24191
rect 27344 24148 27396 24157
rect 27620 24191 27672 24200
rect 27620 24157 27629 24191
rect 27629 24157 27663 24191
rect 27663 24157 27672 24191
rect 27620 24148 27672 24157
rect 27804 24148 27856 24200
rect 28080 24148 28132 24200
rect 28724 24148 28776 24200
rect 28908 24191 28960 24200
rect 28908 24157 28917 24191
rect 28917 24157 28951 24191
rect 28951 24157 28960 24191
rect 28908 24148 28960 24157
rect 29644 24191 29696 24200
rect 29644 24157 29653 24191
rect 29653 24157 29687 24191
rect 29687 24157 29696 24191
rect 29644 24148 29696 24157
rect 32772 24191 32824 24200
rect 24032 24055 24084 24064
rect 24032 24021 24041 24055
rect 24041 24021 24075 24055
rect 24075 24021 24084 24055
rect 24032 24012 24084 24021
rect 24768 24012 24820 24064
rect 24860 24055 24912 24064
rect 24860 24021 24869 24055
rect 24869 24021 24903 24055
rect 24903 24021 24912 24055
rect 24860 24012 24912 24021
rect 25780 24012 25832 24064
rect 27160 24123 27212 24132
rect 27160 24089 27169 24123
rect 27169 24089 27203 24123
rect 27203 24089 27212 24123
rect 27160 24080 27212 24089
rect 26240 24012 26292 24064
rect 27804 24055 27856 24064
rect 27804 24021 27813 24055
rect 27813 24021 27847 24055
rect 27847 24021 27856 24055
rect 27804 24012 27856 24021
rect 28816 24080 28868 24132
rect 29000 24123 29052 24132
rect 29000 24089 29009 24123
rect 29009 24089 29043 24123
rect 29043 24089 29052 24123
rect 29000 24080 29052 24089
rect 29276 24080 29328 24132
rect 32772 24157 32781 24191
rect 32781 24157 32815 24191
rect 32815 24157 32824 24191
rect 32772 24148 32824 24157
rect 30656 24123 30708 24132
rect 30656 24089 30690 24123
rect 30690 24089 30708 24123
rect 30656 24080 30708 24089
rect 33048 24123 33100 24132
rect 33048 24089 33057 24123
rect 33057 24089 33091 24123
rect 33091 24089 33100 24123
rect 33048 24080 33100 24089
rect 33508 24080 33560 24132
rect 28356 24012 28408 24064
rect 34520 24055 34572 24064
rect 34520 24021 34529 24055
rect 34529 24021 34563 24055
rect 34563 24021 34572 24055
rect 34520 24012 34572 24021
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 5448 23808 5500 23860
rect 6644 23808 6696 23860
rect 10140 23808 10192 23860
rect 3792 23672 3844 23724
rect 3884 23715 3936 23724
rect 3884 23681 3893 23715
rect 3893 23681 3927 23715
rect 3927 23681 3936 23715
rect 3884 23672 3936 23681
rect 5264 23672 5316 23724
rect 7196 23672 7248 23724
rect 8300 23715 8352 23724
rect 8300 23681 8309 23715
rect 8309 23681 8343 23715
rect 8343 23681 8352 23715
rect 8300 23672 8352 23681
rect 12716 23808 12768 23860
rect 13268 23851 13320 23860
rect 13268 23817 13277 23851
rect 13277 23817 13311 23851
rect 13311 23817 13320 23851
rect 13268 23808 13320 23817
rect 9036 23672 9088 23724
rect 9772 23672 9824 23724
rect 12440 23672 12492 23724
rect 13176 23672 13228 23724
rect 19156 23808 19208 23860
rect 19524 23808 19576 23860
rect 15752 23740 15804 23792
rect 12716 23604 12768 23656
rect 15936 23672 15988 23724
rect 19340 23740 19392 23792
rect 18052 23672 18104 23724
rect 18972 23715 19024 23724
rect 18972 23681 18981 23715
rect 18981 23681 19015 23715
rect 19015 23681 19024 23715
rect 18972 23672 19024 23681
rect 19064 23672 19116 23724
rect 21732 23740 21784 23792
rect 22008 23808 22060 23860
rect 22468 23808 22520 23860
rect 23848 23808 23900 23860
rect 24308 23808 24360 23860
rect 24676 23808 24728 23860
rect 26516 23808 26568 23860
rect 15844 23647 15896 23656
rect 15844 23613 15853 23647
rect 15853 23613 15887 23647
rect 15887 23613 15896 23647
rect 15844 23604 15896 23613
rect 22100 23672 22152 23724
rect 22284 23672 22336 23724
rect 22560 23715 22612 23724
rect 22560 23681 22569 23715
rect 22569 23681 22603 23715
rect 22603 23681 22612 23715
rect 22560 23672 22612 23681
rect 22836 23715 22888 23724
rect 22836 23681 22870 23715
rect 22870 23681 22888 23715
rect 22836 23672 22888 23681
rect 23204 23672 23256 23724
rect 21640 23604 21692 23656
rect 24768 23672 24820 23724
rect 26332 23672 26384 23724
rect 26608 23604 26660 23656
rect 7656 23536 7708 23588
rect 8208 23536 8260 23588
rect 11336 23579 11388 23588
rect 11336 23545 11345 23579
rect 11345 23545 11379 23579
rect 11379 23545 11388 23579
rect 11336 23536 11388 23545
rect 4620 23468 4672 23520
rect 5264 23511 5316 23520
rect 5264 23477 5273 23511
rect 5273 23477 5307 23511
rect 5307 23477 5316 23511
rect 5264 23468 5316 23477
rect 8024 23511 8076 23520
rect 8024 23477 8033 23511
rect 8033 23477 8067 23511
rect 8067 23477 8076 23511
rect 8024 23468 8076 23477
rect 10232 23468 10284 23520
rect 15752 23468 15804 23520
rect 18420 23468 18472 23520
rect 19248 23468 19300 23520
rect 21732 23468 21784 23520
rect 22468 23468 22520 23520
rect 26148 23468 26200 23520
rect 29644 23808 29696 23860
rect 29920 23808 29972 23860
rect 30656 23851 30708 23860
rect 30656 23817 30665 23851
rect 30665 23817 30699 23851
rect 30699 23817 30708 23851
rect 30656 23808 30708 23817
rect 30932 23808 30984 23860
rect 31760 23808 31812 23860
rect 33048 23808 33100 23860
rect 27988 23740 28040 23792
rect 27252 23715 27304 23724
rect 27252 23681 27286 23715
rect 27286 23681 27304 23715
rect 27252 23672 27304 23681
rect 34796 23783 34848 23792
rect 34796 23749 34805 23783
rect 34805 23749 34839 23783
rect 34839 23749 34848 23783
rect 34796 23740 34848 23749
rect 28908 23715 28960 23724
rect 28908 23681 28942 23715
rect 28942 23681 28960 23715
rect 28908 23672 28960 23681
rect 30656 23672 30708 23724
rect 31300 23672 31352 23724
rect 31392 23672 31444 23724
rect 34244 23672 34296 23724
rect 34520 23715 34572 23724
rect 34520 23681 34529 23715
rect 34529 23681 34563 23715
rect 34563 23681 34572 23715
rect 34520 23672 34572 23681
rect 27160 23468 27212 23520
rect 30932 23604 30984 23656
rect 29644 23468 29696 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 4160 23128 4212 23180
rect 6460 23196 6512 23248
rect 4620 22992 4672 23044
rect 6092 23060 6144 23112
rect 7196 23239 7248 23248
rect 7196 23205 7205 23239
rect 7205 23205 7239 23239
rect 7239 23205 7248 23239
rect 7196 23196 7248 23205
rect 8024 23196 8076 23248
rect 8116 23196 8168 23248
rect 7656 23171 7708 23180
rect 7656 23137 7665 23171
rect 7665 23137 7699 23171
rect 7699 23137 7708 23171
rect 7656 23128 7708 23137
rect 7748 23171 7800 23180
rect 7748 23137 7757 23171
rect 7757 23137 7791 23171
rect 7791 23137 7800 23171
rect 7748 23128 7800 23137
rect 7840 23060 7892 23112
rect 8852 23060 8904 23112
rect 10416 23264 10468 23316
rect 10876 23307 10928 23316
rect 10876 23273 10885 23307
rect 10885 23273 10919 23307
rect 10919 23273 10928 23307
rect 10876 23264 10928 23273
rect 11796 23307 11848 23316
rect 11796 23273 11805 23307
rect 11805 23273 11839 23307
rect 11839 23273 11848 23307
rect 11796 23264 11848 23273
rect 9772 23171 9824 23180
rect 9772 23137 9781 23171
rect 9781 23137 9815 23171
rect 9815 23137 9824 23171
rect 9772 23128 9824 23137
rect 10048 23060 10100 23112
rect 10232 23103 10284 23112
rect 10232 23069 10241 23103
rect 10241 23069 10275 23103
rect 10275 23069 10284 23103
rect 10232 23060 10284 23069
rect 8760 22992 8812 23044
rect 10692 23128 10744 23180
rect 10968 23128 11020 23180
rect 10876 23060 10928 23112
rect 11152 23060 11204 23112
rect 11336 23103 11388 23112
rect 11336 23069 11345 23103
rect 11345 23069 11379 23103
rect 11379 23069 11388 23103
rect 11336 23060 11388 23069
rect 12808 23264 12860 23316
rect 14096 23264 14148 23316
rect 16396 23196 16448 23248
rect 17040 23196 17092 23248
rect 16028 23128 16080 23180
rect 12164 23103 12216 23112
rect 12164 23069 12173 23103
rect 12173 23069 12207 23103
rect 12207 23069 12216 23103
rect 12164 23060 12216 23069
rect 14372 23060 14424 23112
rect 8944 22924 8996 22976
rect 9956 22967 10008 22976
rect 9956 22933 9965 22967
rect 9965 22933 9999 22967
rect 9999 22933 10008 22967
rect 9956 22924 10008 22933
rect 12716 22992 12768 23044
rect 14832 22992 14884 23044
rect 16212 23103 16264 23112
rect 16212 23069 16226 23103
rect 16226 23069 16260 23103
rect 16260 23069 16264 23103
rect 16212 23060 16264 23069
rect 13544 22967 13596 22976
rect 13544 22933 13553 22967
rect 13553 22933 13587 22967
rect 13587 22933 13596 22967
rect 13544 22924 13596 22933
rect 15660 22967 15712 22976
rect 15660 22933 15669 22967
rect 15669 22933 15703 22967
rect 15703 22933 15712 22967
rect 15660 22924 15712 22933
rect 16120 23035 16172 23044
rect 16120 23001 16129 23035
rect 16129 23001 16163 23035
rect 16163 23001 16172 23035
rect 16120 22992 16172 23001
rect 17040 22992 17092 23044
rect 22836 23264 22888 23316
rect 22744 23196 22796 23248
rect 23388 23196 23440 23248
rect 25780 23307 25832 23316
rect 25780 23273 25789 23307
rect 25789 23273 25823 23307
rect 25823 23273 25832 23307
rect 25780 23264 25832 23273
rect 26424 23307 26476 23316
rect 26424 23273 26433 23307
rect 26433 23273 26467 23307
rect 26467 23273 26476 23307
rect 26424 23264 26476 23273
rect 26516 23307 26568 23316
rect 26516 23273 26525 23307
rect 26525 23273 26559 23307
rect 26559 23273 26568 23307
rect 26516 23264 26568 23273
rect 27252 23264 27304 23316
rect 27712 23264 27764 23316
rect 28172 23264 28224 23316
rect 28908 23264 28960 23316
rect 18972 23171 19024 23180
rect 18972 23137 18981 23171
rect 18981 23137 19015 23171
rect 19015 23137 19024 23171
rect 18972 23128 19024 23137
rect 23572 23171 23624 23180
rect 23572 23137 23581 23171
rect 23581 23137 23615 23171
rect 23615 23137 23624 23171
rect 23572 23128 23624 23137
rect 21732 23103 21784 23112
rect 21732 23069 21766 23103
rect 21766 23069 21784 23103
rect 21732 23060 21784 23069
rect 24308 23060 24360 23112
rect 24952 23060 25004 23112
rect 18236 22992 18288 23044
rect 16764 22924 16816 22976
rect 22284 22924 22336 22976
rect 23480 22924 23532 22976
rect 23940 22924 23992 22976
rect 24860 22992 24912 23044
rect 27528 23196 27580 23248
rect 29460 23128 29512 23180
rect 30748 23128 30800 23180
rect 27160 23060 27212 23112
rect 29552 23060 29604 23112
rect 29920 23103 29972 23112
rect 29920 23069 29929 23103
rect 29929 23069 29963 23103
rect 29963 23069 29972 23103
rect 29920 23060 29972 23069
rect 26240 22924 26292 22976
rect 29276 22924 29328 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 3792 22763 3844 22772
rect 3792 22729 3801 22763
rect 3801 22729 3835 22763
rect 3835 22729 3844 22763
rect 3792 22720 3844 22729
rect 4528 22720 4580 22772
rect 4712 22720 4764 22772
rect 1308 22584 1360 22636
rect 7748 22720 7800 22772
rect 8760 22720 8812 22772
rect 8852 22763 8904 22772
rect 8852 22729 8861 22763
rect 8861 22729 8895 22763
rect 8895 22729 8904 22763
rect 8852 22720 8904 22729
rect 9036 22763 9088 22772
rect 9036 22729 9045 22763
rect 9045 22729 9079 22763
rect 9079 22729 9088 22763
rect 9036 22720 9088 22729
rect 10232 22720 10284 22772
rect 12716 22763 12768 22772
rect 12716 22729 12725 22763
rect 12725 22729 12759 22763
rect 12759 22729 12768 22763
rect 12716 22720 12768 22729
rect 14372 22720 14424 22772
rect 14832 22763 14884 22772
rect 14832 22729 14841 22763
rect 14841 22729 14875 22763
rect 14875 22729 14884 22763
rect 14832 22720 14884 22729
rect 15660 22720 15712 22772
rect 5264 22652 5316 22704
rect 9956 22652 10008 22704
rect 10508 22652 10560 22704
rect 5724 22584 5776 22636
rect 8116 22584 8168 22636
rect 8300 22584 8352 22636
rect 9772 22584 9824 22636
rect 10416 22584 10468 22636
rect 13544 22627 13596 22636
rect 13544 22593 13553 22627
rect 13553 22593 13587 22627
rect 13587 22593 13596 22627
rect 13544 22584 13596 22593
rect 13820 22627 13872 22636
rect 13820 22593 13829 22627
rect 13829 22593 13863 22627
rect 13863 22593 13872 22627
rect 13820 22584 13872 22593
rect 16028 22584 16080 22636
rect 16488 22627 16540 22636
rect 16488 22593 16497 22627
rect 16497 22593 16531 22627
rect 16531 22593 16540 22627
rect 16488 22584 16540 22593
rect 17776 22720 17828 22772
rect 18052 22720 18104 22772
rect 18328 22763 18380 22772
rect 18328 22729 18337 22763
rect 18337 22729 18371 22763
rect 18371 22729 18380 22763
rect 18328 22720 18380 22729
rect 18420 22763 18472 22772
rect 18420 22729 18429 22763
rect 18429 22729 18463 22763
rect 18463 22729 18472 22763
rect 18420 22720 18472 22729
rect 19340 22763 19392 22772
rect 19340 22729 19349 22763
rect 19349 22729 19383 22763
rect 19383 22729 19392 22763
rect 19340 22720 19392 22729
rect 19524 22720 19576 22772
rect 16764 22652 16816 22704
rect 17224 22627 17276 22636
rect 17224 22593 17233 22627
rect 17233 22593 17267 22627
rect 17267 22593 17276 22627
rect 17224 22584 17276 22593
rect 21916 22720 21968 22772
rect 25964 22720 26016 22772
rect 26608 22720 26660 22772
rect 27252 22720 27304 22772
rect 1860 22491 1912 22500
rect 1860 22457 1869 22491
rect 1869 22457 1903 22491
rect 1903 22457 1912 22491
rect 1860 22448 1912 22457
rect 4712 22516 4764 22568
rect 5448 22516 5500 22568
rect 5540 22516 5592 22568
rect 9680 22516 9732 22568
rect 13176 22559 13228 22568
rect 13176 22525 13185 22559
rect 13185 22525 13219 22559
rect 13219 22525 13228 22559
rect 13176 22516 13228 22525
rect 13268 22559 13320 22568
rect 13268 22525 13277 22559
rect 13277 22525 13311 22559
rect 13311 22525 13320 22559
rect 13268 22516 13320 22525
rect 13452 22516 13504 22568
rect 15752 22516 15804 22568
rect 16212 22559 16264 22568
rect 16212 22525 16221 22559
rect 16221 22525 16255 22559
rect 16255 22525 16264 22559
rect 16212 22516 16264 22525
rect 16764 22516 16816 22568
rect 4804 22380 4856 22432
rect 5264 22380 5316 22432
rect 5724 22423 5776 22432
rect 5724 22389 5733 22423
rect 5733 22389 5767 22423
rect 5767 22389 5776 22423
rect 5724 22380 5776 22389
rect 17868 22516 17920 22568
rect 20444 22516 20496 22568
rect 23756 22584 23808 22636
rect 24952 22627 25004 22636
rect 24952 22593 24961 22627
rect 24961 22593 24995 22627
rect 24995 22593 25004 22627
rect 24952 22584 25004 22593
rect 25504 22584 25556 22636
rect 26332 22584 26384 22636
rect 27160 22584 27212 22636
rect 22192 22559 22244 22568
rect 22192 22525 22201 22559
rect 22201 22525 22235 22559
rect 22235 22525 22244 22559
rect 22192 22516 22244 22525
rect 22836 22516 22888 22568
rect 29276 22720 29328 22772
rect 29184 22652 29236 22704
rect 28172 22584 28224 22636
rect 29552 22584 29604 22636
rect 30104 22584 30156 22636
rect 30564 22627 30616 22636
rect 30564 22593 30582 22627
rect 30582 22593 30616 22627
rect 30564 22584 30616 22593
rect 31392 22627 31444 22636
rect 31392 22593 31401 22627
rect 31401 22593 31435 22627
rect 31435 22593 31444 22627
rect 31392 22584 31444 22593
rect 34244 22584 34296 22636
rect 34520 22627 34572 22636
rect 34520 22593 34529 22627
rect 34529 22593 34563 22627
rect 34563 22593 34572 22627
rect 34520 22584 34572 22593
rect 29736 22516 29788 22568
rect 34796 22559 34848 22568
rect 34796 22525 34805 22559
rect 34805 22525 34839 22559
rect 34839 22525 34848 22559
rect 34796 22516 34848 22525
rect 8944 22380 8996 22432
rect 11244 22423 11296 22432
rect 11244 22389 11253 22423
rect 11253 22389 11287 22423
rect 11287 22389 11296 22423
rect 11244 22380 11296 22389
rect 12256 22380 12308 22432
rect 23572 22448 23624 22500
rect 29092 22448 29144 22500
rect 17408 22423 17460 22432
rect 17408 22389 17417 22423
rect 17417 22389 17451 22423
rect 17451 22389 17460 22423
rect 17408 22380 17460 22389
rect 19248 22380 19300 22432
rect 20812 22380 20864 22432
rect 22744 22380 22796 22432
rect 29276 22423 29328 22432
rect 29276 22389 29285 22423
rect 29285 22389 29319 22423
rect 29319 22389 29328 22423
rect 29276 22380 29328 22389
rect 29460 22423 29512 22432
rect 29460 22389 29469 22423
rect 29469 22389 29503 22423
rect 29503 22389 29512 22423
rect 29460 22380 29512 22389
rect 29736 22380 29788 22432
rect 33048 22380 33100 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 5356 22176 5408 22228
rect 5632 22176 5684 22228
rect 6184 22176 6236 22228
rect 12072 22176 12124 22228
rect 5172 22108 5224 22160
rect 8944 22108 8996 22160
rect 12900 22176 12952 22228
rect 13268 22176 13320 22228
rect 4528 22040 4580 22092
rect 4712 21972 4764 22024
rect 9864 22040 9916 22092
rect 15476 22108 15528 22160
rect 15752 22108 15804 22160
rect 8484 21972 8536 22024
rect 11244 21972 11296 22024
rect 12164 22015 12216 22024
rect 12164 21981 12173 22015
rect 12173 21981 12207 22015
rect 12207 21981 12216 22015
rect 12164 21972 12216 21981
rect 16856 22176 16908 22228
rect 17408 22176 17460 22228
rect 17224 22108 17276 22160
rect 18972 22108 19024 22160
rect 15936 21972 15988 22024
rect 20444 22040 20496 22092
rect 3148 21836 3200 21888
rect 4160 21879 4212 21888
rect 4160 21845 4169 21879
rect 4169 21845 4203 21879
rect 4203 21845 4212 21879
rect 4160 21836 4212 21845
rect 4528 21836 4580 21888
rect 4712 21836 4764 21888
rect 5540 21904 5592 21956
rect 9680 21904 9732 21956
rect 10416 21879 10468 21888
rect 10416 21845 10425 21879
rect 10425 21845 10459 21879
rect 10459 21845 10468 21879
rect 10416 21836 10468 21845
rect 12808 21904 12860 21956
rect 13176 21904 13228 21956
rect 13820 21836 13872 21888
rect 14832 21879 14884 21888
rect 14832 21845 14841 21879
rect 14841 21845 14875 21879
rect 14875 21845 14884 21879
rect 14832 21836 14884 21845
rect 15200 21879 15252 21888
rect 15200 21845 15209 21879
rect 15209 21845 15243 21879
rect 15243 21845 15252 21879
rect 15200 21836 15252 21845
rect 15844 21879 15896 21888
rect 15844 21845 15853 21879
rect 15853 21845 15887 21879
rect 15887 21845 15896 21879
rect 15844 21836 15896 21845
rect 16672 21904 16724 21956
rect 19248 22015 19300 22024
rect 19248 21981 19257 22015
rect 19257 21981 19291 22015
rect 19291 21981 19300 22015
rect 19248 21972 19300 21981
rect 20076 21972 20128 22024
rect 20260 21904 20312 21956
rect 17040 21836 17092 21888
rect 18696 21836 18748 21888
rect 18788 21879 18840 21888
rect 18788 21845 18797 21879
rect 18797 21845 18831 21879
rect 18831 21845 18840 21879
rect 20720 21972 20772 22024
rect 23664 22108 23716 22160
rect 25504 22219 25556 22228
rect 25504 22185 25513 22219
rect 25513 22185 25547 22219
rect 25547 22185 25556 22219
rect 25504 22176 25556 22185
rect 26516 22176 26568 22228
rect 29092 22176 29144 22228
rect 22836 22083 22888 22092
rect 22836 22049 22845 22083
rect 22845 22049 22879 22083
rect 22879 22049 22888 22083
rect 22836 22040 22888 22049
rect 24032 22040 24084 22092
rect 25780 22040 25832 22092
rect 25964 22083 26016 22092
rect 25964 22049 25973 22083
rect 25973 22049 26007 22083
rect 26007 22049 26016 22083
rect 25964 22040 26016 22049
rect 26148 22083 26200 22092
rect 26148 22049 26157 22083
rect 26157 22049 26191 22083
rect 26191 22049 26200 22083
rect 26148 22040 26200 22049
rect 22468 21972 22520 22024
rect 24308 21972 24360 22024
rect 26608 21972 26660 22024
rect 27068 22015 27120 22024
rect 27068 21981 27077 22015
rect 27077 21981 27111 22015
rect 27111 21981 27120 22015
rect 27068 21972 27120 21981
rect 30564 22219 30616 22228
rect 30564 22185 30573 22219
rect 30573 22185 30607 22219
rect 30607 22185 30616 22219
rect 30564 22176 30616 22185
rect 33048 22219 33100 22228
rect 33048 22185 33078 22219
rect 33078 22185 33100 22219
rect 33048 22176 33100 22185
rect 34520 22219 34572 22228
rect 34520 22185 34529 22219
rect 34529 22185 34563 22219
rect 34563 22185 34572 22219
rect 34520 22176 34572 22185
rect 29368 22108 29420 22160
rect 28540 22015 28592 22024
rect 28540 21981 28549 22015
rect 28549 21981 28583 22015
rect 28583 21981 28592 22015
rect 28540 21972 28592 21981
rect 28632 21972 28684 22024
rect 29460 22040 29512 22092
rect 18788 21836 18840 21845
rect 21180 21836 21232 21888
rect 22744 21947 22796 21956
rect 22744 21913 22753 21947
rect 22753 21913 22787 21947
rect 22787 21913 22796 21947
rect 22744 21904 22796 21913
rect 23020 21836 23072 21888
rect 23388 21836 23440 21888
rect 23664 21836 23716 21888
rect 24032 21879 24084 21888
rect 24032 21845 24041 21879
rect 24041 21845 24075 21879
rect 24075 21845 24084 21879
rect 24032 21836 24084 21845
rect 24860 21904 24912 21956
rect 24952 21904 25004 21956
rect 25228 21947 25280 21956
rect 25228 21913 25237 21947
rect 25237 21913 25271 21947
rect 25271 21913 25280 21947
rect 25228 21904 25280 21913
rect 25320 21904 25372 21956
rect 29276 21972 29328 22024
rect 29368 22015 29420 22024
rect 29368 21981 29377 22015
rect 29377 21981 29411 22015
rect 29411 21981 29420 22015
rect 29368 21972 29420 21981
rect 29552 22015 29604 22024
rect 29552 21981 29561 22015
rect 29561 21981 29595 22015
rect 29595 21981 29604 22015
rect 29552 21972 29604 21981
rect 30380 21972 30432 22024
rect 31024 22040 31076 22092
rect 27620 21904 27672 21956
rect 29644 21904 29696 21956
rect 31392 21972 31444 22024
rect 33140 22040 33192 22092
rect 33508 21904 33560 21956
rect 28816 21836 28868 21888
rect 28908 21836 28960 21888
rect 29000 21836 29052 21888
rect 29460 21836 29512 21888
rect 31024 21879 31076 21888
rect 31024 21845 31033 21879
rect 31033 21845 31067 21879
rect 31067 21845 31076 21879
rect 31024 21836 31076 21845
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 4160 21632 4212 21684
rect 4712 21675 4764 21684
rect 4712 21641 4721 21675
rect 4721 21641 4755 21675
rect 4755 21641 4764 21675
rect 4712 21632 4764 21641
rect 3148 21564 3200 21616
rect 4620 21564 4672 21616
rect 5356 21564 5408 21616
rect 6460 21564 6512 21616
rect 8300 21632 8352 21684
rect 9864 21675 9916 21684
rect 9864 21641 9873 21675
rect 9873 21641 9907 21675
rect 9907 21641 9916 21675
rect 9864 21632 9916 21641
rect 4068 21496 4120 21548
rect 5816 21496 5868 21548
rect 8116 21564 8168 21616
rect 9772 21564 9824 21616
rect 4804 21471 4856 21480
rect 4804 21437 4813 21471
rect 4813 21437 4847 21471
rect 4847 21437 4856 21471
rect 4804 21428 4856 21437
rect 4436 21292 4488 21344
rect 4712 21292 4764 21344
rect 6184 21335 6236 21344
rect 6184 21301 6193 21335
rect 6193 21301 6227 21335
rect 6227 21301 6236 21335
rect 6184 21292 6236 21301
rect 7472 21292 7524 21344
rect 8024 21428 8076 21480
rect 8852 21428 8904 21480
rect 10968 21632 11020 21684
rect 12808 21675 12860 21684
rect 12808 21641 12817 21675
rect 12817 21641 12851 21675
rect 12851 21641 12860 21675
rect 12808 21632 12860 21641
rect 13176 21675 13228 21684
rect 13176 21641 13185 21675
rect 13185 21641 13219 21675
rect 13219 21641 13228 21675
rect 13176 21632 13228 21641
rect 15200 21632 15252 21684
rect 16120 21632 16172 21684
rect 16672 21675 16724 21684
rect 16672 21641 16681 21675
rect 16681 21641 16715 21675
rect 16715 21641 16724 21675
rect 16672 21632 16724 21641
rect 17040 21675 17092 21684
rect 17040 21641 17049 21675
rect 17049 21641 17083 21675
rect 17083 21641 17092 21675
rect 17040 21632 17092 21641
rect 17224 21632 17276 21684
rect 18604 21632 18656 21684
rect 13820 21564 13872 21616
rect 14832 21564 14884 21616
rect 15752 21607 15804 21616
rect 15752 21573 15761 21607
rect 15761 21573 15795 21607
rect 15795 21573 15804 21607
rect 15752 21564 15804 21573
rect 17500 21564 17552 21616
rect 13360 21471 13412 21480
rect 13360 21437 13369 21471
rect 13369 21437 13403 21471
rect 13403 21437 13412 21471
rect 13360 21428 13412 21437
rect 9588 21292 9640 21344
rect 10416 21335 10468 21344
rect 10416 21301 10425 21335
rect 10425 21301 10459 21335
rect 10459 21301 10468 21335
rect 10416 21292 10468 21301
rect 14556 21292 14608 21344
rect 18144 21496 18196 21548
rect 18972 21496 19024 21548
rect 19616 21496 19668 21548
rect 21180 21675 21232 21684
rect 21180 21641 21189 21675
rect 21189 21641 21223 21675
rect 21223 21641 21232 21675
rect 21180 21632 21232 21641
rect 22100 21675 22152 21684
rect 22100 21641 22109 21675
rect 22109 21641 22143 21675
rect 22143 21641 22152 21675
rect 22100 21632 22152 21641
rect 22928 21632 22980 21684
rect 24216 21632 24268 21684
rect 22008 21564 22060 21616
rect 24860 21632 24912 21684
rect 26056 21675 26108 21684
rect 26056 21641 26065 21675
rect 26065 21641 26099 21675
rect 26099 21641 26108 21675
rect 26056 21632 26108 21641
rect 27528 21675 27580 21684
rect 27528 21641 27537 21675
rect 27537 21641 27571 21675
rect 27571 21641 27580 21675
rect 27528 21632 27580 21641
rect 27620 21675 27672 21684
rect 27620 21641 27629 21675
rect 27629 21641 27663 21675
rect 27663 21641 27672 21675
rect 27620 21632 27672 21641
rect 28540 21632 28592 21684
rect 28816 21632 28868 21684
rect 17316 21471 17368 21480
rect 17316 21437 17325 21471
rect 17325 21437 17359 21471
rect 17359 21437 17368 21471
rect 17316 21428 17368 21437
rect 20720 21428 20772 21480
rect 20904 21539 20956 21548
rect 20904 21505 20913 21539
rect 20913 21505 20947 21539
rect 20947 21505 20956 21539
rect 20904 21496 20956 21505
rect 22284 21539 22336 21548
rect 22284 21505 22293 21539
rect 22293 21505 22327 21539
rect 22327 21505 22336 21539
rect 22284 21496 22336 21505
rect 22468 21539 22520 21548
rect 22468 21505 22478 21539
rect 22478 21505 22512 21539
rect 22512 21505 22520 21539
rect 22468 21496 22520 21505
rect 22744 21539 22796 21548
rect 22744 21505 22753 21539
rect 22753 21505 22787 21539
rect 22787 21505 22796 21539
rect 22744 21496 22796 21505
rect 23020 21496 23072 21548
rect 24032 21496 24084 21548
rect 27436 21564 27488 21616
rect 29552 21632 29604 21684
rect 29736 21675 29788 21684
rect 29736 21641 29745 21675
rect 29745 21641 29779 21675
rect 29779 21641 29788 21675
rect 29736 21632 29788 21641
rect 29920 21675 29972 21684
rect 29920 21641 29929 21675
rect 29929 21641 29963 21675
rect 29963 21641 29972 21675
rect 29920 21632 29972 21641
rect 29368 21564 29420 21616
rect 18512 21292 18564 21344
rect 20444 21335 20496 21344
rect 20444 21301 20453 21335
rect 20453 21301 20487 21335
rect 20487 21301 20496 21335
rect 20444 21292 20496 21301
rect 20904 21292 20956 21344
rect 22008 21292 22060 21344
rect 22100 21292 22152 21344
rect 24308 21360 24360 21412
rect 25504 21428 25556 21480
rect 26056 21428 26108 21480
rect 27896 21428 27948 21480
rect 28172 21471 28224 21480
rect 28172 21437 28181 21471
rect 28181 21437 28215 21471
rect 28215 21437 28224 21471
rect 28172 21428 28224 21437
rect 28816 21539 28868 21548
rect 28816 21505 28825 21539
rect 28825 21505 28859 21539
rect 28859 21505 28868 21539
rect 28816 21496 28868 21505
rect 28908 21539 28960 21548
rect 28908 21505 28953 21539
rect 28953 21505 28960 21539
rect 28908 21496 28960 21505
rect 29460 21496 29512 21548
rect 26884 21360 26936 21412
rect 27528 21360 27580 21412
rect 28724 21428 28776 21480
rect 29828 21360 29880 21412
rect 30288 21360 30340 21412
rect 30932 21403 30984 21412
rect 23480 21292 23532 21344
rect 25780 21335 25832 21344
rect 25780 21301 25789 21335
rect 25789 21301 25823 21335
rect 25823 21301 25832 21335
rect 25780 21292 25832 21301
rect 28356 21292 28408 21344
rect 30932 21369 30941 21403
rect 30941 21369 30975 21403
rect 30975 21369 30984 21403
rect 30932 21360 30984 21369
rect 31208 21360 31260 21412
rect 30748 21335 30800 21344
rect 30748 21301 30757 21335
rect 30757 21301 30791 21335
rect 30791 21301 30800 21335
rect 30748 21292 30800 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 4068 21088 4120 21140
rect 5816 21131 5868 21140
rect 5816 21097 5825 21131
rect 5825 21097 5859 21131
rect 5859 21097 5868 21131
rect 5816 21088 5868 21097
rect 7196 21088 7248 21140
rect 7840 21088 7892 21140
rect 8024 21088 8076 21140
rect 8392 21088 8444 21140
rect 6460 21020 6512 21072
rect 14096 21088 14148 21140
rect 15752 21088 15804 21140
rect 18144 21131 18196 21140
rect 18144 21097 18153 21131
rect 18153 21097 18187 21131
rect 18187 21097 18196 21131
rect 18144 21088 18196 21097
rect 19616 21131 19668 21140
rect 19616 21097 19625 21131
rect 19625 21097 19659 21131
rect 19659 21097 19668 21131
rect 19616 21088 19668 21097
rect 6368 20995 6420 21004
rect 6368 20961 6377 20995
rect 6377 20961 6411 20995
rect 6411 20961 6420 20995
rect 6368 20952 6420 20961
rect 4896 20884 4948 20936
rect 6184 20927 6236 20936
rect 6184 20893 6193 20927
rect 6193 20893 6227 20927
rect 6227 20893 6236 20927
rect 6184 20884 6236 20893
rect 7472 20927 7524 20936
rect 7472 20893 7481 20927
rect 7481 20893 7515 20927
rect 7515 20893 7524 20927
rect 7472 20884 7524 20893
rect 8392 20884 8444 20936
rect 9772 20995 9824 21004
rect 9772 20961 9781 20995
rect 9781 20961 9815 20995
rect 9815 20961 9824 20995
rect 9772 20952 9824 20961
rect 18604 20995 18656 21004
rect 18604 20961 18613 20995
rect 18613 20961 18647 20995
rect 18647 20961 18656 20995
rect 18604 20952 18656 20961
rect 18788 21020 18840 21072
rect 20812 21088 20864 21140
rect 25872 21088 25924 21140
rect 20076 21020 20128 21072
rect 22008 21020 22060 21072
rect 23848 21020 23900 21072
rect 24124 21020 24176 21072
rect 27436 21131 27488 21140
rect 27436 21097 27445 21131
rect 27445 21097 27479 21131
rect 27479 21097 27488 21131
rect 27436 21088 27488 21097
rect 29368 21088 29420 21140
rect 30012 21088 30064 21140
rect 30288 21088 30340 21140
rect 31208 21131 31260 21140
rect 31208 21097 31217 21131
rect 31217 21097 31251 21131
rect 31251 21097 31260 21131
rect 31208 21088 31260 21097
rect 29460 21020 29512 21072
rect 9864 20884 9916 20936
rect 12164 20884 12216 20936
rect 12348 20884 12400 20936
rect 14096 20884 14148 20936
rect 17684 20884 17736 20936
rect 19340 20952 19392 21004
rect 23480 20952 23532 21004
rect 20444 20884 20496 20936
rect 23848 20927 23900 20936
rect 23848 20893 23857 20927
rect 23857 20893 23891 20927
rect 23891 20893 23900 20927
rect 23848 20884 23900 20893
rect 4620 20859 4672 20868
rect 4620 20825 4629 20859
rect 4629 20825 4663 20859
rect 4663 20825 4672 20859
rect 4620 20816 4672 20825
rect 7656 20816 7708 20868
rect 8024 20816 8076 20868
rect 10324 20816 10376 20868
rect 12440 20816 12492 20868
rect 14556 20859 14608 20868
rect 14556 20825 14565 20859
rect 14565 20825 14599 20859
rect 14599 20825 14608 20859
rect 14556 20816 14608 20825
rect 17316 20816 17368 20868
rect 20536 20816 20588 20868
rect 20628 20816 20680 20868
rect 6368 20748 6420 20800
rect 8944 20791 8996 20800
rect 8944 20757 8953 20791
rect 8953 20757 8987 20791
rect 8987 20757 8996 20791
rect 8944 20748 8996 20757
rect 9312 20791 9364 20800
rect 9312 20757 9321 20791
rect 9321 20757 9355 20791
rect 9355 20757 9364 20791
rect 9312 20748 9364 20757
rect 9404 20791 9456 20800
rect 9404 20757 9413 20791
rect 9413 20757 9447 20791
rect 9447 20757 9456 20791
rect 9404 20748 9456 20757
rect 11152 20791 11204 20800
rect 11152 20757 11161 20791
rect 11161 20757 11195 20791
rect 11195 20757 11204 20791
rect 11152 20748 11204 20757
rect 13452 20748 13504 20800
rect 18696 20748 18748 20800
rect 19340 20748 19392 20800
rect 20076 20791 20128 20800
rect 20076 20757 20085 20791
rect 20085 20757 20119 20791
rect 20119 20757 20128 20791
rect 20076 20748 20128 20757
rect 22744 20748 22796 20800
rect 22928 20859 22980 20868
rect 22928 20825 22946 20859
rect 22946 20825 22980 20859
rect 22928 20816 22980 20825
rect 24308 20884 24360 20936
rect 27068 20952 27120 21004
rect 29644 20995 29696 21004
rect 25228 20884 25280 20936
rect 29644 20961 29653 20995
rect 29653 20961 29687 20995
rect 29687 20961 29696 20995
rect 29644 20952 29696 20961
rect 29460 20884 29512 20936
rect 29736 20884 29788 20936
rect 29920 20927 29972 20936
rect 29920 20893 29954 20927
rect 29954 20893 29972 20927
rect 29920 20884 29972 20893
rect 23664 20791 23716 20800
rect 23664 20757 23673 20791
rect 23673 20757 23707 20791
rect 23707 20757 23716 20791
rect 23664 20748 23716 20757
rect 24308 20748 24360 20800
rect 24952 20816 25004 20868
rect 25044 20816 25096 20868
rect 25688 20816 25740 20868
rect 26976 20816 27028 20868
rect 27804 20859 27856 20868
rect 27804 20825 27838 20859
rect 27838 20825 27856 20859
rect 27804 20816 27856 20825
rect 31116 20816 31168 20868
rect 34704 20884 34756 20936
rect 31576 20816 31628 20868
rect 35348 20816 35400 20868
rect 25320 20748 25372 20800
rect 26056 20748 26108 20800
rect 27528 20748 27580 20800
rect 28264 20748 28316 20800
rect 28908 20791 28960 20800
rect 28908 20757 28917 20791
rect 28917 20757 28951 20791
rect 28951 20757 28960 20791
rect 28908 20748 28960 20757
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 9312 20544 9364 20596
rect 8944 20476 8996 20528
rect 1308 20408 1360 20460
rect 8116 20451 8168 20460
rect 8116 20417 8125 20451
rect 8125 20417 8159 20451
rect 8159 20417 8168 20451
rect 8116 20408 8168 20417
rect 10324 20587 10376 20596
rect 10324 20553 10333 20587
rect 10333 20553 10367 20587
rect 10367 20553 10376 20587
rect 10324 20544 10376 20553
rect 11152 20544 11204 20596
rect 11612 20544 11664 20596
rect 15568 20544 15620 20596
rect 19984 20587 20036 20596
rect 19984 20553 19993 20587
rect 19993 20553 20027 20587
rect 20027 20553 20036 20587
rect 19984 20544 20036 20553
rect 22744 20544 22796 20596
rect 22928 20544 22980 20596
rect 24400 20544 24452 20596
rect 25320 20587 25372 20596
rect 25320 20553 25329 20587
rect 25329 20553 25363 20587
rect 25363 20553 25372 20587
rect 25320 20544 25372 20553
rect 26056 20544 26108 20596
rect 26424 20587 26476 20596
rect 26424 20553 26433 20587
rect 26433 20553 26467 20587
rect 26467 20553 26476 20587
rect 26424 20544 26476 20553
rect 26976 20587 27028 20596
rect 26976 20553 26985 20587
rect 26985 20553 27019 20587
rect 27019 20553 27028 20587
rect 26976 20544 27028 20553
rect 27436 20544 27488 20596
rect 27804 20587 27856 20596
rect 27804 20553 27813 20587
rect 27813 20553 27847 20587
rect 27847 20553 27856 20587
rect 27804 20544 27856 20553
rect 28908 20544 28960 20596
rect 29368 20587 29420 20596
rect 29368 20553 29377 20587
rect 29377 20553 29411 20587
rect 29411 20553 29420 20587
rect 29368 20544 29420 20553
rect 12348 20476 12400 20528
rect 10324 20408 10376 20460
rect 3792 20204 3844 20256
rect 5540 20204 5592 20256
rect 10416 20340 10468 20392
rect 10232 20247 10284 20256
rect 10232 20213 10241 20247
rect 10241 20213 10275 20247
rect 10275 20213 10284 20247
rect 10232 20204 10284 20213
rect 12348 20383 12400 20392
rect 12348 20349 12357 20383
rect 12357 20349 12391 20383
rect 12391 20349 12400 20383
rect 12348 20340 12400 20349
rect 13452 20408 13504 20460
rect 14556 20476 14608 20528
rect 14096 20408 14148 20460
rect 17040 20451 17092 20460
rect 17040 20417 17049 20451
rect 17049 20417 17083 20451
rect 17083 20417 17092 20451
rect 17040 20408 17092 20417
rect 22100 20476 22152 20528
rect 23756 20476 23808 20528
rect 27896 20476 27948 20528
rect 28724 20476 28776 20528
rect 22652 20408 22704 20460
rect 24032 20451 24084 20460
rect 24032 20417 24041 20451
rect 24041 20417 24075 20451
rect 24075 20417 24084 20451
rect 24032 20408 24084 20417
rect 24216 20408 24268 20460
rect 26608 20408 26660 20460
rect 32220 20476 32272 20528
rect 33508 20476 33560 20528
rect 12900 20383 12952 20392
rect 12900 20349 12909 20383
rect 12909 20349 12943 20383
rect 12943 20349 12952 20383
rect 12900 20340 12952 20349
rect 12992 20340 13044 20392
rect 15936 20340 15988 20392
rect 17224 20383 17276 20392
rect 17224 20349 17233 20383
rect 17233 20349 17267 20383
rect 17267 20349 17276 20383
rect 17224 20340 17276 20349
rect 22468 20383 22520 20392
rect 22468 20349 22477 20383
rect 22477 20349 22511 20383
rect 22511 20349 22520 20383
rect 22468 20340 22520 20349
rect 24124 20383 24176 20392
rect 24124 20349 24133 20383
rect 24133 20349 24167 20383
rect 24167 20349 24176 20383
rect 24124 20340 24176 20349
rect 24952 20340 25004 20392
rect 26056 20340 26108 20392
rect 26424 20340 26476 20392
rect 29828 20451 29880 20460
rect 29828 20417 29837 20451
rect 29837 20417 29871 20451
rect 29871 20417 29880 20451
rect 29828 20408 29880 20417
rect 30288 20408 30340 20460
rect 28356 20383 28408 20392
rect 28356 20349 28365 20383
rect 28365 20349 28399 20383
rect 28399 20349 28408 20383
rect 28356 20340 28408 20349
rect 12440 20315 12492 20324
rect 12440 20281 12449 20315
rect 12449 20281 12483 20315
rect 12483 20281 12492 20315
rect 12440 20272 12492 20281
rect 15844 20272 15896 20324
rect 19432 20272 19484 20324
rect 14648 20204 14700 20256
rect 16672 20247 16724 20256
rect 16672 20213 16681 20247
rect 16681 20213 16715 20247
rect 16715 20213 16724 20247
rect 16672 20204 16724 20213
rect 23572 20204 23624 20256
rect 23664 20204 23716 20256
rect 24308 20204 24360 20256
rect 24860 20204 24912 20256
rect 26608 20315 26660 20324
rect 26608 20281 26617 20315
rect 26617 20281 26651 20315
rect 26651 20281 26660 20315
rect 26608 20272 26660 20281
rect 26792 20272 26844 20324
rect 27804 20204 27856 20256
rect 30380 20247 30432 20256
rect 30380 20213 30389 20247
rect 30389 20213 30423 20247
rect 30423 20213 30432 20247
rect 30380 20204 30432 20213
rect 33140 20408 33192 20460
rect 33968 20340 34020 20392
rect 31392 20204 31444 20256
rect 34704 20204 34756 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 9680 20000 9732 20052
rect 4160 19932 4212 19984
rect 8484 19932 8536 19984
rect 4804 19907 4856 19916
rect 4804 19873 4813 19907
rect 4813 19873 4847 19907
rect 4847 19873 4856 19907
rect 4804 19864 4856 19873
rect 10416 19864 10468 19916
rect 12532 19932 12584 19984
rect 12900 19932 12952 19984
rect 16764 20000 16816 20052
rect 17040 20000 17092 20052
rect 24032 20000 24084 20052
rect 24860 20043 24912 20052
rect 24860 20009 24869 20043
rect 24869 20009 24903 20043
rect 24903 20009 24912 20043
rect 24860 20000 24912 20009
rect 32036 20000 32088 20052
rect 33416 20000 33468 20052
rect 33968 20043 34020 20052
rect 33968 20009 33977 20043
rect 33977 20009 34011 20043
rect 34011 20009 34020 20043
rect 33968 20000 34020 20009
rect 13912 19864 13964 19916
rect 22100 19975 22152 19984
rect 22100 19941 22109 19975
rect 22109 19941 22143 19975
rect 22143 19941 22152 19975
rect 22100 19932 22152 19941
rect 23572 19932 23624 19984
rect 25596 19932 25648 19984
rect 3792 19839 3844 19848
rect 3792 19805 3801 19839
rect 3801 19805 3835 19839
rect 3835 19805 3844 19839
rect 3792 19796 3844 19805
rect 4436 19796 4488 19848
rect 5448 19796 5500 19848
rect 15016 19907 15068 19916
rect 15016 19873 15025 19907
rect 15025 19873 15059 19907
rect 15059 19873 15068 19907
rect 15016 19864 15068 19873
rect 14556 19796 14608 19848
rect 14924 19796 14976 19848
rect 16580 19796 16632 19848
rect 5356 19728 5408 19780
rect 6000 19728 6052 19780
rect 10416 19771 10468 19780
rect 10416 19737 10425 19771
rect 10425 19737 10459 19771
rect 10459 19737 10468 19771
rect 10416 19728 10468 19737
rect 12808 19728 12860 19780
rect 6184 19703 6236 19712
rect 6184 19669 6193 19703
rect 6193 19669 6227 19703
rect 6227 19669 6236 19703
rect 6184 19660 6236 19669
rect 6644 19660 6696 19712
rect 11612 19660 11664 19712
rect 12716 19660 12768 19712
rect 14096 19703 14148 19712
rect 14096 19669 14105 19703
rect 14105 19669 14139 19703
rect 14139 19669 14148 19703
rect 14096 19660 14148 19669
rect 14648 19660 14700 19712
rect 14832 19660 14884 19712
rect 15108 19660 15160 19712
rect 16672 19728 16724 19780
rect 18236 19728 18288 19780
rect 17224 19660 17276 19712
rect 18604 19660 18656 19712
rect 19432 19839 19484 19848
rect 19432 19805 19441 19839
rect 19441 19805 19475 19839
rect 19475 19805 19484 19839
rect 19432 19796 19484 19805
rect 19524 19771 19576 19780
rect 19524 19737 19533 19771
rect 19533 19737 19567 19771
rect 19567 19737 19576 19771
rect 19524 19728 19576 19737
rect 20628 19796 20680 19848
rect 19984 19728 20036 19780
rect 20536 19728 20588 19780
rect 21456 19839 21508 19848
rect 21456 19805 21465 19839
rect 21465 19805 21499 19839
rect 21499 19805 21508 19839
rect 21456 19796 21508 19805
rect 21732 19839 21784 19848
rect 21732 19805 21741 19839
rect 21741 19805 21775 19839
rect 21775 19805 21784 19839
rect 21732 19796 21784 19805
rect 22100 19796 22152 19848
rect 22652 19864 22704 19916
rect 23204 19864 23256 19916
rect 23296 19864 23348 19916
rect 26700 19864 26752 19916
rect 30380 19864 30432 19916
rect 23848 19771 23900 19780
rect 23848 19737 23857 19771
rect 23857 19737 23891 19771
rect 23891 19737 23900 19771
rect 23848 19728 23900 19737
rect 26148 19796 26200 19848
rect 32496 19796 32548 19848
rect 34244 19796 34296 19848
rect 25964 19728 26016 19780
rect 32036 19771 32088 19780
rect 32036 19737 32045 19771
rect 32045 19737 32079 19771
rect 32079 19737 32088 19771
rect 32036 19728 32088 19737
rect 32220 19771 32272 19780
rect 32220 19737 32229 19771
rect 32229 19737 32263 19771
rect 32263 19737 32272 19771
rect 32220 19728 32272 19737
rect 34704 19728 34756 19780
rect 34888 19771 34940 19780
rect 34888 19737 34897 19771
rect 34897 19737 34931 19771
rect 34931 19737 34940 19771
rect 34888 19728 34940 19737
rect 21272 19703 21324 19712
rect 21272 19669 21281 19703
rect 21281 19669 21315 19703
rect 21315 19669 21324 19703
rect 21272 19660 21324 19669
rect 22376 19703 22428 19712
rect 22376 19669 22385 19703
rect 22385 19669 22419 19703
rect 22419 19669 22428 19703
rect 22376 19660 22428 19669
rect 22744 19703 22796 19712
rect 22744 19669 22753 19703
rect 22753 19669 22787 19703
rect 22787 19669 22796 19703
rect 22744 19660 22796 19669
rect 23204 19703 23256 19712
rect 23204 19669 23213 19703
rect 23213 19669 23247 19703
rect 23247 19669 23256 19703
rect 23204 19660 23256 19669
rect 23664 19660 23716 19712
rect 24032 19703 24084 19712
rect 24032 19669 24041 19703
rect 24041 19669 24075 19703
rect 24075 19669 24084 19703
rect 24032 19660 24084 19669
rect 26700 19660 26752 19712
rect 26976 19660 27028 19712
rect 28356 19660 28408 19712
rect 30472 19660 30524 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 3516 19388 3568 19440
rect 4160 19431 4212 19440
rect 4160 19397 4169 19431
rect 4169 19397 4203 19431
rect 4203 19397 4212 19431
rect 4160 19388 4212 19397
rect 4436 19295 4488 19304
rect 4436 19261 4445 19295
rect 4445 19261 4479 19295
rect 4479 19261 4488 19295
rect 4436 19252 4488 19261
rect 4896 19363 4948 19372
rect 4896 19329 4905 19363
rect 4905 19329 4939 19363
rect 4939 19329 4948 19363
rect 4896 19320 4948 19329
rect 4988 19363 5040 19372
rect 4988 19329 4997 19363
rect 4997 19329 5031 19363
rect 5031 19329 5040 19363
rect 4988 19320 5040 19329
rect 5356 19499 5408 19508
rect 5356 19465 5365 19499
rect 5365 19465 5399 19499
rect 5399 19465 5408 19499
rect 5356 19456 5408 19465
rect 5448 19456 5500 19508
rect 12808 19456 12860 19508
rect 6184 19388 6236 19440
rect 6644 19431 6696 19440
rect 6644 19397 6653 19431
rect 6653 19397 6687 19431
rect 6687 19397 6696 19431
rect 6644 19388 6696 19397
rect 7012 19388 7064 19440
rect 5448 19252 5500 19304
rect 6000 19295 6052 19304
rect 6000 19261 6009 19295
rect 6009 19261 6043 19295
rect 6043 19261 6052 19295
rect 6000 19252 6052 19261
rect 5356 19184 5408 19236
rect 7932 19320 7984 19372
rect 7380 19295 7432 19304
rect 7380 19261 7389 19295
rect 7389 19261 7423 19295
rect 7423 19261 7432 19295
rect 7380 19252 7432 19261
rect 8116 19116 8168 19168
rect 8300 19116 8352 19168
rect 9036 19363 9088 19372
rect 9036 19329 9045 19363
rect 9045 19329 9079 19363
rect 9079 19329 9088 19363
rect 9036 19320 9088 19329
rect 9128 19363 9180 19372
rect 9128 19329 9137 19363
rect 9137 19329 9171 19363
rect 9171 19329 9180 19363
rect 9128 19320 9180 19329
rect 10692 19388 10744 19440
rect 14280 19456 14332 19508
rect 9864 19252 9916 19304
rect 10232 19320 10284 19372
rect 10692 19252 10744 19304
rect 9036 19116 9088 19168
rect 9864 19116 9916 19168
rect 11244 19320 11296 19372
rect 12440 19363 12492 19372
rect 12440 19329 12449 19363
rect 12449 19329 12483 19363
rect 12483 19329 12492 19363
rect 12440 19320 12492 19329
rect 12900 19320 12952 19372
rect 13728 19388 13780 19440
rect 13912 19388 13964 19440
rect 14740 19431 14792 19440
rect 14740 19397 14749 19431
rect 14749 19397 14783 19431
rect 14783 19397 14792 19431
rect 14740 19388 14792 19397
rect 14832 19431 14884 19440
rect 14832 19397 14841 19431
rect 14841 19397 14875 19431
rect 14875 19397 14884 19431
rect 14832 19388 14884 19397
rect 16672 19456 16724 19508
rect 15936 19431 15988 19440
rect 15936 19397 15945 19431
rect 15945 19397 15979 19431
rect 15979 19397 15988 19431
rect 15936 19388 15988 19397
rect 17592 19456 17644 19508
rect 20536 19456 20588 19508
rect 21272 19499 21324 19508
rect 21272 19465 21281 19499
rect 21281 19465 21315 19499
rect 21315 19465 21324 19499
rect 21272 19456 21324 19465
rect 21364 19456 21416 19508
rect 21916 19456 21968 19508
rect 22744 19456 22796 19508
rect 12716 19295 12768 19304
rect 12716 19261 12725 19295
rect 12725 19261 12759 19295
rect 12759 19261 12768 19295
rect 12716 19252 12768 19261
rect 12992 19184 13044 19236
rect 13452 19363 13504 19372
rect 13452 19329 13461 19363
rect 13461 19329 13495 19363
rect 13495 19329 13504 19363
rect 13452 19320 13504 19329
rect 14464 19320 14516 19372
rect 14648 19320 14700 19372
rect 15108 19320 15160 19372
rect 16304 19320 16356 19372
rect 16672 19363 16724 19372
rect 16672 19329 16681 19363
rect 16681 19329 16715 19363
rect 16715 19329 16724 19363
rect 16672 19320 16724 19329
rect 17040 19431 17092 19440
rect 17040 19397 17049 19431
rect 17049 19397 17083 19431
rect 17083 19397 17092 19431
rect 17040 19388 17092 19397
rect 18696 19388 18748 19440
rect 20076 19388 20128 19440
rect 17500 19320 17552 19372
rect 18144 19363 18196 19372
rect 18144 19329 18153 19363
rect 18153 19329 18187 19363
rect 18187 19329 18196 19363
rect 18144 19320 18196 19329
rect 19524 19320 19576 19372
rect 20628 19388 20680 19440
rect 21364 19320 21416 19372
rect 22376 19388 22428 19440
rect 24124 19456 24176 19508
rect 23664 19431 23716 19440
rect 23664 19397 23673 19431
rect 23673 19397 23707 19431
rect 23707 19397 23716 19431
rect 23664 19388 23716 19397
rect 23756 19363 23808 19372
rect 23756 19329 23765 19363
rect 23765 19329 23799 19363
rect 23799 19329 23808 19363
rect 23756 19320 23808 19329
rect 24860 19456 24912 19508
rect 26240 19456 26292 19508
rect 28080 19456 28132 19508
rect 28724 19456 28776 19508
rect 29092 19499 29144 19508
rect 29092 19465 29101 19499
rect 29101 19465 29135 19499
rect 29135 19465 29144 19499
rect 29092 19456 29144 19465
rect 29920 19456 29972 19508
rect 31208 19456 31260 19508
rect 13636 19252 13688 19304
rect 14372 19252 14424 19304
rect 14740 19252 14792 19304
rect 16028 19295 16080 19304
rect 16028 19261 16037 19295
rect 16037 19261 16071 19295
rect 16071 19261 16080 19295
rect 16028 19252 16080 19261
rect 16212 19252 16264 19304
rect 20444 19252 20496 19304
rect 21640 19252 21692 19304
rect 11060 19116 11112 19168
rect 12072 19159 12124 19168
rect 12072 19125 12081 19159
rect 12081 19125 12115 19159
rect 12115 19125 12124 19159
rect 12072 19116 12124 19125
rect 13360 19116 13412 19168
rect 15476 19159 15528 19168
rect 15476 19125 15485 19159
rect 15485 19125 15519 19159
rect 15519 19125 15528 19159
rect 15476 19116 15528 19125
rect 16028 19116 16080 19168
rect 17132 19116 17184 19168
rect 17500 19116 17552 19168
rect 18144 19116 18196 19168
rect 19616 19159 19668 19168
rect 19616 19125 19625 19159
rect 19625 19125 19659 19159
rect 19659 19125 19668 19159
rect 19616 19116 19668 19125
rect 20536 19116 20588 19168
rect 23112 19252 23164 19304
rect 25412 19320 25464 19372
rect 26424 19388 26476 19440
rect 28264 19388 28316 19440
rect 26608 19329 26625 19346
rect 26625 19329 26660 19346
rect 25964 19252 26016 19304
rect 26608 19294 26660 19329
rect 26792 19320 26844 19372
rect 29184 19388 29236 19440
rect 24032 19184 24084 19236
rect 22192 19116 22244 19168
rect 24400 19116 24452 19168
rect 25228 19184 25280 19236
rect 27804 19184 27856 19236
rect 25688 19116 25740 19168
rect 25872 19116 25924 19168
rect 26332 19116 26384 19168
rect 26424 19159 26476 19168
rect 26424 19125 26433 19159
rect 26433 19125 26467 19159
rect 26467 19125 26476 19159
rect 26424 19116 26476 19125
rect 27344 19159 27396 19168
rect 27344 19125 27353 19159
rect 27353 19125 27387 19159
rect 27387 19125 27396 19159
rect 27344 19116 27396 19125
rect 27896 19116 27948 19168
rect 28540 19252 28592 19304
rect 29000 19252 29052 19304
rect 29644 19363 29696 19372
rect 29644 19329 29653 19363
rect 29653 19329 29687 19363
rect 29687 19329 29696 19363
rect 29644 19320 29696 19329
rect 32128 19363 32180 19372
rect 32128 19329 32137 19363
rect 32137 19329 32171 19363
rect 32171 19329 32180 19363
rect 32128 19320 32180 19329
rect 29828 19252 29880 19304
rect 29092 19184 29144 19236
rect 30472 19295 30524 19304
rect 30472 19261 30481 19295
rect 30481 19261 30515 19295
rect 30515 19261 30524 19295
rect 30472 19252 30524 19261
rect 32864 19252 32916 19304
rect 34888 19252 34940 19304
rect 30564 19184 30616 19236
rect 29368 19116 29420 19168
rect 31024 19116 31076 19168
rect 32772 19116 32824 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 5448 18912 5500 18964
rect 7012 18955 7064 18964
rect 7012 18921 7021 18955
rect 7021 18921 7055 18955
rect 7055 18921 7064 18955
rect 7012 18912 7064 18921
rect 7932 18955 7984 18964
rect 7932 18921 7941 18955
rect 7941 18921 7975 18955
rect 7975 18921 7984 18955
rect 7932 18912 7984 18921
rect 12900 18955 12952 18964
rect 12900 18921 12909 18955
rect 12909 18921 12943 18955
rect 12943 18921 12952 18955
rect 12900 18912 12952 18921
rect 14280 18955 14332 18964
rect 14280 18921 14289 18955
rect 14289 18921 14323 18955
rect 14323 18921 14332 18955
rect 14280 18912 14332 18921
rect 14372 18912 14424 18964
rect 16212 18912 16264 18964
rect 16304 18955 16356 18964
rect 16304 18921 16313 18955
rect 16313 18921 16347 18955
rect 16347 18921 16356 18955
rect 16304 18912 16356 18921
rect 18236 18955 18288 18964
rect 18236 18921 18245 18955
rect 18245 18921 18279 18955
rect 18279 18921 18288 18955
rect 18236 18912 18288 18921
rect 19524 18912 19576 18964
rect 20444 18912 20496 18964
rect 21824 18955 21876 18964
rect 21824 18921 21833 18955
rect 21833 18921 21867 18955
rect 21867 18921 21876 18955
rect 21824 18912 21876 18921
rect 21916 18912 21968 18964
rect 23664 18912 23716 18964
rect 23756 18912 23808 18964
rect 25412 18955 25464 18964
rect 25412 18921 25421 18955
rect 25421 18921 25455 18955
rect 25455 18921 25464 18955
rect 25412 18912 25464 18921
rect 26240 18955 26292 18964
rect 26240 18921 26249 18955
rect 26249 18921 26283 18955
rect 26283 18921 26292 18955
rect 26240 18912 26292 18921
rect 26332 18955 26384 18964
rect 26332 18921 26341 18955
rect 26341 18921 26375 18955
rect 26375 18921 26384 18955
rect 26332 18912 26384 18921
rect 27344 18912 27396 18964
rect 27436 18955 27488 18964
rect 27436 18921 27445 18955
rect 27445 18921 27479 18955
rect 27479 18921 27488 18955
rect 27436 18912 27488 18921
rect 29000 18912 29052 18964
rect 30196 18912 30248 18964
rect 16028 18844 16080 18896
rect 19340 18844 19392 18896
rect 22652 18844 22704 18896
rect 23848 18844 23900 18896
rect 7932 18776 7984 18828
rect 9312 18776 9364 18828
rect 9404 18819 9456 18828
rect 9404 18785 9413 18819
rect 9413 18785 9447 18819
rect 9447 18785 9456 18819
rect 9404 18776 9456 18785
rect 9588 18819 9640 18828
rect 9588 18785 9597 18819
rect 9597 18785 9631 18819
rect 9631 18785 9640 18819
rect 9588 18776 9640 18785
rect 14924 18819 14976 18828
rect 14924 18785 14933 18819
rect 14933 18785 14967 18819
rect 14967 18785 14976 18819
rect 14924 18776 14976 18785
rect 17224 18819 17276 18828
rect 17224 18785 17233 18819
rect 17233 18785 17267 18819
rect 17267 18785 17276 18819
rect 17224 18776 17276 18785
rect 1308 18708 1360 18760
rect 3516 18708 3568 18760
rect 7012 18708 7064 18760
rect 3884 18640 3936 18692
rect 1768 18615 1820 18624
rect 1768 18581 1777 18615
rect 1777 18581 1811 18615
rect 1811 18581 1820 18615
rect 1768 18572 1820 18581
rect 4160 18572 4212 18624
rect 4896 18572 4948 18624
rect 5356 18615 5408 18624
rect 5356 18581 5365 18615
rect 5365 18581 5399 18615
rect 5399 18581 5408 18615
rect 5356 18572 5408 18581
rect 8300 18683 8352 18692
rect 8300 18649 8309 18683
rect 8309 18649 8343 18683
rect 8343 18649 8352 18683
rect 8300 18640 8352 18649
rect 8944 18615 8996 18624
rect 8944 18581 8953 18615
rect 8953 18581 8987 18615
rect 8987 18581 8996 18615
rect 8944 18572 8996 18581
rect 9128 18640 9180 18692
rect 9404 18640 9456 18692
rect 12072 18708 12124 18760
rect 12348 18708 12400 18760
rect 15476 18708 15528 18760
rect 10324 18640 10376 18692
rect 9680 18572 9732 18624
rect 12992 18640 13044 18692
rect 10692 18572 10744 18624
rect 13728 18572 13780 18624
rect 15844 18572 15896 18624
rect 17132 18751 17184 18760
rect 17132 18717 17141 18751
rect 17141 18717 17175 18751
rect 17175 18717 17184 18751
rect 17132 18708 17184 18717
rect 17408 18708 17460 18760
rect 17684 18683 17736 18692
rect 17684 18649 17693 18683
rect 17693 18649 17727 18683
rect 17727 18649 17736 18683
rect 17684 18640 17736 18649
rect 17960 18640 18012 18692
rect 18696 18819 18748 18828
rect 18696 18785 18705 18819
rect 18705 18785 18739 18819
rect 18739 18785 18748 18819
rect 18696 18776 18748 18785
rect 18880 18819 18932 18828
rect 18880 18785 18889 18819
rect 18889 18785 18923 18819
rect 18923 18785 18932 18819
rect 18880 18776 18932 18785
rect 18604 18751 18656 18760
rect 18604 18717 18613 18751
rect 18613 18717 18647 18751
rect 18647 18717 18656 18751
rect 18604 18708 18656 18717
rect 20536 18708 20588 18760
rect 20628 18751 20680 18760
rect 20628 18717 20637 18751
rect 20637 18717 20671 18751
rect 20671 18717 20680 18751
rect 20628 18708 20680 18717
rect 21548 18708 21600 18760
rect 22192 18751 22244 18760
rect 22192 18717 22201 18751
rect 22201 18717 22235 18751
rect 22235 18717 22244 18751
rect 22192 18708 22244 18717
rect 22284 18708 22336 18760
rect 25964 18776 26016 18828
rect 26424 18819 26476 18828
rect 26424 18785 26433 18819
rect 26433 18785 26467 18819
rect 26467 18785 26476 18819
rect 26424 18776 26476 18785
rect 26792 18776 26844 18828
rect 26700 18751 26752 18760
rect 26700 18717 26709 18751
rect 26709 18717 26743 18751
rect 26743 18717 26752 18751
rect 26700 18708 26752 18717
rect 27344 18776 27396 18828
rect 21548 18615 21600 18624
rect 21548 18581 21557 18615
rect 21557 18581 21591 18615
rect 21591 18581 21600 18615
rect 21548 18572 21600 18581
rect 21640 18572 21692 18624
rect 23296 18640 23348 18692
rect 26056 18683 26108 18692
rect 26056 18649 26065 18683
rect 26065 18649 26099 18683
rect 26099 18649 26108 18683
rect 26056 18640 26108 18649
rect 26240 18640 26292 18692
rect 27436 18751 27488 18760
rect 27436 18717 27445 18751
rect 27445 18717 27479 18751
rect 27479 18717 27488 18751
rect 27436 18708 27488 18717
rect 29184 18844 29236 18896
rect 29644 18776 29696 18828
rect 28540 18751 28592 18760
rect 28540 18717 28549 18751
rect 28549 18717 28583 18751
rect 28583 18717 28592 18751
rect 28540 18708 28592 18717
rect 29184 18708 29236 18760
rect 30380 18844 30432 18896
rect 32496 18955 32548 18964
rect 32496 18921 32505 18955
rect 32505 18921 32539 18955
rect 32539 18921 32548 18955
rect 32496 18912 32548 18921
rect 27896 18683 27948 18692
rect 23020 18572 23072 18624
rect 25964 18572 26016 18624
rect 26516 18572 26568 18624
rect 26792 18615 26844 18624
rect 26792 18581 26801 18615
rect 26801 18581 26835 18615
rect 26835 18581 26844 18615
rect 26792 18572 26844 18581
rect 27896 18649 27905 18683
rect 27905 18649 27939 18683
rect 27939 18649 27948 18683
rect 27896 18640 27948 18649
rect 28724 18640 28776 18692
rect 30472 18708 30524 18760
rect 28448 18615 28500 18624
rect 28448 18581 28457 18615
rect 28457 18581 28491 18615
rect 28491 18581 28500 18615
rect 28448 18572 28500 18581
rect 28908 18615 28960 18624
rect 28908 18581 28917 18615
rect 28917 18581 28951 18615
rect 28951 18581 28960 18615
rect 28908 18572 28960 18581
rect 29368 18640 29420 18692
rect 29552 18572 29604 18624
rect 30012 18572 30064 18624
rect 30104 18572 30156 18624
rect 30288 18572 30340 18624
rect 31024 18819 31076 18828
rect 31024 18785 31033 18819
rect 31033 18785 31067 18819
rect 31067 18785 31076 18819
rect 31024 18776 31076 18785
rect 32220 18776 32272 18828
rect 32588 18776 32640 18828
rect 30748 18751 30800 18760
rect 30748 18717 30757 18751
rect 30757 18717 30791 18751
rect 30791 18717 30800 18751
rect 30748 18708 30800 18717
rect 32772 18751 32824 18760
rect 32772 18717 32781 18751
rect 32781 18717 32815 18751
rect 32815 18717 32824 18751
rect 32772 18708 32824 18717
rect 34152 18751 34204 18760
rect 34152 18717 34161 18751
rect 34161 18717 34195 18751
rect 34195 18717 34204 18751
rect 34152 18708 34204 18717
rect 31760 18572 31812 18624
rect 33692 18572 33744 18624
rect 33784 18572 33836 18624
rect 34520 18572 34572 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 3884 18368 3936 18420
rect 4160 18411 4212 18420
rect 4160 18377 4169 18411
rect 4169 18377 4203 18411
rect 4203 18377 4212 18411
rect 4160 18368 4212 18377
rect 5448 18368 5500 18420
rect 7104 18368 7156 18420
rect 6000 18300 6052 18352
rect 7380 18232 7432 18284
rect 8944 18300 8996 18352
rect 9128 18411 9180 18420
rect 9128 18377 9137 18411
rect 9137 18377 9171 18411
rect 9171 18377 9180 18411
rect 9128 18368 9180 18377
rect 9588 18368 9640 18420
rect 10324 18411 10376 18420
rect 10324 18377 10333 18411
rect 10333 18377 10367 18411
rect 10367 18377 10376 18411
rect 10324 18368 10376 18377
rect 10692 18411 10744 18420
rect 10692 18377 10701 18411
rect 10701 18377 10735 18411
rect 10735 18377 10744 18411
rect 10692 18368 10744 18377
rect 10784 18411 10836 18420
rect 10784 18377 10793 18411
rect 10793 18377 10827 18411
rect 10827 18377 10836 18411
rect 10784 18368 10836 18377
rect 12716 18368 12768 18420
rect 10416 18300 10468 18352
rect 13360 18343 13412 18352
rect 10324 18232 10376 18284
rect 4712 18164 4764 18216
rect 5264 18164 5316 18216
rect 13360 18309 13394 18343
rect 13394 18309 13412 18343
rect 13360 18300 13412 18309
rect 14004 18300 14056 18352
rect 14464 18411 14516 18420
rect 14464 18377 14473 18411
rect 14473 18377 14507 18411
rect 14507 18377 14516 18411
rect 14464 18368 14516 18377
rect 21548 18368 21600 18420
rect 22192 18368 22244 18420
rect 22468 18368 22520 18420
rect 22652 18411 22704 18420
rect 22652 18377 22661 18411
rect 22661 18377 22695 18411
rect 22695 18377 22704 18411
rect 22652 18368 22704 18377
rect 23204 18411 23256 18420
rect 23204 18377 23213 18411
rect 23213 18377 23247 18411
rect 23247 18377 23256 18411
rect 23204 18368 23256 18377
rect 23296 18411 23348 18420
rect 23296 18377 23305 18411
rect 23305 18377 23339 18411
rect 23339 18377 23348 18411
rect 23296 18368 23348 18377
rect 23664 18411 23716 18420
rect 23664 18377 23673 18411
rect 23673 18377 23707 18411
rect 23707 18377 23716 18411
rect 23664 18368 23716 18377
rect 23756 18411 23808 18420
rect 23756 18377 23765 18411
rect 23765 18377 23799 18411
rect 23799 18377 23808 18411
rect 23756 18368 23808 18377
rect 25412 18368 25464 18420
rect 25688 18368 25740 18420
rect 12072 18164 12124 18216
rect 13084 18207 13136 18216
rect 13084 18173 13093 18207
rect 13093 18173 13127 18207
rect 13127 18173 13136 18207
rect 13084 18164 13136 18173
rect 9864 18096 9916 18148
rect 7932 18028 7984 18080
rect 9312 18071 9364 18080
rect 9312 18037 9321 18071
rect 9321 18037 9355 18071
rect 9355 18037 9364 18071
rect 9312 18028 9364 18037
rect 9588 18028 9640 18080
rect 14096 18096 14148 18148
rect 14372 18096 14424 18148
rect 15108 18164 15160 18216
rect 14004 18028 14056 18080
rect 16580 18232 16632 18284
rect 16948 18275 17000 18284
rect 16948 18241 16982 18275
rect 16982 18241 17000 18275
rect 16948 18232 17000 18241
rect 21732 18300 21784 18352
rect 22928 18300 22980 18352
rect 21548 18207 21600 18216
rect 21548 18173 21557 18207
rect 21557 18173 21591 18207
rect 21591 18173 21600 18207
rect 21548 18164 21600 18173
rect 22744 18207 22796 18216
rect 22744 18173 22753 18207
rect 22753 18173 22787 18207
rect 22787 18173 22796 18207
rect 22744 18164 22796 18173
rect 23020 18164 23072 18216
rect 25136 18300 25188 18352
rect 24860 18232 24912 18284
rect 25228 18275 25280 18284
rect 25228 18241 25237 18275
rect 25237 18241 25271 18275
rect 25271 18241 25280 18275
rect 25228 18232 25280 18241
rect 26056 18300 26108 18352
rect 26332 18411 26384 18420
rect 26332 18377 26341 18411
rect 26341 18377 26375 18411
rect 26375 18377 26384 18411
rect 26332 18368 26384 18377
rect 29092 18368 29144 18420
rect 25320 18207 25372 18216
rect 25320 18173 25329 18207
rect 25329 18173 25363 18207
rect 25363 18173 25372 18207
rect 25320 18164 25372 18173
rect 19616 18096 19668 18148
rect 24768 18096 24820 18148
rect 24860 18096 24912 18148
rect 26608 18300 26660 18352
rect 27068 18300 27120 18352
rect 27436 18300 27488 18352
rect 29644 18368 29696 18420
rect 29552 18300 29604 18352
rect 30932 18300 30984 18352
rect 27620 18275 27672 18284
rect 27620 18241 27629 18275
rect 27629 18241 27663 18275
rect 27663 18241 27672 18275
rect 27620 18232 27672 18241
rect 28908 18232 28960 18284
rect 29092 18232 29144 18284
rect 30012 18232 30064 18284
rect 25412 18096 25464 18148
rect 25872 18096 25924 18148
rect 28540 18164 28592 18216
rect 26700 18096 26752 18148
rect 30104 18207 30156 18216
rect 30104 18173 30113 18207
rect 30113 18173 30147 18207
rect 30147 18173 30156 18207
rect 30104 18164 30156 18173
rect 32128 18368 32180 18420
rect 31760 18300 31812 18352
rect 32772 18368 32824 18420
rect 33140 18300 33192 18352
rect 33692 18343 33744 18352
rect 33692 18309 33701 18343
rect 33701 18309 33735 18343
rect 33735 18309 33744 18343
rect 33692 18300 33744 18309
rect 31668 18275 31720 18284
rect 31668 18241 31677 18275
rect 31677 18241 31711 18275
rect 31711 18241 31720 18275
rect 31668 18232 31720 18241
rect 34520 18275 34572 18284
rect 34520 18241 34529 18275
rect 34529 18241 34563 18275
rect 34563 18241 34572 18275
rect 34520 18232 34572 18241
rect 34796 18275 34848 18284
rect 34796 18241 34805 18275
rect 34805 18241 34839 18275
rect 34839 18241 34848 18275
rect 34796 18232 34848 18241
rect 30564 18096 30616 18148
rect 31576 18096 31628 18148
rect 16304 18028 16356 18080
rect 17316 18028 17368 18080
rect 18880 18028 18932 18080
rect 22100 18028 22152 18080
rect 22192 18028 22244 18080
rect 24584 18028 24636 18080
rect 24676 18028 24728 18080
rect 28724 18071 28776 18080
rect 28724 18037 28733 18071
rect 28733 18037 28767 18071
rect 28767 18037 28776 18071
rect 28724 18028 28776 18037
rect 29276 18028 29328 18080
rect 29644 18028 29696 18080
rect 29828 18028 29880 18080
rect 31300 18028 31352 18080
rect 32680 18028 32732 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1768 17824 1820 17876
rect 7196 17756 7248 17808
rect 11888 17756 11940 17808
rect 15108 17756 15160 17808
rect 16948 17824 17000 17876
rect 17132 17824 17184 17876
rect 10324 17688 10376 17740
rect 16856 17688 16908 17740
rect 17132 17688 17184 17740
rect 17316 17731 17368 17740
rect 17316 17697 17325 17731
rect 17325 17697 17359 17731
rect 17359 17697 17368 17731
rect 17316 17688 17368 17697
rect 17592 17688 17644 17740
rect 7748 17620 7800 17672
rect 10692 17552 10744 17604
rect 7380 17484 7432 17536
rect 9312 17484 9364 17536
rect 9864 17527 9916 17536
rect 9864 17493 9873 17527
rect 9873 17493 9907 17527
rect 9907 17493 9916 17527
rect 9864 17484 9916 17493
rect 10876 17484 10928 17536
rect 11152 17595 11204 17604
rect 11152 17561 11161 17595
rect 11161 17561 11195 17595
rect 11195 17561 11204 17595
rect 11152 17552 11204 17561
rect 11428 17527 11480 17536
rect 11428 17493 11437 17527
rect 11437 17493 11471 17527
rect 11471 17493 11480 17527
rect 11428 17484 11480 17493
rect 11612 17527 11664 17536
rect 11612 17493 11621 17527
rect 11621 17493 11655 17527
rect 11655 17493 11664 17527
rect 11612 17484 11664 17493
rect 12440 17527 12492 17536
rect 12440 17493 12449 17527
rect 12449 17493 12483 17527
rect 12483 17493 12492 17527
rect 14924 17620 14976 17672
rect 16764 17620 16816 17672
rect 22376 17824 22428 17876
rect 25412 17824 25464 17876
rect 24860 17688 24912 17740
rect 25228 17756 25280 17808
rect 14648 17552 14700 17604
rect 17500 17552 17552 17604
rect 22284 17663 22336 17672
rect 22284 17629 22293 17663
rect 22293 17629 22327 17663
rect 22327 17629 22336 17663
rect 22284 17620 22336 17629
rect 19892 17552 19944 17604
rect 12440 17484 12492 17493
rect 12992 17484 13044 17536
rect 14280 17484 14332 17536
rect 14832 17484 14884 17536
rect 17592 17484 17644 17536
rect 18972 17484 19024 17536
rect 22468 17552 22520 17604
rect 24952 17552 25004 17604
rect 25136 17731 25188 17740
rect 25136 17697 25145 17731
rect 25145 17697 25179 17731
rect 25179 17697 25188 17731
rect 25136 17688 25188 17697
rect 25872 17824 25924 17876
rect 25964 17867 26016 17876
rect 25964 17833 25973 17867
rect 25973 17833 26007 17867
rect 26007 17833 26016 17867
rect 25964 17824 26016 17833
rect 26148 17824 26200 17876
rect 29184 17824 29236 17876
rect 34520 17867 34572 17876
rect 34520 17833 34529 17867
rect 34529 17833 34563 17867
rect 34563 17833 34572 17867
rect 34520 17824 34572 17833
rect 26332 17688 26384 17740
rect 28264 17756 28316 17808
rect 27068 17731 27120 17740
rect 27068 17697 27077 17731
rect 27077 17697 27111 17731
rect 27111 17697 27120 17731
rect 27068 17688 27120 17697
rect 27344 17731 27396 17740
rect 27344 17697 27353 17731
rect 27353 17697 27387 17731
rect 27387 17697 27396 17731
rect 27344 17688 27396 17697
rect 26424 17620 26476 17672
rect 20720 17527 20772 17536
rect 20720 17493 20729 17527
rect 20729 17493 20763 17527
rect 20763 17493 20772 17527
rect 20720 17484 20772 17493
rect 22100 17484 22152 17536
rect 22744 17484 22796 17536
rect 23940 17484 23992 17536
rect 24124 17484 24176 17536
rect 25136 17484 25188 17536
rect 25320 17484 25372 17536
rect 27620 17688 27672 17740
rect 27712 17620 27764 17672
rect 29552 17688 29604 17740
rect 30012 17731 30064 17740
rect 30012 17697 30021 17731
rect 30021 17697 30055 17731
rect 30055 17697 30064 17731
rect 30012 17688 30064 17697
rect 28448 17620 28500 17672
rect 27712 17527 27764 17536
rect 27712 17493 27721 17527
rect 27721 17493 27755 17527
rect 27755 17493 27764 17527
rect 27712 17484 27764 17493
rect 28264 17552 28316 17604
rect 29644 17620 29696 17672
rect 29828 17620 29880 17672
rect 30196 17663 30248 17672
rect 30196 17629 30205 17663
rect 30205 17629 30239 17663
rect 30239 17629 30248 17663
rect 30196 17620 30248 17629
rect 30932 17620 30984 17672
rect 31208 17756 31260 17808
rect 33784 17688 33836 17740
rect 31576 17663 31628 17672
rect 31576 17629 31585 17663
rect 31585 17629 31619 17663
rect 31619 17629 31628 17663
rect 31576 17620 31628 17629
rect 32128 17620 32180 17672
rect 32680 17620 32732 17672
rect 31300 17595 31352 17604
rect 31300 17561 31309 17595
rect 31309 17561 31343 17595
rect 31343 17561 31352 17595
rect 31300 17552 31352 17561
rect 33140 17552 33192 17604
rect 29000 17484 29052 17536
rect 31024 17484 31076 17536
rect 31484 17527 31536 17536
rect 31484 17493 31493 17527
rect 31493 17493 31527 17527
rect 31527 17493 31536 17527
rect 31484 17484 31536 17493
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 4620 17212 4672 17264
rect 4988 17280 5040 17332
rect 5264 17280 5316 17332
rect 4068 17144 4120 17196
rect 6736 17187 6788 17196
rect 6736 17153 6745 17187
rect 6745 17153 6779 17187
rect 6779 17153 6788 17187
rect 7748 17323 7800 17332
rect 7748 17289 7757 17323
rect 7757 17289 7791 17323
rect 7791 17289 7800 17323
rect 7748 17280 7800 17289
rect 9496 17280 9548 17332
rect 10692 17323 10744 17332
rect 10692 17289 10701 17323
rect 10701 17289 10735 17323
rect 10735 17289 10744 17323
rect 10692 17280 10744 17289
rect 11152 17280 11204 17332
rect 12256 17280 12308 17332
rect 14280 17323 14332 17332
rect 14280 17289 14289 17323
rect 14289 17289 14323 17323
rect 14323 17289 14332 17323
rect 14280 17280 14332 17289
rect 14648 17323 14700 17332
rect 14648 17289 14657 17323
rect 14657 17289 14691 17323
rect 14691 17289 14700 17323
rect 14648 17280 14700 17289
rect 14740 17280 14792 17332
rect 15108 17280 15160 17332
rect 9864 17212 9916 17264
rect 6736 17144 6788 17153
rect 3516 17119 3568 17128
rect 3516 17085 3525 17119
rect 3525 17085 3559 17119
rect 3559 17085 3568 17119
rect 3516 17076 3568 17085
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 7012 17119 7064 17128
rect 7012 17085 7021 17119
rect 7021 17085 7055 17119
rect 7055 17085 7064 17119
rect 7012 17076 7064 17085
rect 5724 17008 5776 17060
rect 9312 17187 9364 17196
rect 9312 17153 9321 17187
rect 9321 17153 9355 17187
rect 9355 17153 9364 17187
rect 9312 17144 9364 17153
rect 13084 17212 13136 17264
rect 14188 17212 14240 17264
rect 19892 17323 19944 17332
rect 19892 17289 19901 17323
rect 19901 17289 19935 17323
rect 19935 17289 19944 17323
rect 19892 17280 19944 17289
rect 21548 17280 21600 17332
rect 11796 17187 11848 17196
rect 11796 17153 11830 17187
rect 11830 17153 11848 17187
rect 11796 17144 11848 17153
rect 12072 17144 12124 17196
rect 14648 17144 14700 17196
rect 14740 17187 14792 17196
rect 14740 17153 14749 17187
rect 14749 17153 14783 17187
rect 14783 17153 14792 17187
rect 14740 17144 14792 17153
rect 11520 17119 11572 17128
rect 11520 17085 11529 17119
rect 11529 17085 11563 17119
rect 11563 17085 11572 17119
rect 11520 17076 11572 17085
rect 13820 17076 13872 17128
rect 14096 17119 14148 17128
rect 14096 17085 14105 17119
rect 14105 17085 14139 17119
rect 14139 17085 14148 17119
rect 14096 17076 14148 17085
rect 14188 17119 14240 17128
rect 14188 17085 14197 17119
rect 14197 17085 14231 17119
rect 14231 17085 14240 17119
rect 14188 17076 14240 17085
rect 14556 17076 14608 17128
rect 15752 17144 15804 17196
rect 17500 17187 17552 17196
rect 17500 17153 17509 17187
rect 17509 17153 17543 17187
rect 17543 17153 17552 17187
rect 17500 17144 17552 17153
rect 18052 17144 18104 17196
rect 8484 17051 8536 17060
rect 6368 16983 6420 16992
rect 6368 16949 6377 16983
rect 6377 16949 6411 16983
rect 6411 16949 6420 16983
rect 6368 16940 6420 16949
rect 8484 17017 8493 17051
rect 8493 17017 8527 17051
rect 8527 17017 8536 17051
rect 8484 17008 8536 17017
rect 9036 17008 9088 17060
rect 10324 16940 10376 16992
rect 13084 17008 13136 17060
rect 16580 17008 16632 17060
rect 19340 17212 19392 17264
rect 20536 17212 20588 17264
rect 18972 17187 19024 17196
rect 18972 17153 18981 17187
rect 18981 17153 19015 17187
rect 19015 17153 19024 17187
rect 18972 17144 19024 17153
rect 20720 17144 20772 17196
rect 19800 17076 19852 17128
rect 21548 17051 21600 17060
rect 21548 17017 21557 17051
rect 21557 17017 21591 17051
rect 21591 17017 21600 17051
rect 21548 17008 21600 17017
rect 16488 16983 16540 16992
rect 16488 16949 16497 16983
rect 16497 16949 16531 16983
rect 16531 16949 16540 16983
rect 16488 16940 16540 16949
rect 18880 16983 18932 16992
rect 18880 16949 18889 16983
rect 18889 16949 18923 16983
rect 18923 16949 18932 16983
rect 18880 16940 18932 16949
rect 20168 16940 20220 16992
rect 20996 16940 21048 16992
rect 22100 17255 22152 17264
rect 22100 17221 22109 17255
rect 22109 17221 22143 17255
rect 22143 17221 22152 17255
rect 22100 17212 22152 17221
rect 22652 17280 22704 17332
rect 24860 17280 24912 17332
rect 27068 17280 27120 17332
rect 24584 17212 24636 17264
rect 26608 17212 26660 17264
rect 27252 17212 27304 17264
rect 23112 17144 23164 17196
rect 23388 17187 23440 17196
rect 23388 17153 23397 17187
rect 23397 17153 23431 17187
rect 23431 17153 23440 17187
rect 23388 17144 23440 17153
rect 22376 17076 22428 17128
rect 23940 17119 23992 17128
rect 23940 17085 23949 17119
rect 23949 17085 23983 17119
rect 23983 17085 23992 17119
rect 23940 17076 23992 17085
rect 24032 17119 24084 17128
rect 24032 17085 24041 17119
rect 24041 17085 24075 17119
rect 24075 17085 24084 17119
rect 24032 17076 24084 17085
rect 24584 17076 24636 17128
rect 25136 17187 25188 17196
rect 25136 17153 25145 17187
rect 25145 17153 25179 17187
rect 25179 17153 25188 17187
rect 25136 17144 25188 17153
rect 26332 17144 26384 17196
rect 24952 17076 25004 17128
rect 27344 17076 27396 17128
rect 22376 16983 22428 16992
rect 22376 16949 22385 16983
rect 22385 16949 22419 16983
rect 22419 16949 22428 16983
rect 22376 16940 22428 16949
rect 23480 16983 23532 16992
rect 23480 16949 23489 16983
rect 23489 16949 23523 16983
rect 23523 16949 23532 16983
rect 23480 16940 23532 16949
rect 23848 16940 23900 16992
rect 26884 17008 26936 17060
rect 24308 16983 24360 16992
rect 24308 16949 24317 16983
rect 24317 16949 24351 16983
rect 24351 16949 24360 16983
rect 24308 16940 24360 16949
rect 25596 16940 25648 16992
rect 27804 17076 27856 17128
rect 28632 17119 28684 17128
rect 28632 17085 28641 17119
rect 28641 17085 28675 17119
rect 28675 17085 28684 17119
rect 28632 17076 28684 17085
rect 30104 17323 30156 17332
rect 30104 17289 30113 17323
rect 30113 17289 30147 17323
rect 30147 17289 30156 17323
rect 30104 17280 30156 17289
rect 30932 17280 30984 17332
rect 31300 17280 31352 17332
rect 29828 17076 29880 17128
rect 29276 16940 29328 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 5356 16736 5408 16788
rect 5540 16736 5592 16788
rect 6736 16779 6788 16788
rect 6736 16745 6745 16779
rect 6745 16745 6779 16779
rect 6779 16745 6788 16779
rect 6736 16736 6788 16745
rect 7012 16736 7064 16788
rect 9680 16736 9732 16788
rect 5356 16643 5408 16652
rect 1400 16575 1452 16584
rect 1400 16541 1409 16575
rect 1409 16541 1443 16575
rect 1443 16541 1452 16575
rect 1400 16532 1452 16541
rect 2780 16464 2832 16516
rect 3516 16464 3568 16516
rect 5356 16609 5365 16643
rect 5365 16609 5399 16643
rect 5399 16609 5408 16643
rect 5356 16600 5408 16609
rect 7380 16643 7432 16652
rect 7380 16609 7389 16643
rect 7389 16609 7423 16643
rect 7423 16609 7432 16643
rect 7380 16600 7432 16609
rect 9312 16600 9364 16652
rect 11520 16600 11572 16652
rect 12440 16736 12492 16788
rect 13636 16711 13688 16720
rect 13636 16677 13645 16711
rect 13645 16677 13679 16711
rect 13679 16677 13688 16711
rect 13636 16668 13688 16677
rect 6368 16532 6420 16584
rect 1584 16439 1636 16448
rect 1584 16405 1593 16439
rect 1593 16405 1627 16439
rect 1627 16405 1636 16439
rect 1584 16396 1636 16405
rect 11888 16600 11940 16652
rect 13820 16600 13872 16652
rect 14004 16736 14056 16788
rect 14556 16736 14608 16788
rect 14648 16736 14700 16788
rect 14188 16668 14240 16720
rect 15016 16668 15068 16720
rect 15292 16711 15344 16720
rect 15292 16677 15301 16711
rect 15301 16677 15335 16711
rect 15335 16677 15344 16711
rect 15292 16668 15344 16677
rect 14740 16600 14792 16652
rect 15752 16779 15804 16788
rect 15752 16745 15761 16779
rect 15761 16745 15795 16779
rect 15795 16745 15804 16779
rect 15752 16736 15804 16745
rect 18052 16779 18104 16788
rect 18052 16745 18061 16779
rect 18061 16745 18095 16779
rect 18095 16745 18104 16779
rect 18052 16736 18104 16745
rect 19340 16668 19392 16720
rect 19156 16600 19208 16652
rect 19892 16600 19944 16652
rect 13636 16532 13688 16584
rect 8024 16464 8076 16516
rect 11152 16464 11204 16516
rect 14556 16575 14608 16584
rect 14556 16541 14565 16575
rect 14565 16541 14599 16575
rect 14599 16541 14608 16575
rect 14556 16532 14608 16541
rect 14648 16532 14700 16584
rect 14832 16575 14884 16584
rect 14832 16541 14841 16575
rect 14841 16541 14875 16575
rect 14875 16541 14884 16575
rect 14832 16532 14884 16541
rect 15108 16532 15160 16584
rect 15936 16532 15988 16584
rect 16488 16532 16540 16584
rect 16580 16575 16632 16584
rect 16580 16541 16589 16575
rect 16589 16541 16623 16575
rect 16623 16541 16632 16575
rect 17224 16575 17276 16584
rect 16580 16532 16632 16541
rect 17224 16541 17233 16575
rect 17233 16541 17267 16575
rect 17267 16541 17276 16575
rect 17224 16532 17276 16541
rect 18880 16532 18932 16584
rect 21456 16736 21508 16788
rect 22100 16736 22152 16788
rect 27068 16779 27120 16788
rect 27068 16745 27077 16779
rect 27077 16745 27111 16779
rect 27111 16745 27120 16779
rect 27068 16736 27120 16745
rect 28632 16736 28684 16788
rect 29736 16779 29788 16788
rect 29736 16745 29745 16779
rect 29745 16745 29779 16779
rect 29779 16745 29788 16779
rect 29736 16736 29788 16745
rect 30196 16779 30248 16788
rect 30196 16745 30205 16779
rect 30205 16745 30239 16779
rect 30239 16745 30248 16779
rect 30196 16736 30248 16745
rect 30840 16736 30892 16788
rect 23940 16668 23992 16720
rect 25320 16668 25372 16720
rect 20628 16600 20680 16652
rect 24032 16600 24084 16652
rect 24400 16643 24452 16652
rect 24400 16609 24409 16643
rect 24409 16609 24443 16643
rect 24443 16609 24452 16643
rect 24400 16600 24452 16609
rect 6460 16396 6512 16448
rect 8944 16396 8996 16448
rect 15200 16396 15252 16448
rect 16212 16439 16264 16448
rect 16212 16405 16221 16439
rect 16221 16405 16255 16439
rect 16255 16405 16264 16439
rect 16212 16396 16264 16405
rect 16764 16439 16816 16448
rect 16764 16405 16773 16439
rect 16773 16405 16807 16439
rect 16807 16405 16816 16439
rect 16764 16396 16816 16405
rect 19340 16396 19392 16448
rect 22192 16532 22244 16584
rect 22284 16575 22336 16584
rect 22284 16541 22293 16575
rect 22293 16541 22327 16575
rect 22327 16541 22336 16575
rect 22284 16532 22336 16541
rect 23480 16532 23532 16584
rect 24492 16532 24544 16584
rect 25320 16575 25372 16584
rect 25320 16541 25329 16575
rect 25329 16541 25363 16575
rect 25363 16541 25372 16575
rect 25320 16532 25372 16541
rect 25596 16600 25648 16652
rect 26148 16668 26200 16720
rect 26608 16643 26660 16652
rect 26608 16609 26617 16643
rect 26617 16609 26651 16643
rect 26651 16609 26660 16643
rect 26608 16600 26660 16609
rect 29000 16600 29052 16652
rect 26516 16532 26568 16584
rect 27344 16532 27396 16584
rect 28080 16532 28132 16584
rect 28724 16532 28776 16584
rect 28908 16575 28960 16584
rect 28908 16541 28917 16575
rect 28917 16541 28951 16575
rect 28951 16541 28960 16575
rect 28908 16532 28960 16541
rect 29552 16575 29604 16584
rect 29552 16541 29561 16575
rect 29561 16541 29595 16575
rect 29595 16541 29604 16575
rect 29552 16532 29604 16541
rect 30012 16575 30064 16584
rect 30012 16541 30021 16575
rect 30021 16541 30055 16575
rect 30055 16541 30064 16575
rect 31484 16600 31536 16652
rect 30012 16532 30064 16541
rect 30380 16532 30432 16584
rect 30748 16575 30800 16584
rect 30748 16541 30757 16575
rect 30757 16541 30791 16575
rect 30791 16541 30800 16575
rect 30748 16532 30800 16541
rect 32864 16532 32916 16584
rect 34060 16575 34112 16584
rect 34060 16541 34069 16575
rect 34069 16541 34103 16575
rect 34103 16541 34112 16575
rect 34060 16532 34112 16541
rect 23388 16464 23440 16516
rect 23940 16507 23992 16516
rect 23940 16473 23949 16507
rect 23949 16473 23983 16507
rect 23983 16473 23992 16507
rect 23940 16464 23992 16473
rect 22100 16396 22152 16448
rect 25412 16464 25464 16516
rect 24584 16396 24636 16448
rect 25872 16439 25924 16448
rect 25872 16405 25881 16439
rect 25881 16405 25915 16439
rect 25915 16405 25924 16439
rect 25872 16396 25924 16405
rect 26056 16439 26108 16448
rect 26056 16405 26065 16439
rect 26065 16405 26099 16439
rect 26099 16405 26108 16439
rect 26056 16396 26108 16405
rect 26424 16439 26476 16448
rect 26424 16405 26433 16439
rect 26433 16405 26467 16439
rect 26467 16405 26476 16439
rect 26424 16396 26476 16405
rect 27436 16439 27488 16448
rect 27436 16405 27445 16439
rect 27445 16405 27479 16439
rect 27479 16405 27488 16439
rect 27436 16396 27488 16405
rect 29092 16439 29144 16448
rect 29092 16405 29101 16439
rect 29101 16405 29135 16439
rect 29135 16405 29144 16439
rect 29092 16396 29144 16405
rect 29276 16439 29328 16448
rect 29276 16405 29285 16439
rect 29285 16405 29319 16439
rect 29319 16405 29328 16439
rect 29276 16396 29328 16405
rect 30932 16464 30984 16516
rect 33140 16464 33192 16516
rect 34336 16507 34388 16516
rect 34336 16473 34345 16507
rect 34345 16473 34379 16507
rect 34379 16473 34388 16507
rect 34336 16464 34388 16473
rect 31668 16396 31720 16448
rect 32588 16439 32640 16448
rect 32588 16405 32597 16439
rect 32597 16405 32631 16439
rect 32631 16405 32640 16439
rect 32588 16396 32640 16405
rect 32956 16439 33008 16448
rect 32956 16405 32965 16439
rect 32965 16405 32999 16439
rect 32999 16405 33008 16439
rect 32956 16396 33008 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 4068 16235 4120 16244
rect 4068 16201 4077 16235
rect 4077 16201 4111 16235
rect 4111 16201 4120 16235
rect 4068 16192 4120 16201
rect 4620 16192 4672 16244
rect 8024 16235 8076 16244
rect 8024 16201 8033 16235
rect 8033 16201 8067 16235
rect 8067 16201 8076 16235
rect 8024 16192 8076 16201
rect 11152 16192 11204 16244
rect 11796 16235 11848 16244
rect 11796 16201 11805 16235
rect 11805 16201 11839 16235
rect 11839 16201 11848 16235
rect 11796 16192 11848 16201
rect 12256 16235 12308 16244
rect 12256 16201 12265 16235
rect 12265 16201 12299 16235
rect 12299 16201 12308 16235
rect 12256 16192 12308 16201
rect 12716 16235 12768 16244
rect 12716 16201 12725 16235
rect 12725 16201 12759 16235
rect 12759 16201 12768 16235
rect 12716 16192 12768 16201
rect 1584 16056 1636 16108
rect 5356 16056 5408 16108
rect 6644 16099 6696 16108
rect 6644 16065 6678 16099
rect 6678 16065 6696 16099
rect 6644 16056 6696 16065
rect 7564 16056 7616 16108
rect 8944 16099 8996 16108
rect 8944 16065 8954 16099
rect 8954 16065 8988 16099
rect 8988 16065 8996 16099
rect 8944 16056 8996 16065
rect 4068 15852 4120 15904
rect 4712 16031 4764 16040
rect 4712 15997 4721 16031
rect 4721 15997 4755 16031
rect 4755 15997 4764 16031
rect 4712 15988 4764 15997
rect 9036 15988 9088 16040
rect 9220 16099 9272 16108
rect 9220 16065 9229 16099
rect 9229 16065 9263 16099
rect 9263 16065 9272 16099
rect 9220 16056 9272 16065
rect 9404 16056 9456 16108
rect 10876 16099 10928 16108
rect 10876 16065 10885 16099
rect 10885 16065 10919 16099
rect 10919 16065 10928 16099
rect 10876 16056 10928 16065
rect 11152 16099 11204 16108
rect 11152 16065 11161 16099
rect 11161 16065 11195 16099
rect 11195 16065 11204 16099
rect 11152 16056 11204 16065
rect 6736 15852 6788 15904
rect 7748 15895 7800 15904
rect 7748 15861 7757 15895
rect 7757 15861 7791 15895
rect 7791 15861 7800 15895
rect 7748 15852 7800 15861
rect 11336 15920 11388 15972
rect 9772 15852 9824 15904
rect 13084 16099 13136 16108
rect 13084 16065 13093 16099
rect 13093 16065 13127 16099
rect 13127 16065 13136 16099
rect 13084 16056 13136 16065
rect 15108 16192 15160 16244
rect 15660 16192 15712 16244
rect 16120 16192 16172 16244
rect 17960 16192 18012 16244
rect 15936 16167 15988 16176
rect 15936 16133 15945 16167
rect 15945 16133 15979 16167
rect 15979 16133 15988 16167
rect 15936 16124 15988 16133
rect 22100 16192 22152 16244
rect 22376 16192 22428 16244
rect 22468 16192 22520 16244
rect 25412 16192 25464 16244
rect 13728 16056 13780 16108
rect 14096 16056 14148 16108
rect 12716 15988 12768 16040
rect 14556 16056 14608 16108
rect 15200 16056 15252 16108
rect 15660 16099 15712 16108
rect 15660 16065 15670 16099
rect 15670 16065 15704 16099
rect 15704 16065 15712 16099
rect 15660 16056 15712 16065
rect 15016 16031 15068 16040
rect 15016 15997 15025 16031
rect 15025 15997 15059 16031
rect 15059 15997 15068 16031
rect 15016 15988 15068 15997
rect 15108 16031 15160 16040
rect 15108 15997 15117 16031
rect 15117 15997 15151 16031
rect 15151 15997 15160 16031
rect 15108 15988 15160 15997
rect 15384 15988 15436 16040
rect 16764 16056 16816 16108
rect 17500 16056 17552 16108
rect 18788 16099 18840 16108
rect 18788 16065 18795 16099
rect 18795 16065 18840 16099
rect 18788 16056 18840 16065
rect 18972 16099 19024 16108
rect 18972 16065 18981 16099
rect 18981 16065 19015 16099
rect 19015 16065 19024 16099
rect 18972 16056 19024 16065
rect 19248 16056 19300 16108
rect 20076 16056 20128 16108
rect 21456 16056 21508 16108
rect 22284 16124 22336 16176
rect 19340 15988 19392 16040
rect 19432 15988 19484 16040
rect 22192 16099 22244 16108
rect 22192 16065 22201 16099
rect 22201 16065 22235 16099
rect 22235 16065 22244 16099
rect 22468 16099 22520 16108
rect 22192 16056 22244 16065
rect 22468 16065 22477 16099
rect 22477 16065 22511 16099
rect 22511 16065 22520 16099
rect 22468 16056 22520 16065
rect 22928 16056 22980 16108
rect 24676 16124 24728 16176
rect 24768 16124 24820 16176
rect 25872 16124 25924 16176
rect 24308 16056 24360 16108
rect 25320 16056 25372 16108
rect 26332 16056 26384 16108
rect 26884 16124 26936 16176
rect 29552 16192 29604 16244
rect 28908 16124 28960 16176
rect 29276 16167 29328 16176
rect 29276 16133 29285 16167
rect 29285 16133 29319 16167
rect 29319 16133 29328 16167
rect 29276 16124 29328 16133
rect 31208 16124 31260 16176
rect 33140 16124 33192 16176
rect 27068 16099 27120 16108
rect 27068 16065 27078 16099
rect 27078 16065 27112 16099
rect 27112 16065 27120 16099
rect 27068 16056 27120 16065
rect 22560 15988 22612 16040
rect 26424 15988 26476 16040
rect 11704 15895 11756 15904
rect 11704 15861 11713 15895
rect 11713 15861 11747 15895
rect 11747 15861 11756 15895
rect 11704 15852 11756 15861
rect 14280 15852 14332 15904
rect 15844 15852 15896 15904
rect 19340 15895 19392 15904
rect 19340 15861 19349 15895
rect 19349 15861 19383 15895
rect 19383 15861 19392 15895
rect 19340 15852 19392 15861
rect 19524 15852 19576 15904
rect 20720 15852 20772 15904
rect 23112 15852 23164 15904
rect 24584 15920 24636 15972
rect 25780 15920 25832 15972
rect 27252 15920 27304 15972
rect 28448 16056 28500 16108
rect 30840 16056 30892 16108
rect 31392 16099 31444 16108
rect 31392 16065 31401 16099
rect 31401 16065 31435 16099
rect 31435 16065 31444 16099
rect 31392 16056 31444 16065
rect 27804 16031 27856 16040
rect 27804 15997 27813 16031
rect 27813 15997 27847 16031
rect 27847 15997 27856 16031
rect 27804 15988 27856 15997
rect 30380 15988 30432 16040
rect 30564 15988 30616 16040
rect 31116 16031 31168 16040
rect 31116 15997 31125 16031
rect 31125 15997 31159 16031
rect 31159 15997 31168 16031
rect 31116 15988 31168 15997
rect 29092 15920 29144 15972
rect 29460 15920 29512 15972
rect 32128 15988 32180 16040
rect 32680 16031 32732 16040
rect 32680 15997 32689 16031
rect 32689 15997 32723 16031
rect 32723 15997 32732 16031
rect 32680 15988 32732 15997
rect 29000 15852 29052 15904
rect 29184 15895 29236 15904
rect 29184 15861 29193 15895
rect 29193 15861 29227 15895
rect 29227 15861 29236 15895
rect 29184 15852 29236 15861
rect 30656 15852 30708 15904
rect 31484 15895 31536 15904
rect 31484 15861 31493 15895
rect 31493 15861 31527 15895
rect 31527 15861 31536 15895
rect 31484 15852 31536 15861
rect 31852 15895 31904 15904
rect 31852 15861 31861 15895
rect 31861 15861 31895 15895
rect 31895 15861 31904 15895
rect 31852 15852 31904 15861
rect 31944 15852 31996 15904
rect 33416 15852 33468 15904
rect 34060 15852 34112 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 6644 15648 6696 15700
rect 7564 15691 7616 15700
rect 7564 15657 7573 15691
rect 7573 15657 7607 15691
rect 7607 15657 7616 15691
rect 7564 15648 7616 15657
rect 7656 15691 7708 15700
rect 7656 15657 7665 15691
rect 7665 15657 7699 15691
rect 7699 15657 7708 15691
rect 7656 15648 7708 15657
rect 8116 15648 8168 15700
rect 5448 15512 5500 15564
rect 2780 15444 2832 15496
rect 2872 15376 2924 15428
rect 3240 15308 3292 15360
rect 5540 15487 5592 15496
rect 5540 15453 5549 15487
rect 5549 15453 5583 15487
rect 5583 15453 5592 15487
rect 5540 15444 5592 15453
rect 6276 15555 6328 15564
rect 6276 15521 6285 15555
rect 6285 15521 6319 15555
rect 6319 15521 6328 15555
rect 6276 15512 6328 15521
rect 4160 15376 4212 15428
rect 5356 15376 5408 15428
rect 4620 15308 4672 15360
rect 5540 15308 5592 15360
rect 5632 15308 5684 15360
rect 7748 15512 7800 15564
rect 7656 15444 7708 15496
rect 9128 15555 9180 15564
rect 9128 15521 9137 15555
rect 9137 15521 9171 15555
rect 9171 15521 9180 15555
rect 9128 15512 9180 15521
rect 9312 15512 9364 15564
rect 12900 15648 12952 15700
rect 15108 15580 15160 15632
rect 16488 15580 16540 15632
rect 18972 15648 19024 15700
rect 20076 15691 20128 15700
rect 20076 15657 20085 15691
rect 20085 15657 20119 15691
rect 20119 15657 20128 15691
rect 20076 15648 20128 15657
rect 22560 15648 22612 15700
rect 23572 15648 23624 15700
rect 24124 15648 24176 15700
rect 24216 15648 24268 15700
rect 26424 15648 26476 15700
rect 26884 15648 26936 15700
rect 28448 15691 28500 15700
rect 28448 15657 28457 15691
rect 28457 15657 28491 15691
rect 28491 15657 28500 15691
rect 28448 15648 28500 15657
rect 30196 15691 30248 15700
rect 30196 15657 30205 15691
rect 30205 15657 30239 15691
rect 30239 15657 30248 15691
rect 30196 15648 30248 15657
rect 31392 15648 31444 15700
rect 19340 15580 19392 15632
rect 22468 15580 22520 15632
rect 13084 15555 13136 15564
rect 13084 15521 13093 15555
rect 13093 15521 13127 15555
rect 13127 15521 13136 15555
rect 13084 15512 13136 15521
rect 13728 15512 13780 15564
rect 6828 15376 6880 15428
rect 7012 15351 7064 15360
rect 7012 15317 7021 15351
rect 7021 15317 7055 15351
rect 7055 15317 7064 15351
rect 7012 15308 7064 15317
rect 7932 15351 7984 15360
rect 7932 15317 7941 15351
rect 7941 15317 7975 15351
rect 7975 15317 7984 15351
rect 7932 15308 7984 15317
rect 9220 15376 9272 15428
rect 9956 15376 10008 15428
rect 11704 15444 11756 15496
rect 12256 15444 12308 15496
rect 15384 15444 15436 15496
rect 15752 15444 15804 15496
rect 15844 15487 15896 15496
rect 15844 15453 15853 15487
rect 15853 15453 15887 15487
rect 15887 15453 15896 15487
rect 15844 15444 15896 15453
rect 16120 15444 16172 15496
rect 17500 15555 17552 15564
rect 17500 15521 17509 15555
rect 17509 15521 17543 15555
rect 17543 15521 17552 15555
rect 17500 15512 17552 15521
rect 20536 15555 20588 15564
rect 20536 15521 20545 15555
rect 20545 15521 20579 15555
rect 20579 15521 20588 15555
rect 20536 15512 20588 15521
rect 20996 15512 21048 15564
rect 22928 15512 22980 15564
rect 23940 15555 23992 15564
rect 23940 15521 23949 15555
rect 23949 15521 23983 15555
rect 23983 15521 23992 15555
rect 23940 15512 23992 15521
rect 24032 15512 24084 15564
rect 26516 15580 26568 15632
rect 24400 15512 24452 15564
rect 26792 15512 26844 15564
rect 27252 15512 27304 15564
rect 27436 15512 27488 15564
rect 29092 15555 29144 15564
rect 29092 15521 29101 15555
rect 29101 15521 29135 15555
rect 29135 15521 29144 15555
rect 29092 15512 29144 15521
rect 18052 15444 18104 15496
rect 19064 15444 19116 15496
rect 9036 15351 9088 15360
rect 9036 15317 9045 15351
rect 9045 15317 9079 15351
rect 9079 15317 9088 15351
rect 9036 15308 9088 15317
rect 10784 15351 10836 15360
rect 10784 15317 10793 15351
rect 10793 15317 10827 15351
rect 10827 15317 10836 15351
rect 10784 15308 10836 15317
rect 11520 15351 11572 15360
rect 11520 15317 11529 15351
rect 11529 15317 11563 15351
rect 11563 15317 11572 15351
rect 11520 15308 11572 15317
rect 12624 15376 12676 15428
rect 14740 15376 14792 15428
rect 17960 15376 18012 15428
rect 19432 15444 19484 15496
rect 21364 15444 21416 15496
rect 24676 15444 24728 15496
rect 27804 15444 27856 15496
rect 30380 15487 30432 15496
rect 30380 15453 30389 15487
rect 30389 15453 30423 15487
rect 30423 15453 30432 15487
rect 30380 15444 30432 15453
rect 12440 15308 12492 15360
rect 12900 15308 12952 15360
rect 16396 15351 16448 15360
rect 16396 15317 16405 15351
rect 16405 15317 16439 15351
rect 16439 15317 16448 15351
rect 16396 15308 16448 15317
rect 20720 15376 20772 15428
rect 21824 15376 21876 15428
rect 23940 15376 23992 15428
rect 25320 15376 25372 15428
rect 26056 15376 26108 15428
rect 29184 15376 29236 15428
rect 30656 15487 30708 15496
rect 30656 15453 30690 15487
rect 30690 15453 30708 15487
rect 30656 15444 30708 15453
rect 30840 15376 30892 15428
rect 31208 15376 31260 15428
rect 33048 15419 33100 15428
rect 33048 15385 33057 15419
rect 33057 15385 33091 15419
rect 33091 15385 33100 15419
rect 34796 15444 34848 15496
rect 33048 15376 33100 15385
rect 34704 15376 34756 15428
rect 20812 15308 20864 15360
rect 20996 15351 21048 15360
rect 20996 15317 21005 15351
rect 21005 15317 21039 15351
rect 21039 15317 21048 15351
rect 20996 15308 21048 15317
rect 21916 15308 21968 15360
rect 24124 15308 24176 15360
rect 24768 15308 24820 15360
rect 25504 15308 25556 15360
rect 29276 15351 29328 15360
rect 29276 15317 29285 15351
rect 29285 15317 29319 15351
rect 29319 15317 29328 15351
rect 29276 15308 29328 15317
rect 30380 15308 30432 15360
rect 30564 15308 30616 15360
rect 31484 15308 31536 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 2872 15147 2924 15156
rect 2872 15113 2881 15147
rect 2881 15113 2915 15147
rect 2915 15113 2924 15147
rect 2872 15104 2924 15113
rect 3240 15147 3292 15156
rect 3240 15113 3249 15147
rect 3249 15113 3283 15147
rect 3283 15113 3292 15147
rect 3240 15104 3292 15113
rect 3700 15147 3752 15156
rect 3700 15113 3709 15147
rect 3709 15113 3743 15147
rect 3743 15113 3752 15147
rect 3700 15104 3752 15113
rect 4160 15147 4212 15156
rect 4160 15113 4169 15147
rect 4169 15113 4203 15147
rect 4203 15113 4212 15147
rect 4160 15104 4212 15113
rect 4620 15147 4672 15156
rect 4620 15113 4629 15147
rect 4629 15113 4663 15147
rect 4663 15113 4672 15147
rect 4620 15104 4672 15113
rect 9220 15104 9272 15156
rect 9956 15147 10008 15156
rect 9956 15113 9965 15147
rect 9965 15113 9999 15147
rect 9999 15113 10008 15147
rect 9956 15104 10008 15113
rect 10784 15104 10836 15156
rect 4068 15036 4120 15088
rect 1308 14968 1360 15020
rect 9312 15036 9364 15088
rect 10876 15036 10928 15088
rect 11336 15036 11388 15088
rect 7932 14968 7984 15020
rect 8024 14968 8076 15020
rect 3700 14900 3752 14952
rect 5356 14900 5408 14952
rect 11244 14968 11296 15020
rect 12624 15104 12676 15156
rect 12808 15104 12860 15156
rect 14924 15104 14976 15156
rect 15660 15104 15712 15156
rect 16212 15104 16264 15156
rect 17960 15147 18012 15156
rect 17960 15113 17969 15147
rect 17969 15113 18003 15147
rect 18003 15113 18012 15147
rect 17960 15104 18012 15113
rect 18972 15104 19024 15156
rect 16396 15036 16448 15088
rect 20536 15104 20588 15156
rect 20720 15104 20772 15156
rect 21456 15147 21508 15156
rect 21456 15113 21465 15147
rect 21465 15113 21499 15147
rect 21499 15113 21508 15147
rect 21456 15104 21508 15113
rect 21824 15147 21876 15156
rect 21824 15113 21833 15147
rect 21833 15113 21867 15147
rect 21867 15113 21876 15147
rect 21824 15104 21876 15113
rect 22560 15104 22612 15156
rect 23572 15147 23624 15156
rect 23572 15113 23581 15147
rect 23581 15113 23615 15147
rect 23615 15113 23624 15147
rect 23572 15104 23624 15113
rect 24032 15104 24084 15156
rect 24216 15104 24268 15156
rect 26240 15104 26292 15156
rect 27068 15104 27120 15156
rect 29736 15147 29788 15156
rect 29736 15113 29745 15147
rect 29745 15113 29779 15147
rect 29779 15113 29788 15147
rect 29736 15104 29788 15113
rect 30012 15147 30064 15156
rect 30012 15113 30021 15147
rect 30021 15113 30055 15147
rect 30055 15113 30064 15147
rect 30012 15104 30064 15113
rect 30564 15147 30616 15156
rect 30564 15113 30573 15147
rect 30573 15113 30607 15147
rect 30607 15113 30616 15147
rect 30564 15104 30616 15113
rect 30932 15104 30984 15156
rect 14648 14968 14700 15020
rect 11428 14900 11480 14952
rect 12624 14943 12676 14952
rect 12624 14909 12633 14943
rect 12633 14909 12667 14943
rect 12667 14909 12676 14943
rect 12624 14900 12676 14909
rect 12808 14943 12860 14952
rect 12808 14909 12817 14943
rect 12817 14909 12851 14943
rect 12851 14909 12860 14943
rect 12808 14900 12860 14909
rect 3700 14764 3752 14816
rect 4804 14764 4856 14816
rect 5356 14764 5408 14816
rect 5448 14764 5500 14816
rect 6368 14764 6420 14816
rect 11244 14807 11296 14816
rect 11244 14773 11253 14807
rect 11253 14773 11287 14807
rect 11287 14773 11296 14807
rect 11244 14764 11296 14773
rect 11520 14807 11572 14816
rect 11520 14773 11529 14807
rect 11529 14773 11563 14807
rect 11563 14773 11572 14807
rect 11520 14764 11572 14773
rect 13728 14832 13780 14884
rect 14004 14764 14056 14816
rect 16120 14900 16172 14952
rect 17776 14832 17828 14884
rect 19524 14968 19576 15020
rect 20904 15011 20956 15020
rect 20904 14977 20914 15011
rect 20914 14977 20948 15011
rect 20948 14977 20956 15011
rect 20904 14968 20956 14977
rect 21088 15011 21140 15020
rect 21088 14977 21097 15011
rect 21097 14977 21131 15011
rect 21131 14977 21140 15011
rect 21088 14968 21140 14977
rect 21732 14968 21784 15020
rect 20536 14943 20588 14952
rect 20536 14909 20545 14943
rect 20545 14909 20579 14943
rect 20579 14909 20588 14943
rect 20536 14900 20588 14909
rect 22652 14968 22704 15020
rect 23480 14968 23532 15020
rect 24124 14968 24176 15020
rect 24216 15011 24268 15020
rect 24216 14977 24225 15011
rect 24225 14977 24259 15011
rect 24259 14977 24268 15011
rect 24216 14968 24268 14977
rect 24676 15011 24728 15020
rect 24676 14977 24685 15011
rect 24685 14977 24719 15011
rect 24719 14977 24728 15011
rect 24676 14968 24728 14977
rect 25228 14968 25280 15020
rect 26884 14968 26936 15020
rect 27068 14968 27120 15020
rect 22468 14943 22520 14952
rect 22468 14909 22477 14943
rect 22477 14909 22511 14943
rect 22511 14909 22520 14943
rect 22468 14900 22520 14909
rect 26976 14943 27028 14952
rect 26976 14909 26985 14943
rect 26985 14909 27019 14943
rect 27019 14909 27028 14943
rect 26976 14900 27028 14909
rect 28908 15036 28960 15088
rect 28540 14968 28592 15020
rect 28724 14968 28776 15020
rect 29920 15079 29972 15088
rect 29920 15045 29929 15079
rect 29929 15045 29963 15079
rect 29963 15045 29972 15079
rect 29920 15036 29972 15045
rect 30472 15079 30524 15088
rect 30472 15045 30481 15079
rect 30481 15045 30515 15079
rect 30515 15045 30524 15079
rect 30472 15036 30524 15045
rect 29184 15011 29236 15020
rect 29184 14977 29194 15011
rect 29194 14977 29228 15011
rect 29228 14977 29236 15011
rect 29184 14968 29236 14977
rect 29368 15011 29420 15020
rect 29368 14977 29377 15011
rect 29377 14977 29411 15011
rect 29411 14977 29420 15011
rect 29368 14968 29420 14977
rect 29460 15011 29512 15020
rect 29460 14977 29469 15011
rect 29469 14977 29503 15011
rect 29503 14977 29512 15011
rect 29460 14968 29512 14977
rect 29552 14968 29604 15020
rect 30196 14968 30248 15020
rect 31024 15036 31076 15088
rect 32680 15147 32732 15156
rect 32680 15113 32689 15147
rect 32689 15113 32723 15147
rect 32723 15113 32732 15147
rect 32680 15104 32732 15113
rect 33140 15104 33192 15156
rect 33416 15036 33468 15088
rect 31852 14968 31904 15020
rect 32588 14968 32640 15020
rect 15108 14764 15160 14816
rect 15752 14764 15804 14816
rect 16488 14807 16540 14816
rect 16488 14773 16497 14807
rect 16497 14773 16531 14807
rect 16531 14773 16540 14807
rect 16488 14764 16540 14773
rect 16764 14764 16816 14816
rect 17592 14807 17644 14816
rect 17592 14773 17601 14807
rect 17601 14773 17635 14807
rect 17635 14773 17644 14807
rect 17592 14764 17644 14773
rect 19984 14807 20036 14816
rect 19984 14773 19993 14807
rect 19993 14773 20027 14807
rect 20027 14773 20036 14807
rect 19984 14764 20036 14773
rect 20536 14764 20588 14816
rect 24032 14832 24084 14884
rect 28172 14832 28224 14884
rect 28632 14875 28684 14884
rect 28632 14841 28641 14875
rect 28641 14841 28675 14875
rect 28675 14841 28684 14875
rect 28632 14832 28684 14841
rect 29368 14832 29420 14884
rect 32036 14832 32088 14884
rect 32128 14832 32180 14884
rect 33048 14832 33100 14884
rect 33968 14900 34020 14952
rect 22468 14764 22520 14816
rect 23204 14764 23256 14816
rect 26332 14807 26384 14816
rect 26332 14773 26341 14807
rect 26341 14773 26375 14807
rect 26375 14773 26384 14807
rect 26516 14807 26568 14816
rect 26332 14764 26384 14773
rect 26516 14773 26525 14807
rect 26525 14773 26559 14807
rect 26559 14773 26568 14807
rect 26516 14764 26568 14773
rect 27988 14764 28040 14816
rect 28448 14764 28500 14816
rect 28724 14764 28776 14816
rect 30012 14764 30064 14816
rect 31484 14764 31536 14816
rect 34796 14764 34848 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3424 14560 3476 14612
rect 6368 14492 6420 14544
rect 11980 14492 12032 14544
rect 12164 14560 12216 14612
rect 14648 14603 14700 14612
rect 14648 14569 14657 14603
rect 14657 14569 14691 14603
rect 14691 14569 14700 14603
rect 14648 14560 14700 14569
rect 10416 14467 10468 14476
rect 10416 14433 10425 14467
rect 10425 14433 10459 14467
rect 10459 14433 10468 14467
rect 10416 14424 10468 14433
rect 11060 14424 11112 14476
rect 12256 14424 12308 14476
rect 12716 14424 12768 14476
rect 15016 14492 15068 14544
rect 16120 14560 16172 14612
rect 16396 14560 16448 14612
rect 20904 14560 20956 14612
rect 21732 14560 21784 14612
rect 22008 14560 22060 14612
rect 24492 14560 24544 14612
rect 25228 14603 25280 14612
rect 25228 14569 25237 14603
rect 25237 14569 25271 14603
rect 25271 14569 25280 14603
rect 25228 14560 25280 14569
rect 26148 14560 26200 14612
rect 27068 14560 27120 14612
rect 27896 14603 27948 14612
rect 27896 14569 27905 14603
rect 27905 14569 27939 14603
rect 27939 14569 27948 14603
rect 27896 14560 27948 14569
rect 14556 14424 14608 14476
rect 7748 14356 7800 14408
rect 6368 14288 6420 14340
rect 9496 14288 9548 14340
rect 5540 14220 5592 14272
rect 6736 14263 6788 14272
rect 6736 14229 6745 14263
rect 6745 14229 6779 14263
rect 6779 14229 6788 14263
rect 6736 14220 6788 14229
rect 9864 14263 9916 14272
rect 9864 14229 9873 14263
rect 9873 14229 9907 14263
rect 9907 14229 9916 14263
rect 9864 14220 9916 14229
rect 10692 14288 10744 14340
rect 10784 14220 10836 14272
rect 11152 14331 11204 14340
rect 11152 14297 11161 14331
rect 11161 14297 11195 14331
rect 11195 14297 11204 14331
rect 11152 14288 11204 14297
rect 11980 14356 12032 14408
rect 12256 14220 12308 14272
rect 12348 14220 12400 14272
rect 15660 14356 15712 14408
rect 22468 14492 22520 14544
rect 17500 14424 17552 14476
rect 16764 14399 16816 14408
rect 16764 14365 16782 14399
rect 16782 14365 16816 14399
rect 16764 14356 16816 14365
rect 19432 14399 19484 14408
rect 19432 14365 19441 14399
rect 19441 14365 19475 14399
rect 19475 14365 19484 14399
rect 19432 14356 19484 14365
rect 19984 14356 20036 14408
rect 22376 14356 22428 14408
rect 24768 14492 24820 14544
rect 24584 14424 24636 14476
rect 26148 14424 26200 14476
rect 27436 14467 27488 14476
rect 27436 14433 27445 14467
rect 27445 14433 27479 14467
rect 27479 14433 27488 14467
rect 27436 14424 27488 14433
rect 24676 14356 24728 14408
rect 26240 14356 26292 14408
rect 27988 14399 28040 14408
rect 27988 14365 27997 14399
rect 27997 14365 28031 14399
rect 28031 14365 28040 14399
rect 27988 14356 28040 14365
rect 13084 14220 13136 14272
rect 20904 14288 20956 14340
rect 16672 14220 16724 14272
rect 20628 14220 20680 14272
rect 21088 14220 21140 14272
rect 24124 14220 24176 14272
rect 24492 14220 24544 14272
rect 24952 14220 25004 14272
rect 25688 14220 25740 14272
rect 26148 14263 26200 14272
rect 26148 14229 26157 14263
rect 26157 14229 26191 14263
rect 26191 14229 26200 14263
rect 26148 14220 26200 14229
rect 27988 14220 28040 14272
rect 28264 14424 28316 14476
rect 32036 14560 32088 14612
rect 28172 14331 28224 14340
rect 28172 14297 28181 14331
rect 28181 14297 28215 14331
rect 28215 14297 28224 14331
rect 28172 14288 28224 14297
rect 28264 14331 28316 14340
rect 28264 14297 28273 14331
rect 28273 14297 28307 14331
rect 28307 14297 28316 14331
rect 28264 14288 28316 14297
rect 28632 14492 28684 14544
rect 29276 14492 29328 14544
rect 28724 14424 28776 14476
rect 30288 14424 30340 14476
rect 30840 14492 30892 14544
rect 30564 14467 30616 14476
rect 30564 14433 30573 14467
rect 30573 14433 30607 14467
rect 30607 14433 30616 14467
rect 30564 14424 30616 14433
rect 28632 14399 28684 14408
rect 28632 14365 28647 14399
rect 28647 14365 28681 14399
rect 28681 14365 28684 14399
rect 28632 14356 28684 14365
rect 28816 14356 28868 14408
rect 29276 14356 29328 14408
rect 29460 14356 29512 14408
rect 31116 14356 31168 14408
rect 33968 14603 34020 14612
rect 33968 14569 33977 14603
rect 33977 14569 34011 14603
rect 34011 14569 34020 14603
rect 33968 14560 34020 14569
rect 34428 14399 34480 14408
rect 34428 14365 34437 14399
rect 34437 14365 34471 14399
rect 34471 14365 34480 14399
rect 34428 14356 34480 14365
rect 28908 14288 28960 14340
rect 34796 14288 34848 14340
rect 28724 14220 28776 14272
rect 28816 14263 28868 14272
rect 28816 14229 28825 14263
rect 28825 14229 28859 14263
rect 28859 14229 28868 14263
rect 28816 14220 28868 14229
rect 30012 14263 30064 14272
rect 30012 14229 30021 14263
rect 30021 14229 30055 14263
rect 30055 14229 30064 14263
rect 30012 14220 30064 14229
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 6276 14016 6328 14068
rect 6368 14059 6420 14068
rect 6368 14025 6377 14059
rect 6377 14025 6411 14059
rect 6411 14025 6420 14059
rect 6368 14016 6420 14025
rect 6736 14059 6788 14068
rect 6736 14025 6745 14059
rect 6745 14025 6779 14059
rect 6779 14025 6788 14059
rect 6736 14016 6788 14025
rect 7748 14059 7800 14068
rect 7748 14025 7757 14059
rect 7757 14025 7791 14059
rect 7791 14025 7800 14059
rect 7748 14016 7800 14025
rect 5448 13948 5500 14000
rect 2872 13880 2924 13932
rect 3424 13923 3476 13932
rect 3424 13889 3433 13923
rect 3433 13889 3467 13923
rect 3467 13889 3476 13923
rect 3424 13880 3476 13889
rect 4160 13880 4212 13932
rect 4620 13923 4672 13932
rect 4620 13889 4629 13923
rect 4629 13889 4663 13923
rect 4663 13889 4672 13923
rect 4620 13880 4672 13889
rect 5264 13880 5316 13932
rect 6920 13948 6972 14000
rect 7656 13948 7708 14000
rect 8392 14016 8444 14068
rect 8760 14016 8812 14068
rect 10692 14059 10744 14068
rect 10692 14025 10701 14059
rect 10701 14025 10735 14059
rect 10735 14025 10744 14059
rect 10692 14016 10744 14025
rect 11152 14016 11204 14068
rect 11888 14016 11940 14068
rect 13268 14016 13320 14068
rect 14556 14016 14608 14068
rect 16580 14016 16632 14068
rect 9864 13948 9916 14000
rect 10416 13948 10468 14000
rect 14004 13948 14056 14000
rect 7012 13855 7064 13864
rect 7012 13821 7021 13855
rect 7021 13821 7055 13855
rect 7055 13821 7064 13855
rect 7012 13812 7064 13821
rect 9312 13923 9364 13932
rect 9312 13889 9321 13923
rect 9321 13889 9355 13923
rect 9355 13889 9364 13923
rect 9312 13880 9364 13889
rect 11980 13880 12032 13932
rect 12440 13880 12492 13932
rect 12624 13923 12676 13932
rect 12624 13889 12658 13923
rect 12658 13889 12676 13923
rect 12624 13880 12676 13889
rect 12992 13880 13044 13932
rect 7656 13812 7708 13864
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 14188 13923 14240 13932
rect 14188 13889 14197 13923
rect 14197 13889 14231 13923
rect 14231 13889 14240 13923
rect 14188 13880 14240 13889
rect 14280 13880 14332 13932
rect 14648 13855 14700 13864
rect 3700 13676 3752 13728
rect 6828 13676 6880 13728
rect 9496 13676 9548 13728
rect 11520 13719 11572 13728
rect 11520 13685 11529 13719
rect 11529 13685 11563 13719
rect 11563 13685 11572 13719
rect 11520 13676 11572 13685
rect 14648 13821 14657 13855
rect 14657 13821 14691 13855
rect 14691 13821 14700 13855
rect 14648 13812 14700 13821
rect 15108 13880 15160 13932
rect 17316 13880 17368 13932
rect 17500 13880 17552 13932
rect 19156 13880 19208 13932
rect 24124 14016 24176 14068
rect 24860 14016 24912 14068
rect 26424 14016 26476 14068
rect 27068 14059 27120 14068
rect 27068 14025 27077 14059
rect 27077 14025 27111 14059
rect 27111 14025 27120 14059
rect 27068 14016 27120 14025
rect 27896 14016 27948 14068
rect 28264 14016 28316 14068
rect 28816 14016 28868 14068
rect 31116 14059 31168 14068
rect 31116 14025 31125 14059
rect 31125 14025 31159 14059
rect 31159 14025 31168 14059
rect 31116 14016 31168 14025
rect 22284 13880 22336 13932
rect 15016 13812 15068 13864
rect 22376 13855 22428 13864
rect 22376 13821 22385 13855
rect 22385 13821 22419 13855
rect 22419 13821 22428 13855
rect 22376 13812 22428 13821
rect 25412 13948 25464 14000
rect 26148 13948 26200 14000
rect 28448 13991 28500 14000
rect 28448 13957 28482 13991
rect 28482 13957 28500 13991
rect 28448 13948 28500 13957
rect 24676 13923 24728 13932
rect 24676 13889 24685 13923
rect 24685 13889 24719 13923
rect 24719 13889 24728 13923
rect 24676 13880 24728 13889
rect 24860 13923 24912 13932
rect 24860 13889 24869 13923
rect 24869 13889 24903 13923
rect 24903 13889 24912 13923
rect 24860 13880 24912 13889
rect 12716 13676 12768 13728
rect 13544 13676 13596 13728
rect 13728 13719 13780 13728
rect 13728 13685 13737 13719
rect 13737 13685 13771 13719
rect 13771 13685 13780 13719
rect 13728 13676 13780 13685
rect 16488 13676 16540 13728
rect 17960 13676 18012 13728
rect 21732 13744 21784 13796
rect 18696 13676 18748 13728
rect 19708 13719 19760 13728
rect 19708 13685 19717 13719
rect 19717 13685 19751 13719
rect 19751 13685 19760 13719
rect 19708 13676 19760 13685
rect 22100 13676 22152 13728
rect 24400 13855 24452 13864
rect 24400 13821 24409 13855
rect 24409 13821 24443 13855
rect 24443 13821 24452 13855
rect 24400 13812 24452 13821
rect 24768 13812 24820 13864
rect 26056 13880 26108 13932
rect 26976 13880 27028 13932
rect 27804 13880 27856 13932
rect 27252 13812 27304 13864
rect 29552 13880 29604 13932
rect 32128 13948 32180 14000
rect 30012 13923 30064 13932
rect 30012 13889 30046 13923
rect 30046 13889 30064 13923
rect 30012 13880 30064 13889
rect 29736 13855 29788 13864
rect 29736 13821 29745 13855
rect 29745 13821 29779 13855
rect 29779 13821 29788 13855
rect 29736 13812 29788 13821
rect 26516 13744 26568 13796
rect 25688 13719 25740 13728
rect 25688 13685 25697 13719
rect 25697 13685 25731 13719
rect 25731 13685 25740 13719
rect 25688 13676 25740 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 4068 13472 4120 13524
rect 6920 13515 6972 13524
rect 6920 13481 6929 13515
rect 6929 13481 6963 13515
rect 6963 13481 6972 13515
rect 6920 13472 6972 13481
rect 7012 13472 7064 13524
rect 11888 13515 11940 13524
rect 11888 13481 11897 13515
rect 11897 13481 11931 13515
rect 11931 13481 11940 13515
rect 11888 13472 11940 13481
rect 12256 13515 12308 13524
rect 12256 13481 12265 13515
rect 12265 13481 12299 13515
rect 12299 13481 12308 13515
rect 12256 13472 12308 13481
rect 12624 13472 12676 13524
rect 14924 13515 14976 13524
rect 14924 13481 14933 13515
rect 14933 13481 14967 13515
rect 14967 13481 14976 13515
rect 14924 13472 14976 13481
rect 17316 13515 17368 13524
rect 17316 13481 17325 13515
rect 17325 13481 17359 13515
rect 17359 13481 17368 13515
rect 17316 13472 17368 13481
rect 19156 13472 19208 13524
rect 12716 13404 12768 13456
rect 13176 13404 13228 13456
rect 13636 13447 13688 13456
rect 5540 13379 5592 13388
rect 5540 13345 5549 13379
rect 5549 13345 5583 13379
rect 5583 13345 5592 13379
rect 5540 13336 5592 13345
rect 9128 13336 9180 13388
rect 9588 13336 9640 13388
rect 13268 13336 13320 13388
rect 13636 13413 13645 13447
rect 13645 13413 13679 13447
rect 13679 13413 13688 13447
rect 13636 13404 13688 13413
rect 14188 13336 14240 13388
rect 14832 13336 14884 13388
rect 17592 13404 17644 13456
rect 15108 13379 15160 13388
rect 15108 13345 15117 13379
rect 15117 13345 15151 13379
rect 15151 13345 15160 13379
rect 15108 13336 15160 13345
rect 18512 13404 18564 13456
rect 22192 13404 22244 13456
rect 24400 13472 24452 13524
rect 24584 13472 24636 13524
rect 26332 13472 26384 13524
rect 27252 13515 27304 13524
rect 27252 13481 27261 13515
rect 27261 13481 27295 13515
rect 27295 13481 27304 13515
rect 27252 13472 27304 13481
rect 27528 13515 27580 13524
rect 27528 13481 27537 13515
rect 27537 13481 27571 13515
rect 27571 13481 27580 13515
rect 27528 13472 27580 13481
rect 2780 13268 2832 13320
rect 9312 13268 9364 13320
rect 11520 13268 11572 13320
rect 12256 13311 12308 13320
rect 12256 13277 12265 13311
rect 12265 13277 12299 13311
rect 12299 13277 12308 13311
rect 12256 13268 12308 13277
rect 13728 13268 13780 13320
rect 2964 13200 3016 13252
rect 4068 13243 4120 13252
rect 4068 13209 4102 13243
rect 4102 13209 4120 13243
rect 4068 13200 4120 13209
rect 6368 13200 6420 13252
rect 4344 13132 4396 13184
rect 4620 13132 4672 13184
rect 8852 13132 8904 13184
rect 9496 13200 9548 13252
rect 11980 13200 12032 13252
rect 12440 13200 12492 13252
rect 9036 13132 9088 13184
rect 12624 13175 12676 13184
rect 12624 13141 12633 13175
rect 12633 13141 12667 13175
rect 12667 13141 12676 13175
rect 12624 13132 12676 13141
rect 12900 13132 12952 13184
rect 13176 13132 13228 13184
rect 14096 13175 14148 13184
rect 14096 13141 14105 13175
rect 14105 13141 14139 13175
rect 14139 13141 14148 13175
rect 14096 13132 14148 13141
rect 16580 13311 16632 13320
rect 16580 13277 16589 13311
rect 16589 13277 16623 13311
rect 16623 13277 16632 13311
rect 16580 13268 16632 13277
rect 17960 13268 18012 13320
rect 19616 13336 19668 13388
rect 22376 13336 22428 13388
rect 15660 13200 15712 13252
rect 19432 13268 19484 13320
rect 20996 13268 21048 13320
rect 23848 13268 23900 13320
rect 26424 13311 26476 13320
rect 26424 13277 26433 13311
rect 26433 13277 26467 13311
rect 26467 13277 26476 13311
rect 26424 13268 26476 13277
rect 26884 13404 26936 13456
rect 28448 13515 28500 13524
rect 28448 13481 28457 13515
rect 28457 13481 28491 13515
rect 28491 13481 28500 13515
rect 28448 13472 28500 13481
rect 29276 13515 29328 13524
rect 29276 13481 29285 13515
rect 29285 13481 29319 13515
rect 29319 13481 29328 13515
rect 29276 13472 29328 13481
rect 30564 13404 30616 13456
rect 28080 13336 28132 13388
rect 16028 13132 16080 13184
rect 16764 13175 16816 13184
rect 16764 13141 16773 13175
rect 16773 13141 16807 13175
rect 16807 13141 16816 13175
rect 16764 13132 16816 13141
rect 17500 13132 17552 13184
rect 20536 13200 20588 13252
rect 21824 13200 21876 13252
rect 19708 13175 19760 13184
rect 19708 13141 19717 13175
rect 19717 13141 19751 13175
rect 19751 13141 19760 13175
rect 19708 13132 19760 13141
rect 25504 13200 25556 13252
rect 27252 13268 27304 13320
rect 27344 13311 27396 13320
rect 27344 13277 27353 13311
rect 27353 13277 27387 13311
rect 27387 13277 27396 13311
rect 27344 13268 27396 13277
rect 27896 13268 27948 13320
rect 28816 13311 28868 13320
rect 28816 13277 28825 13311
rect 28825 13277 28859 13311
rect 28859 13277 28868 13311
rect 28816 13268 28868 13277
rect 27804 13200 27856 13252
rect 28632 13200 28684 13252
rect 22836 13132 22888 13184
rect 23388 13132 23440 13184
rect 24124 13132 24176 13184
rect 26332 13175 26384 13184
rect 26332 13141 26341 13175
rect 26341 13141 26375 13175
rect 26375 13141 26384 13175
rect 26332 13132 26384 13141
rect 26608 13132 26660 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 2872 12928 2924 12980
rect 2964 12971 3016 12980
rect 2964 12937 2973 12971
rect 2973 12937 3007 12971
rect 3007 12937 3016 12971
rect 2964 12928 3016 12937
rect 4068 12928 4120 12980
rect 4344 12971 4396 12980
rect 4344 12937 4353 12971
rect 4353 12937 4387 12971
rect 4387 12937 4396 12971
rect 4344 12928 4396 12937
rect 6368 12971 6420 12980
rect 6368 12937 6377 12971
rect 6377 12937 6411 12971
rect 6411 12937 6420 12971
rect 6368 12928 6420 12937
rect 6920 12928 6972 12980
rect 12256 12928 12308 12980
rect 14188 12928 14240 12980
rect 15660 12971 15712 12980
rect 15660 12937 15669 12971
rect 15669 12937 15703 12971
rect 15703 12937 15712 12971
rect 15660 12928 15712 12937
rect 16028 12971 16080 12980
rect 16028 12937 16037 12971
rect 16037 12937 16071 12971
rect 16071 12937 16080 12971
rect 16028 12928 16080 12937
rect 16764 12928 16816 12980
rect 4160 12860 4212 12912
rect 6276 12860 6328 12912
rect 9404 12903 9456 12912
rect 1308 12792 1360 12844
rect 3700 12792 3752 12844
rect 6828 12835 6880 12844
rect 6828 12801 6837 12835
rect 6837 12801 6871 12835
rect 6871 12801 6880 12835
rect 6828 12792 6880 12801
rect 4712 12724 4764 12776
rect 5264 12724 5316 12776
rect 7196 12767 7248 12776
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 8208 12724 8260 12776
rect 8852 12792 8904 12844
rect 9404 12869 9413 12903
rect 9413 12869 9447 12903
rect 9447 12869 9456 12903
rect 9404 12860 9456 12869
rect 11152 12860 11204 12912
rect 14096 12860 14148 12912
rect 9680 12792 9732 12844
rect 10048 12792 10100 12844
rect 16948 12860 17000 12912
rect 24768 12928 24820 12980
rect 25504 12971 25556 12980
rect 25504 12937 25513 12971
rect 25513 12937 25547 12971
rect 25547 12937 25556 12971
rect 25504 12928 25556 12937
rect 26332 12928 26384 12980
rect 26884 12928 26936 12980
rect 27804 12928 27856 12980
rect 17960 12860 18012 12912
rect 12532 12724 12584 12776
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 6460 12656 6512 12708
rect 16580 12724 16632 12776
rect 17592 12792 17644 12844
rect 5356 12588 5408 12640
rect 12716 12588 12768 12640
rect 15936 12588 15988 12640
rect 16856 12588 16908 12640
rect 20996 12860 21048 12912
rect 18420 12835 18472 12844
rect 18420 12801 18429 12835
rect 18429 12801 18463 12835
rect 18463 12801 18472 12835
rect 18420 12792 18472 12801
rect 18512 12835 18564 12844
rect 18512 12801 18526 12835
rect 18526 12801 18560 12835
rect 18560 12801 18564 12835
rect 18512 12792 18564 12801
rect 18788 12835 18840 12844
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 18788 12792 18840 12801
rect 19064 12835 19116 12844
rect 19064 12801 19073 12835
rect 19073 12801 19107 12835
rect 19107 12801 19116 12835
rect 19064 12792 19116 12801
rect 19156 12835 19208 12844
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 19708 12792 19760 12844
rect 20904 12835 20956 12844
rect 20904 12801 20913 12835
rect 20913 12801 20947 12835
rect 20947 12801 20956 12835
rect 20904 12792 20956 12801
rect 21088 12835 21140 12844
rect 21088 12801 21097 12835
rect 21097 12801 21131 12835
rect 21131 12801 21140 12835
rect 21088 12792 21140 12801
rect 19248 12724 19300 12776
rect 22192 12860 22244 12912
rect 18788 12656 18840 12708
rect 20628 12656 20680 12708
rect 20812 12656 20864 12708
rect 21732 12792 21784 12844
rect 19524 12631 19576 12640
rect 19524 12597 19533 12631
rect 19533 12597 19567 12631
rect 19567 12597 19576 12631
rect 19524 12588 19576 12597
rect 19708 12588 19760 12640
rect 23296 12835 23348 12844
rect 23296 12801 23306 12835
rect 23306 12801 23340 12835
rect 23340 12801 23348 12835
rect 23296 12792 23348 12801
rect 23388 12792 23440 12844
rect 23572 12835 23624 12844
rect 23572 12801 23581 12835
rect 23581 12801 23615 12835
rect 23615 12801 23624 12835
rect 23572 12792 23624 12801
rect 23664 12835 23716 12844
rect 24676 12860 24728 12912
rect 26700 12860 26752 12912
rect 27344 12860 27396 12912
rect 33140 12860 33192 12912
rect 23664 12801 23678 12835
rect 23678 12801 23712 12835
rect 23712 12801 23716 12835
rect 23664 12792 23716 12801
rect 26516 12835 26568 12844
rect 26516 12801 26525 12835
rect 26525 12801 26559 12835
rect 26559 12801 26568 12835
rect 26516 12792 26568 12801
rect 26976 12835 27028 12844
rect 26976 12801 26985 12835
rect 26985 12801 27019 12835
rect 27019 12801 27028 12835
rect 26976 12792 27028 12801
rect 27252 12835 27304 12844
rect 27252 12801 27286 12835
rect 27286 12801 27304 12835
rect 27252 12792 27304 12801
rect 32128 12835 32180 12844
rect 32128 12801 32137 12835
rect 32137 12801 32171 12835
rect 32171 12801 32180 12835
rect 32128 12792 32180 12801
rect 33876 12792 33928 12844
rect 22560 12724 22612 12776
rect 25228 12724 25280 12776
rect 22744 12656 22796 12708
rect 24952 12656 25004 12708
rect 26148 12767 26200 12776
rect 26148 12733 26157 12767
rect 26157 12733 26191 12767
rect 26191 12733 26200 12767
rect 26148 12724 26200 12733
rect 32404 12767 32456 12776
rect 32404 12733 32413 12767
rect 32413 12733 32447 12767
rect 32447 12733 32456 12767
rect 32404 12724 32456 12733
rect 35348 12724 35400 12776
rect 26424 12656 26476 12708
rect 24860 12631 24912 12640
rect 24860 12597 24869 12631
rect 24869 12597 24903 12631
rect 24903 12597 24912 12631
rect 24860 12588 24912 12597
rect 25596 12588 25648 12640
rect 28632 12631 28684 12640
rect 28632 12597 28641 12631
rect 28641 12597 28675 12631
rect 28675 12597 28684 12631
rect 28632 12588 28684 12597
rect 33876 12631 33928 12640
rect 33876 12597 33885 12631
rect 33885 12597 33919 12631
rect 33919 12597 33928 12631
rect 33876 12588 33928 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 12992 12427 13044 12436
rect 12992 12393 13001 12427
rect 13001 12393 13035 12427
rect 13035 12393 13044 12427
rect 12992 12384 13044 12393
rect 13912 12384 13964 12436
rect 16304 12384 16356 12436
rect 20996 12384 21048 12436
rect 21088 12384 21140 12436
rect 21824 12427 21876 12436
rect 21824 12393 21833 12427
rect 21833 12393 21867 12427
rect 21867 12393 21876 12427
rect 21824 12384 21876 12393
rect 22100 12384 22152 12436
rect 22744 12384 22796 12436
rect 23572 12384 23624 12436
rect 25780 12427 25832 12436
rect 25780 12393 25789 12427
rect 25789 12393 25823 12427
rect 25823 12393 25832 12427
rect 25780 12384 25832 12393
rect 26608 12427 26660 12436
rect 26608 12393 26617 12427
rect 26617 12393 26651 12427
rect 26651 12393 26660 12427
rect 26608 12384 26660 12393
rect 27068 12384 27120 12436
rect 27252 12427 27304 12436
rect 27252 12393 27261 12427
rect 27261 12393 27295 12427
rect 27295 12393 27304 12427
rect 27252 12384 27304 12393
rect 29460 12384 29512 12436
rect 29828 12384 29880 12436
rect 8484 12316 8536 12368
rect 10140 12316 10192 12368
rect 10324 12316 10376 12368
rect 19616 12316 19668 12368
rect 20904 12316 20956 12368
rect 21272 12316 21324 12368
rect 23848 12316 23900 12368
rect 24124 12316 24176 12368
rect 24492 12359 24544 12368
rect 24492 12325 24501 12359
rect 24501 12325 24535 12359
rect 24535 12325 24544 12359
rect 24492 12316 24544 12325
rect 26240 12316 26292 12368
rect 7932 12248 7984 12300
rect 5540 12180 5592 12232
rect 6000 12155 6052 12164
rect 6000 12121 6009 12155
rect 6009 12121 6043 12155
rect 6043 12121 6052 12155
rect 6000 12112 6052 12121
rect 6460 12112 6512 12164
rect 6736 12155 6788 12164
rect 6736 12121 6745 12155
rect 6745 12121 6779 12155
rect 6779 12121 6788 12155
rect 6736 12112 6788 12121
rect 8116 12180 8168 12232
rect 13176 12291 13228 12300
rect 8760 12180 8812 12232
rect 11336 12180 11388 12232
rect 13176 12257 13185 12291
rect 13185 12257 13219 12291
rect 13219 12257 13228 12291
rect 13176 12248 13228 12257
rect 13728 12248 13780 12300
rect 18604 12248 18656 12300
rect 19340 12291 19392 12300
rect 14004 12180 14056 12232
rect 14280 12180 14332 12232
rect 14832 12180 14884 12232
rect 17040 12180 17092 12232
rect 17684 12180 17736 12232
rect 19340 12257 19349 12291
rect 19349 12257 19383 12291
rect 19383 12257 19392 12291
rect 19340 12248 19392 12257
rect 19432 12248 19484 12300
rect 20812 12248 20864 12300
rect 22100 12248 22152 12300
rect 24952 12248 25004 12300
rect 9404 12112 9456 12164
rect 7012 12087 7064 12096
rect 7012 12053 7021 12087
rect 7021 12053 7055 12087
rect 7055 12053 7064 12087
rect 7012 12044 7064 12053
rect 7380 12087 7432 12096
rect 7380 12053 7389 12087
rect 7389 12053 7423 12087
rect 7423 12053 7432 12087
rect 7380 12044 7432 12053
rect 7472 12087 7524 12096
rect 7472 12053 7481 12087
rect 7481 12053 7515 12087
rect 7515 12053 7524 12087
rect 7472 12044 7524 12053
rect 7932 12087 7984 12096
rect 7932 12053 7941 12087
rect 7941 12053 7975 12087
rect 7975 12053 7984 12087
rect 7932 12044 7984 12053
rect 8392 12044 8444 12096
rect 10692 12044 10744 12096
rect 13176 12112 13228 12164
rect 16580 12112 16632 12164
rect 17316 12112 17368 12164
rect 20352 12112 20404 12164
rect 22008 12180 22060 12232
rect 22192 12223 22244 12232
rect 22192 12189 22201 12223
rect 22201 12189 22235 12223
rect 22235 12189 22244 12223
rect 22192 12180 22244 12189
rect 22468 12180 22520 12232
rect 22928 12180 22980 12232
rect 23664 12180 23716 12232
rect 23480 12112 23532 12164
rect 19616 12044 19668 12096
rect 20168 12044 20220 12096
rect 22652 12044 22704 12096
rect 25780 12180 25832 12232
rect 26332 12180 26384 12232
rect 29644 12316 29696 12368
rect 32404 12384 32456 12436
rect 33140 12384 33192 12436
rect 32864 12359 32916 12368
rect 32864 12325 32873 12359
rect 32873 12325 32907 12359
rect 32907 12325 32916 12359
rect 32864 12316 32916 12325
rect 27528 12248 27580 12300
rect 29736 12248 29788 12300
rect 27896 12180 27948 12232
rect 27068 12112 27120 12164
rect 30104 12155 30156 12164
rect 30104 12121 30138 12155
rect 30138 12121 30156 12155
rect 30104 12112 30156 12121
rect 31392 12180 31444 12232
rect 33876 12248 33928 12300
rect 34428 12180 34480 12232
rect 32864 12112 32916 12164
rect 24860 12087 24912 12096
rect 24860 12053 24869 12087
rect 24869 12053 24903 12087
rect 24903 12053 24912 12087
rect 24860 12044 24912 12053
rect 25872 12087 25924 12096
rect 25872 12053 25881 12087
rect 25881 12053 25915 12087
rect 25915 12053 25924 12087
rect 25872 12044 25924 12053
rect 26424 12044 26476 12096
rect 27528 12044 27580 12096
rect 28264 12087 28316 12096
rect 28264 12053 28273 12087
rect 28273 12053 28307 12087
rect 28307 12053 28316 12087
rect 28264 12044 28316 12053
rect 30932 12044 30984 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 7932 11840 7984 11892
rect 11244 11840 11296 11892
rect 11336 11883 11388 11892
rect 11336 11849 11345 11883
rect 11345 11849 11379 11883
rect 11379 11849 11388 11883
rect 11336 11840 11388 11849
rect 13176 11883 13228 11892
rect 13176 11849 13185 11883
rect 13185 11849 13219 11883
rect 13219 11849 13228 11883
rect 13176 11840 13228 11849
rect 13544 11840 13596 11892
rect 16948 11840 17000 11892
rect 17132 11840 17184 11892
rect 18420 11840 18472 11892
rect 20352 11883 20404 11892
rect 20352 11849 20361 11883
rect 20361 11849 20395 11883
rect 20395 11849 20404 11883
rect 20352 11840 20404 11849
rect 20720 11883 20772 11892
rect 20720 11849 20729 11883
rect 20729 11849 20763 11883
rect 20763 11849 20772 11883
rect 20720 11840 20772 11849
rect 21088 11840 21140 11892
rect 3240 11772 3292 11824
rect 3700 11704 3752 11756
rect 5540 11772 5592 11824
rect 4896 11704 4948 11756
rect 6736 11704 6788 11756
rect 7656 11704 7708 11756
rect 9312 11704 9364 11756
rect 11152 11772 11204 11824
rect 10968 11704 11020 11756
rect 12348 11704 12400 11756
rect 12532 11772 12584 11824
rect 15476 11772 15528 11824
rect 14648 11747 14700 11756
rect 14648 11713 14657 11747
rect 14657 11713 14691 11747
rect 14691 11713 14700 11747
rect 14648 11704 14700 11713
rect 4620 11500 4672 11552
rect 5264 11500 5316 11552
rect 6092 11500 6144 11552
rect 8392 11543 8444 11552
rect 8392 11509 8401 11543
rect 8401 11509 8435 11543
rect 8435 11509 8444 11543
rect 8392 11500 8444 11509
rect 9772 11500 9824 11552
rect 10324 11500 10376 11552
rect 13912 11636 13964 11688
rect 14924 11747 14976 11756
rect 14924 11713 14933 11747
rect 14933 11713 14967 11747
rect 14967 11713 14976 11747
rect 14924 11704 14976 11713
rect 16580 11704 16632 11756
rect 17316 11704 17368 11756
rect 17500 11704 17552 11756
rect 17684 11772 17736 11824
rect 17868 11747 17920 11756
rect 17868 11713 17902 11747
rect 17902 11713 17920 11747
rect 17868 11704 17920 11713
rect 16672 11636 16724 11688
rect 20076 11636 20128 11688
rect 21364 11636 21416 11688
rect 22468 11772 22520 11824
rect 22100 11747 22152 11756
rect 22100 11713 22134 11747
rect 22134 11713 22152 11747
rect 22100 11704 22152 11713
rect 23480 11883 23532 11892
rect 23480 11849 23489 11883
rect 23489 11849 23523 11883
rect 23523 11849 23532 11883
rect 23480 11840 23532 11849
rect 23848 11883 23900 11892
rect 23848 11849 23857 11883
rect 23857 11849 23891 11883
rect 23891 11849 23900 11883
rect 23848 11840 23900 11849
rect 25044 11840 25096 11892
rect 25872 11840 25924 11892
rect 27252 11883 27304 11892
rect 27252 11849 27261 11883
rect 27261 11849 27295 11883
rect 27295 11849 27304 11883
rect 27252 11840 27304 11849
rect 23664 11772 23716 11824
rect 12532 11500 12584 11552
rect 12716 11500 12768 11552
rect 13544 11500 13596 11552
rect 14648 11500 14700 11552
rect 16948 11568 17000 11620
rect 17592 11568 17644 11620
rect 20352 11568 20404 11620
rect 23940 11679 23992 11688
rect 23940 11645 23949 11679
rect 23949 11645 23983 11679
rect 23983 11645 23992 11679
rect 23940 11636 23992 11645
rect 24676 11704 24728 11756
rect 25044 11747 25096 11756
rect 25044 11713 25053 11747
rect 25053 11713 25087 11747
rect 25087 11713 25096 11747
rect 25044 11704 25096 11713
rect 26148 11815 26200 11824
rect 26148 11781 26157 11815
rect 26157 11781 26191 11815
rect 26191 11781 26200 11815
rect 26148 11772 26200 11781
rect 23296 11568 23348 11620
rect 24400 11568 24452 11620
rect 26056 11636 26108 11688
rect 26516 11704 26568 11756
rect 27712 11747 27764 11756
rect 27712 11713 27721 11747
rect 27721 11713 27755 11747
rect 27755 11713 27764 11747
rect 27712 11704 27764 11713
rect 28172 11772 28224 11824
rect 30104 11883 30156 11892
rect 30104 11849 30113 11883
rect 30113 11849 30147 11883
rect 30147 11849 30156 11883
rect 30104 11840 30156 11849
rect 31392 11883 31444 11892
rect 31392 11849 31401 11883
rect 31401 11849 31435 11883
rect 31435 11849 31444 11883
rect 31392 11840 31444 11849
rect 31484 11883 31536 11892
rect 31484 11849 31493 11883
rect 31493 11849 31527 11883
rect 31527 11849 31536 11883
rect 31484 11840 31536 11849
rect 28724 11704 28776 11756
rect 29092 11747 29144 11756
rect 29092 11713 29110 11747
rect 29110 11713 29144 11747
rect 29092 11704 29144 11713
rect 30288 11704 30340 11756
rect 30932 11747 30984 11756
rect 30932 11713 30941 11747
rect 30941 11713 30975 11747
rect 30975 11713 30984 11747
rect 30932 11704 30984 11713
rect 31300 11704 31352 11756
rect 34520 11747 34572 11756
rect 34520 11713 34529 11747
rect 34529 11713 34563 11747
rect 34563 11713 34572 11747
rect 34520 11704 34572 11713
rect 26792 11636 26844 11688
rect 27620 11636 27672 11688
rect 28356 11636 28408 11688
rect 29828 11636 29880 11688
rect 30656 11679 30708 11688
rect 30656 11645 30665 11679
rect 30665 11645 30699 11679
rect 30699 11645 30708 11679
rect 30656 11636 30708 11645
rect 34796 11679 34848 11688
rect 34796 11645 34805 11679
rect 34805 11645 34839 11679
rect 34839 11645 34848 11679
rect 34796 11636 34848 11645
rect 27988 11611 28040 11620
rect 27988 11577 27997 11611
rect 27997 11577 28031 11611
rect 28031 11577 28040 11611
rect 27988 11568 28040 11577
rect 15200 11543 15252 11552
rect 15200 11509 15209 11543
rect 15209 11509 15243 11543
rect 15243 11509 15252 11543
rect 15200 11500 15252 11509
rect 16672 11543 16724 11552
rect 16672 11509 16681 11543
rect 16681 11509 16715 11543
rect 16715 11509 16724 11543
rect 16672 11500 16724 11509
rect 20720 11500 20772 11552
rect 22560 11500 22612 11552
rect 25504 11500 25556 11552
rect 26516 11543 26568 11552
rect 26516 11509 26525 11543
rect 26525 11509 26559 11543
rect 26559 11509 26568 11543
rect 26516 11500 26568 11509
rect 26700 11500 26752 11552
rect 29552 11500 29604 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 3700 11296 3752 11348
rect 4896 11339 4948 11348
rect 4896 11305 4905 11339
rect 4905 11305 4939 11339
rect 4939 11305 4948 11339
rect 4896 11296 4948 11305
rect 5080 11228 5132 11280
rect 4252 11203 4304 11212
rect 4252 11169 4261 11203
rect 4261 11169 4295 11203
rect 4295 11169 4304 11203
rect 4252 11160 4304 11169
rect 1308 11092 1360 11144
rect 4620 11092 4672 11144
rect 5264 11135 5316 11144
rect 5264 11101 5273 11135
rect 5273 11101 5307 11135
rect 5307 11101 5316 11135
rect 5264 11092 5316 11101
rect 6092 11228 6144 11280
rect 6736 11092 6788 11144
rect 3148 11067 3200 11076
rect 3148 11033 3157 11067
rect 3157 11033 3191 11067
rect 3191 11033 3200 11067
rect 3148 11024 3200 11033
rect 5080 11024 5132 11076
rect 7012 11024 7064 11076
rect 7380 11296 7432 11348
rect 7656 11339 7708 11348
rect 7656 11305 7665 11339
rect 7665 11305 7699 11339
rect 7699 11305 7708 11339
rect 7656 11296 7708 11305
rect 9312 11296 9364 11348
rect 7472 11160 7524 11212
rect 8208 11203 8260 11212
rect 8208 11169 8217 11203
rect 8217 11169 8251 11203
rect 8251 11169 8260 11203
rect 8208 11160 8260 11169
rect 8392 11092 8444 11144
rect 10416 11296 10468 11348
rect 10876 11296 10928 11348
rect 10968 11339 11020 11348
rect 10968 11305 10977 11339
rect 10977 11305 11011 11339
rect 11011 11305 11020 11339
rect 10968 11296 11020 11305
rect 12348 11339 12400 11348
rect 12348 11305 12357 11339
rect 12357 11305 12391 11339
rect 12391 11305 12400 11339
rect 12348 11296 12400 11305
rect 13912 11339 13964 11348
rect 13912 11305 13921 11339
rect 13921 11305 13955 11339
rect 13955 11305 13964 11339
rect 13912 11296 13964 11305
rect 14924 11296 14976 11348
rect 16120 11296 16172 11348
rect 17132 11296 17184 11348
rect 17592 11339 17644 11348
rect 17592 11305 17601 11339
rect 17601 11305 17635 11339
rect 17635 11305 17644 11339
rect 17592 11296 17644 11305
rect 17868 11296 17920 11348
rect 19616 11296 19668 11348
rect 20996 11296 21048 11348
rect 21732 11296 21784 11348
rect 22100 11296 22152 11348
rect 9680 11160 9732 11212
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 10140 11160 10192 11212
rect 12716 11228 12768 11280
rect 16948 11228 17000 11280
rect 26056 11296 26108 11348
rect 26332 11339 26384 11348
rect 26332 11305 26341 11339
rect 26341 11305 26375 11339
rect 26375 11305 26384 11339
rect 26332 11296 26384 11305
rect 26516 11296 26568 11348
rect 28540 11296 28592 11348
rect 29092 11339 29144 11348
rect 29092 11305 29101 11339
rect 29101 11305 29135 11339
rect 29135 11305 29144 11339
rect 29092 11296 29144 11305
rect 30656 11296 30708 11348
rect 27712 11228 27764 11280
rect 11244 11160 11296 11212
rect 12808 11160 12860 11212
rect 9772 11135 9824 11144
rect 9772 11101 9781 11135
rect 9781 11101 9815 11135
rect 9815 11101 9824 11135
rect 9772 11092 9824 11101
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 10416 11135 10468 11144
rect 10416 11101 10425 11135
rect 10425 11101 10459 11135
rect 10459 11101 10468 11135
rect 10416 11092 10468 11101
rect 10692 11135 10744 11144
rect 10692 11101 10701 11135
rect 10701 11101 10735 11135
rect 10735 11101 10744 11135
rect 10692 11092 10744 11101
rect 11152 11092 11204 11144
rect 11336 11135 11388 11144
rect 11336 11101 11345 11135
rect 11345 11101 11379 11135
rect 11379 11101 11388 11135
rect 11336 11092 11388 11101
rect 13176 11092 13228 11144
rect 13360 11135 13412 11144
rect 13360 11101 13369 11135
rect 13369 11101 13403 11135
rect 13403 11101 13412 11135
rect 13360 11092 13412 11101
rect 13544 11135 13596 11144
rect 13544 11101 13553 11135
rect 13553 11101 13587 11135
rect 13587 11101 13596 11135
rect 13544 11092 13596 11101
rect 13728 11135 13780 11144
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 17316 11160 17368 11212
rect 19616 11160 19668 11212
rect 22100 11160 22152 11212
rect 22928 11160 22980 11212
rect 15108 11092 15160 11144
rect 16672 11092 16724 11144
rect 18420 11135 18472 11144
rect 18420 11101 18429 11135
rect 18429 11101 18463 11135
rect 18463 11101 18472 11135
rect 18420 11092 18472 11101
rect 12440 11024 12492 11076
rect 13912 11024 13964 11076
rect 15476 11024 15528 11076
rect 15752 11024 15804 11076
rect 19616 11067 19668 11076
rect 19616 11033 19625 11067
rect 19625 11033 19659 11067
rect 19659 11033 19668 11067
rect 22468 11092 22520 11144
rect 23296 11092 23348 11144
rect 23388 11092 23440 11144
rect 26148 11092 26200 11144
rect 27620 11160 27672 11212
rect 27804 11203 27856 11212
rect 27804 11169 27813 11203
rect 27813 11169 27847 11203
rect 27847 11169 27856 11203
rect 27804 11160 27856 11169
rect 27436 11092 27488 11144
rect 27712 11092 27764 11144
rect 28080 11160 28132 11212
rect 28632 11160 28684 11212
rect 30748 11160 30800 11212
rect 27988 11092 28040 11144
rect 29552 11135 29604 11144
rect 29552 11101 29561 11135
rect 29561 11101 29595 11135
rect 29595 11101 29604 11135
rect 29552 11092 29604 11101
rect 29644 11092 29696 11144
rect 30196 11092 30248 11144
rect 34152 11135 34204 11144
rect 34152 11101 34161 11135
rect 34161 11101 34195 11135
rect 34195 11101 34204 11135
rect 34152 11092 34204 11101
rect 34428 11135 34480 11144
rect 34428 11101 34437 11135
rect 34437 11101 34471 11135
rect 34471 11101 34480 11135
rect 34428 11092 34480 11101
rect 19616 11024 19668 11033
rect 22100 11067 22152 11076
rect 22100 11033 22109 11067
rect 22109 11033 22143 11067
rect 22143 11033 22152 11067
rect 22100 11024 22152 11033
rect 22652 11067 22704 11076
rect 22652 11033 22661 11067
rect 22661 11033 22695 11067
rect 22695 11033 22704 11067
rect 22652 11024 22704 11033
rect 23940 11024 23992 11076
rect 24952 11024 25004 11076
rect 4344 10956 4396 11008
rect 5172 10956 5224 11008
rect 5448 10956 5500 11008
rect 8668 10956 8720 11008
rect 14004 10956 14056 11008
rect 14832 10956 14884 11008
rect 17776 10956 17828 11008
rect 20628 10956 20680 11008
rect 22376 10956 22428 11008
rect 25504 10956 25556 11008
rect 27160 11024 27212 11076
rect 27528 11024 27580 11076
rect 27620 11067 27672 11076
rect 27620 11033 27629 11067
rect 27629 11033 27663 11067
rect 27663 11033 27672 11067
rect 27620 11024 27672 11033
rect 26976 10999 27028 11008
rect 26976 10965 26985 10999
rect 26985 10965 27019 10999
rect 27019 10965 27028 10999
rect 26976 10956 27028 10965
rect 34520 11024 34572 11076
rect 34980 11024 35032 11076
rect 28080 10999 28132 11008
rect 28080 10965 28089 10999
rect 28089 10965 28123 10999
rect 28123 10965 28132 10999
rect 28080 10956 28132 10965
rect 28264 10956 28316 11008
rect 33508 10956 33560 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 3608 10752 3660 10804
rect 4252 10752 4304 10804
rect 3240 10659 3292 10668
rect 3240 10625 3249 10659
rect 3249 10625 3283 10659
rect 3283 10625 3292 10659
rect 3240 10616 3292 10625
rect 4160 10659 4212 10668
rect 4160 10625 4169 10659
rect 4169 10625 4203 10659
rect 4203 10625 4212 10659
rect 4160 10616 4212 10625
rect 4252 10548 4304 10600
rect 5080 10752 5132 10804
rect 5264 10727 5316 10736
rect 5264 10693 5273 10727
rect 5273 10693 5307 10727
rect 5307 10693 5316 10727
rect 5264 10684 5316 10693
rect 5724 10795 5776 10804
rect 5724 10761 5733 10795
rect 5733 10761 5767 10795
rect 5767 10761 5776 10795
rect 5724 10752 5776 10761
rect 8760 10752 8812 10804
rect 10048 10752 10100 10804
rect 10416 10752 10468 10804
rect 11152 10795 11204 10804
rect 11152 10761 11161 10795
rect 11161 10761 11195 10795
rect 11195 10761 11204 10795
rect 11152 10752 11204 10761
rect 12808 10752 12860 10804
rect 14832 10752 14884 10804
rect 15752 10795 15804 10804
rect 15752 10761 15761 10795
rect 15761 10761 15795 10795
rect 15795 10761 15804 10795
rect 15752 10752 15804 10761
rect 16120 10795 16172 10804
rect 16120 10761 16129 10795
rect 16129 10761 16163 10795
rect 16163 10761 16172 10795
rect 16120 10752 16172 10761
rect 12440 10684 12492 10736
rect 14740 10727 14792 10736
rect 14740 10693 14749 10727
rect 14749 10693 14783 10727
rect 14783 10693 14792 10727
rect 14740 10684 14792 10693
rect 15476 10727 15528 10736
rect 15476 10693 15485 10727
rect 15485 10693 15519 10727
rect 15519 10693 15528 10727
rect 15476 10684 15528 10693
rect 17132 10727 17184 10736
rect 17132 10693 17141 10727
rect 17141 10693 17175 10727
rect 17175 10693 17184 10727
rect 17132 10684 17184 10693
rect 19432 10684 19484 10736
rect 4620 10548 4672 10600
rect 5724 10548 5776 10600
rect 5908 10616 5960 10668
rect 4804 10480 4856 10532
rect 4896 10412 4948 10464
rect 5540 10455 5592 10464
rect 5540 10421 5549 10455
rect 5549 10421 5583 10455
rect 5583 10421 5592 10455
rect 5540 10412 5592 10421
rect 10048 10548 10100 10600
rect 12256 10548 12308 10600
rect 14556 10548 14608 10600
rect 16764 10616 16816 10668
rect 16948 10616 17000 10668
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 18328 10616 18380 10668
rect 16856 10548 16908 10600
rect 20352 10616 20404 10668
rect 23388 10752 23440 10804
rect 24952 10795 25004 10804
rect 24952 10761 24961 10795
rect 24961 10761 24995 10795
rect 24995 10761 25004 10795
rect 24952 10752 25004 10761
rect 26056 10752 26108 10804
rect 26976 10795 27028 10804
rect 26976 10761 26985 10795
rect 26985 10761 27019 10795
rect 27019 10761 27028 10795
rect 26976 10752 27028 10761
rect 23848 10684 23900 10736
rect 23940 10684 23992 10736
rect 20628 10548 20680 10600
rect 21364 10659 21416 10668
rect 21364 10625 21373 10659
rect 21373 10625 21407 10659
rect 21407 10625 21416 10659
rect 21364 10616 21416 10625
rect 21732 10616 21784 10668
rect 10048 10412 10100 10464
rect 10784 10412 10836 10464
rect 12164 10412 12216 10464
rect 13820 10412 13872 10464
rect 16028 10412 16080 10464
rect 21916 10548 21968 10600
rect 25596 10616 25648 10668
rect 25504 10591 25556 10600
rect 25504 10557 25513 10591
rect 25513 10557 25547 10591
rect 25547 10557 25556 10591
rect 25504 10548 25556 10557
rect 29000 10752 29052 10804
rect 29644 10752 29696 10804
rect 27528 10616 27580 10668
rect 29092 10684 29144 10736
rect 30288 10752 30340 10804
rect 34980 10795 35032 10804
rect 34980 10761 34989 10795
rect 34989 10761 35023 10795
rect 35023 10761 35032 10795
rect 34980 10752 35032 10761
rect 30196 10684 30248 10736
rect 29000 10616 29052 10668
rect 29276 10616 29328 10668
rect 29828 10591 29880 10600
rect 29828 10557 29837 10591
rect 29837 10557 29871 10591
rect 29871 10557 29880 10591
rect 29828 10548 29880 10557
rect 20812 10412 20864 10464
rect 21088 10455 21140 10464
rect 21088 10421 21097 10455
rect 21097 10421 21131 10455
rect 21131 10421 21140 10455
rect 21088 10412 21140 10421
rect 21824 10412 21876 10464
rect 23848 10412 23900 10464
rect 29184 10412 29236 10464
rect 33508 10727 33560 10736
rect 33508 10693 33517 10727
rect 33517 10693 33551 10727
rect 33551 10693 33560 10727
rect 33508 10684 33560 10693
rect 34520 10684 34572 10736
rect 32772 10548 32824 10600
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 3608 10251 3660 10260
rect 3608 10217 3617 10251
rect 3617 10217 3651 10251
rect 3651 10217 3660 10251
rect 3608 10208 3660 10217
rect 4896 10251 4948 10260
rect 4896 10217 4905 10251
rect 4905 10217 4939 10251
rect 4939 10217 4948 10251
rect 4896 10208 4948 10217
rect 5632 10208 5684 10260
rect 8668 10251 8720 10260
rect 8668 10217 8677 10251
rect 8677 10217 8711 10251
rect 8711 10217 8720 10251
rect 8668 10208 8720 10217
rect 8760 10208 8812 10260
rect 10416 10208 10468 10260
rect 11520 10208 11572 10260
rect 4712 10183 4764 10192
rect 4344 10072 4396 10124
rect 4712 10149 4721 10183
rect 4721 10149 4755 10183
rect 4755 10149 4764 10183
rect 4712 10140 4764 10149
rect 4252 10004 4304 10056
rect 4712 10004 4764 10056
rect 5080 10047 5132 10056
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 5080 10004 5132 10013
rect 9956 10140 10008 10192
rect 3792 9911 3844 9920
rect 3792 9877 3801 9911
rect 3801 9877 3835 9911
rect 3835 9877 3844 9911
rect 3792 9868 3844 9877
rect 4804 9936 4856 9988
rect 5724 10004 5776 10056
rect 5632 9936 5684 9988
rect 6368 9979 6420 9988
rect 6368 9945 6377 9979
rect 6377 9945 6411 9979
rect 6411 9945 6420 9979
rect 6368 9936 6420 9945
rect 5908 9868 5960 9920
rect 7840 10047 7892 10056
rect 7840 10013 7847 10047
rect 7847 10013 7892 10047
rect 7840 10004 7892 10013
rect 8668 10004 8720 10056
rect 9772 10072 9824 10124
rect 10876 10115 10928 10124
rect 10876 10081 10885 10115
rect 10885 10081 10919 10115
rect 10919 10081 10928 10115
rect 10876 10072 10928 10081
rect 10048 10004 10100 10056
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 10508 10047 10560 10056
rect 10508 10013 10553 10047
rect 10553 10013 10560 10047
rect 10508 10004 10560 10013
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 11796 10208 11848 10260
rect 13912 10251 13964 10260
rect 13912 10217 13921 10251
rect 13921 10217 13955 10251
rect 13955 10217 13964 10251
rect 13912 10208 13964 10217
rect 14464 10208 14516 10260
rect 17040 10208 17092 10260
rect 12164 10115 12216 10124
rect 12164 10081 12173 10115
rect 12173 10081 12207 10115
rect 12207 10081 12216 10115
rect 12164 10072 12216 10081
rect 12256 10115 12308 10124
rect 12256 10081 12265 10115
rect 12265 10081 12299 10115
rect 12299 10081 12308 10115
rect 12256 10072 12308 10081
rect 12532 10115 12584 10124
rect 12532 10081 12541 10115
rect 12541 10081 12575 10115
rect 12575 10081 12584 10115
rect 12532 10072 12584 10081
rect 13820 10072 13872 10124
rect 14556 10115 14608 10124
rect 14556 10081 14565 10115
rect 14565 10081 14599 10115
rect 14599 10081 14608 10115
rect 14556 10072 14608 10081
rect 14832 10072 14884 10124
rect 15476 10072 15528 10124
rect 13636 10004 13688 10056
rect 8024 9979 8076 9988
rect 8024 9945 8033 9979
rect 8033 9945 8067 9979
rect 8067 9945 8076 9979
rect 8024 9936 8076 9945
rect 9404 9936 9456 9988
rect 10140 9936 10192 9988
rect 9588 9868 9640 9920
rect 10048 9911 10100 9920
rect 10048 9877 10057 9911
rect 10057 9877 10091 9911
rect 10091 9877 10100 9911
rect 10048 9868 10100 9877
rect 11704 9911 11756 9920
rect 11704 9877 11713 9911
rect 11713 9877 11747 9911
rect 11747 9877 11756 9911
rect 11704 9868 11756 9877
rect 14464 10047 14516 10056
rect 14464 10013 14473 10047
rect 14473 10013 14507 10047
rect 14507 10013 14516 10047
rect 14464 10004 14516 10013
rect 16028 10047 16080 10056
rect 16028 10013 16062 10047
rect 16062 10013 16080 10047
rect 16028 10004 16080 10013
rect 17776 10208 17828 10260
rect 17408 10140 17460 10192
rect 18420 10140 18472 10192
rect 22284 10208 22336 10260
rect 23572 10208 23624 10260
rect 17408 10047 17460 10056
rect 17408 10013 17417 10047
rect 17417 10013 17451 10047
rect 17451 10013 17460 10047
rect 17408 10004 17460 10013
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 13360 9868 13412 9920
rect 18788 9936 18840 9988
rect 17316 9868 17368 9920
rect 18328 9868 18380 9920
rect 25504 10140 25556 10192
rect 26792 10208 26844 10260
rect 27160 10208 27212 10260
rect 27528 10208 27580 10260
rect 27712 10251 27764 10260
rect 27712 10217 27721 10251
rect 27721 10217 27755 10251
rect 27755 10217 27764 10251
rect 27712 10208 27764 10217
rect 27804 10208 27856 10260
rect 28632 10208 28684 10260
rect 29092 10208 29144 10260
rect 29828 10208 29880 10260
rect 28172 10140 28224 10192
rect 20352 10115 20404 10124
rect 20352 10081 20361 10115
rect 20361 10081 20395 10115
rect 20395 10081 20404 10115
rect 20352 10072 20404 10081
rect 22468 10072 22520 10124
rect 19800 10004 19852 10056
rect 22376 10004 22428 10056
rect 22560 10004 22612 10056
rect 20628 9979 20680 9988
rect 20628 9945 20662 9979
rect 20662 9945 20680 9979
rect 20628 9936 20680 9945
rect 21916 9936 21968 9988
rect 20996 9868 21048 9920
rect 21364 9868 21416 9920
rect 23020 10047 23072 10056
rect 23020 10013 23029 10047
rect 23029 10013 23063 10047
rect 23063 10013 23072 10047
rect 23020 10004 23072 10013
rect 26792 10115 26844 10124
rect 26792 10081 26801 10115
rect 26801 10081 26835 10115
rect 26835 10081 26844 10115
rect 26792 10072 26844 10081
rect 23296 10047 23348 10056
rect 23296 10013 23305 10047
rect 23305 10013 23339 10047
rect 23339 10013 23348 10047
rect 23296 10004 23348 10013
rect 23480 10047 23532 10056
rect 23480 10013 23489 10047
rect 23489 10013 23523 10047
rect 23523 10013 23532 10047
rect 23480 10004 23532 10013
rect 24400 10047 24452 10056
rect 24400 10013 24409 10047
rect 24409 10013 24443 10047
rect 24443 10013 24452 10047
rect 24400 10004 24452 10013
rect 24768 10004 24820 10056
rect 26976 10004 27028 10056
rect 27160 10004 27212 10056
rect 28080 10004 28132 10056
rect 28816 10047 28868 10056
rect 28816 10013 28820 10047
rect 28820 10013 28854 10047
rect 28854 10013 28868 10047
rect 28816 10004 28868 10013
rect 29000 10047 29052 10056
rect 29000 10013 29009 10047
rect 29009 10013 29043 10047
rect 29043 10013 29052 10047
rect 29000 10004 29052 10013
rect 29184 10047 29236 10056
rect 29184 10013 29192 10047
rect 29192 10013 29226 10047
rect 29226 10013 29236 10047
rect 29184 10004 29236 10013
rect 29276 10047 29328 10056
rect 29276 10013 29285 10047
rect 29285 10013 29319 10047
rect 29319 10013 29328 10047
rect 29276 10004 29328 10013
rect 29644 10047 29696 10056
rect 29644 10013 29653 10047
rect 29653 10013 29687 10047
rect 29687 10013 29696 10047
rect 29644 10004 29696 10013
rect 29828 10004 29880 10056
rect 23204 9868 23256 9920
rect 27896 9936 27948 9988
rect 28908 9979 28960 9988
rect 28908 9945 28917 9979
rect 28917 9945 28951 9979
rect 28951 9945 28960 9979
rect 28908 9936 28960 9945
rect 31208 9979 31260 9988
rect 31208 9945 31217 9979
rect 31217 9945 31251 9979
rect 31251 9945 31260 9979
rect 31208 9936 31260 9945
rect 32772 9936 32824 9988
rect 27252 9868 27304 9920
rect 28264 9868 28316 9920
rect 28540 9868 28592 9920
rect 29736 9911 29788 9920
rect 29736 9877 29745 9911
rect 29745 9877 29779 9911
rect 29779 9877 29788 9911
rect 30472 9911 30524 9920
rect 29736 9868 29788 9877
rect 30472 9877 30481 9911
rect 30481 9877 30515 9911
rect 30515 9877 30524 9911
rect 30472 9868 30524 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 4344 9707 4396 9716
rect 4344 9673 4353 9707
rect 4353 9673 4387 9707
rect 4387 9673 4396 9707
rect 4344 9664 4396 9673
rect 5632 9664 5684 9716
rect 3792 9596 3844 9648
rect 3976 9528 4028 9580
rect 5540 9596 5592 9648
rect 5724 9596 5776 9648
rect 7840 9664 7892 9716
rect 9772 9707 9824 9716
rect 9772 9673 9781 9707
rect 9781 9673 9815 9707
rect 9815 9673 9824 9707
rect 9772 9664 9824 9673
rect 10508 9664 10560 9716
rect 13360 9664 13412 9716
rect 14832 9664 14884 9716
rect 20628 9707 20680 9716
rect 20628 9673 20637 9707
rect 20637 9673 20671 9707
rect 20671 9673 20680 9707
rect 20628 9664 20680 9673
rect 20996 9707 21048 9716
rect 20996 9673 21005 9707
rect 21005 9673 21039 9707
rect 21039 9673 21048 9707
rect 20996 9664 21048 9673
rect 4620 9528 4672 9580
rect 3884 9503 3936 9512
rect 3884 9469 3893 9503
rect 3893 9469 3927 9503
rect 3927 9469 3936 9503
rect 3884 9460 3936 9469
rect 4252 9460 4304 9512
rect 6368 9528 6420 9580
rect 6644 9571 6696 9580
rect 6644 9537 6653 9571
rect 6653 9537 6687 9571
rect 6687 9537 6696 9571
rect 6644 9528 6696 9537
rect 6736 9528 6788 9580
rect 7380 9528 7432 9580
rect 8944 9528 8996 9580
rect 11060 9571 11112 9580
rect 11060 9537 11078 9571
rect 11078 9537 11112 9571
rect 11060 9528 11112 9537
rect 11704 9596 11756 9648
rect 14372 9596 14424 9648
rect 20352 9596 20404 9648
rect 20720 9596 20772 9648
rect 22560 9664 22612 9716
rect 23296 9664 23348 9716
rect 22468 9596 22520 9648
rect 22652 9596 22704 9648
rect 24308 9664 24360 9716
rect 23480 9596 23532 9648
rect 24216 9639 24268 9648
rect 24216 9605 24225 9639
rect 24225 9605 24259 9639
rect 24259 9605 24268 9639
rect 24216 9596 24268 9605
rect 4068 9392 4120 9444
rect 5908 9503 5960 9512
rect 5908 9469 5917 9503
rect 5917 9469 5951 9503
rect 5951 9469 5960 9503
rect 5908 9460 5960 9469
rect 6092 9503 6144 9512
rect 6092 9469 6101 9503
rect 6101 9469 6135 9503
rect 6135 9469 6144 9503
rect 6092 9460 6144 9469
rect 8208 9460 8260 9512
rect 11520 9460 11572 9512
rect 15200 9528 15252 9580
rect 15476 9528 15528 9580
rect 17684 9571 17736 9580
rect 17684 9537 17718 9571
rect 17718 9537 17736 9571
rect 17684 9528 17736 9537
rect 19892 9528 19944 9580
rect 16764 9503 16816 9512
rect 3976 9367 4028 9376
rect 3976 9333 3985 9367
rect 3985 9333 4019 9367
rect 4019 9333 4028 9367
rect 3976 9324 4028 9333
rect 5448 9367 5500 9376
rect 5448 9333 5457 9367
rect 5457 9333 5491 9367
rect 5491 9333 5500 9367
rect 5448 9324 5500 9333
rect 9404 9392 9456 9444
rect 16764 9469 16773 9503
rect 16773 9469 16807 9503
rect 16807 9469 16816 9503
rect 16764 9460 16816 9469
rect 7472 9324 7524 9376
rect 10140 9324 10192 9376
rect 18788 9435 18840 9444
rect 18788 9401 18797 9435
rect 18797 9401 18831 9435
rect 18831 9401 18840 9435
rect 18788 9392 18840 9401
rect 14924 9367 14976 9376
rect 14924 9333 14933 9367
rect 14933 9333 14967 9367
rect 14967 9333 14976 9367
rect 14924 9324 14976 9333
rect 19984 9324 20036 9376
rect 22376 9528 22428 9580
rect 23020 9528 23072 9580
rect 23204 9571 23256 9580
rect 23204 9537 23213 9571
rect 23213 9537 23247 9571
rect 23247 9537 23256 9571
rect 23204 9528 23256 9537
rect 23572 9528 23624 9580
rect 24124 9571 24176 9580
rect 24124 9537 24133 9571
rect 24133 9537 24167 9571
rect 24167 9537 24176 9571
rect 24124 9528 24176 9537
rect 24400 9571 24452 9580
rect 24400 9537 24409 9571
rect 24409 9537 24443 9571
rect 24443 9537 24452 9571
rect 24400 9528 24452 9537
rect 20536 9460 20588 9512
rect 20996 9460 21048 9512
rect 21824 9503 21876 9512
rect 21824 9469 21833 9503
rect 21833 9469 21867 9503
rect 21867 9469 21876 9503
rect 21824 9460 21876 9469
rect 25228 9639 25280 9648
rect 25228 9605 25237 9639
rect 25237 9605 25271 9639
rect 25271 9605 25280 9639
rect 25228 9596 25280 9605
rect 26608 9596 26660 9648
rect 25136 9571 25188 9580
rect 25136 9537 25145 9571
rect 25145 9537 25179 9571
rect 25179 9537 25188 9571
rect 25136 9528 25188 9537
rect 25320 9571 25372 9580
rect 25320 9537 25329 9571
rect 25329 9537 25363 9571
rect 25363 9537 25372 9571
rect 25320 9528 25372 9537
rect 23112 9392 23164 9444
rect 22100 9324 22152 9376
rect 22652 9324 22704 9376
rect 24032 9392 24084 9444
rect 25504 9460 25556 9512
rect 26516 9571 26568 9580
rect 26516 9537 26525 9571
rect 26525 9537 26559 9571
rect 26559 9537 26568 9571
rect 26516 9528 26568 9537
rect 26884 9596 26936 9648
rect 27620 9596 27672 9648
rect 31208 9664 31260 9716
rect 28908 9596 28960 9648
rect 28264 9528 28316 9580
rect 27804 9460 27856 9512
rect 29828 9571 29880 9580
rect 29828 9537 29837 9571
rect 29837 9537 29871 9571
rect 29871 9537 29880 9571
rect 29828 9528 29880 9537
rect 34060 9571 34112 9580
rect 34060 9537 34069 9571
rect 34069 9537 34103 9571
rect 34103 9537 34112 9571
rect 34060 9528 34112 9537
rect 34244 9571 34296 9580
rect 34244 9537 34253 9571
rect 34253 9537 34287 9571
rect 34287 9537 34296 9571
rect 34244 9528 34296 9537
rect 34428 9528 34480 9580
rect 25412 9392 25464 9444
rect 26332 9435 26384 9444
rect 26332 9401 26341 9435
rect 26341 9401 26375 9435
rect 26375 9401 26384 9435
rect 26332 9392 26384 9401
rect 28172 9392 28224 9444
rect 30288 9460 30340 9512
rect 30472 9503 30524 9512
rect 30472 9469 30481 9503
rect 30481 9469 30515 9503
rect 30515 9469 30524 9503
rect 30472 9460 30524 9469
rect 23756 9324 23808 9376
rect 23848 9367 23900 9376
rect 23848 9333 23857 9367
rect 23857 9333 23891 9367
rect 23891 9333 23900 9367
rect 23848 9324 23900 9333
rect 24124 9324 24176 9376
rect 25504 9324 25556 9376
rect 26792 9324 26844 9376
rect 27804 9324 27856 9376
rect 28080 9324 28132 9376
rect 33048 9324 33100 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 4712 9120 4764 9172
rect 5540 9120 5592 9172
rect 6368 9120 6420 9172
rect 7380 9163 7432 9172
rect 7380 9129 7389 9163
rect 7389 9129 7423 9163
rect 7423 9129 7432 9163
rect 7380 9120 7432 9129
rect 8944 9163 8996 9172
rect 8944 9129 8953 9163
rect 8953 9129 8987 9163
rect 8987 9129 8996 9163
rect 8944 9120 8996 9129
rect 10048 9163 10100 9172
rect 10048 9129 10057 9163
rect 10057 9129 10091 9163
rect 10091 9129 10100 9163
rect 10048 9120 10100 9129
rect 6644 8984 6696 9036
rect 9404 9052 9456 9104
rect 11060 9120 11112 9172
rect 13084 9120 13136 9172
rect 13636 9163 13688 9172
rect 13636 9129 13645 9163
rect 13645 9129 13679 9163
rect 13679 9129 13688 9163
rect 13636 9120 13688 9129
rect 14924 9163 14976 9172
rect 14924 9129 14933 9163
rect 14933 9129 14967 9163
rect 14967 9129 14976 9163
rect 14924 9120 14976 9129
rect 17684 9120 17736 9172
rect 19984 9120 20036 9172
rect 21824 9120 21876 9172
rect 22008 9120 22060 9172
rect 22652 9120 22704 9172
rect 15568 9052 15620 9104
rect 25320 9120 25372 9172
rect 29276 9120 29328 9172
rect 34244 9120 34296 9172
rect 9680 8984 9732 9036
rect 1308 8916 1360 8968
rect 3884 8916 3936 8968
rect 4068 8959 4120 8968
rect 4068 8925 4102 8959
rect 4102 8925 4120 8959
rect 4068 8916 4120 8925
rect 5448 8848 5500 8900
rect 6828 8959 6880 8968
rect 6828 8925 6837 8959
rect 6837 8925 6871 8959
rect 6871 8925 6880 8959
rect 6828 8916 6880 8925
rect 7840 8916 7892 8968
rect 9772 8916 9824 8968
rect 10232 8984 10284 9036
rect 10508 9027 10560 9036
rect 10508 8993 10517 9027
rect 10517 8993 10551 9027
rect 10551 8993 10560 9027
rect 10508 8984 10560 8993
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 10140 8916 10192 8968
rect 12716 8959 12768 8968
rect 12716 8925 12725 8959
rect 12725 8925 12759 8959
rect 12759 8925 12768 8959
rect 12716 8916 12768 8925
rect 12808 8916 12860 8968
rect 13084 8959 13136 8968
rect 13084 8925 13093 8959
rect 13093 8925 13127 8959
rect 13127 8925 13136 8959
rect 13084 8916 13136 8925
rect 10876 8848 10928 8900
rect 16396 8984 16448 9036
rect 16856 8984 16908 9036
rect 18328 9027 18380 9036
rect 18328 8993 18337 9027
rect 18337 8993 18371 9027
rect 18371 8993 18380 9027
rect 18328 8984 18380 8993
rect 20812 8984 20864 9036
rect 6736 8780 6788 8832
rect 7472 8780 7524 8832
rect 7748 8780 7800 8832
rect 9588 8780 9640 8832
rect 9680 8780 9732 8832
rect 10324 8780 10376 8832
rect 10508 8780 10560 8832
rect 10784 8780 10836 8832
rect 11336 8780 11388 8832
rect 13176 8780 13228 8832
rect 14464 8959 14516 8968
rect 14464 8925 14471 8959
rect 14471 8925 14516 8959
rect 14464 8916 14516 8925
rect 14648 8959 14700 8968
rect 14648 8925 14657 8959
rect 14657 8925 14691 8959
rect 14691 8925 14700 8959
rect 14648 8916 14700 8925
rect 15016 8916 15068 8968
rect 17868 8916 17920 8968
rect 18788 8916 18840 8968
rect 18880 8916 18932 8968
rect 14004 8848 14056 8900
rect 20720 8916 20772 8968
rect 20996 8984 21048 9036
rect 21272 9027 21324 9036
rect 21272 8993 21281 9027
rect 21281 8993 21315 9027
rect 21315 8993 21324 9027
rect 21272 8984 21324 8993
rect 21824 9027 21876 9036
rect 21824 8993 21833 9027
rect 21833 8993 21867 9027
rect 21867 8993 21876 9027
rect 21824 8984 21876 8993
rect 22008 8984 22060 9036
rect 22376 8984 22428 9036
rect 21640 8916 21692 8968
rect 21732 8959 21784 8968
rect 21732 8925 21741 8959
rect 21741 8925 21775 8959
rect 21775 8925 21784 8959
rect 21732 8916 21784 8925
rect 24400 9095 24452 9104
rect 24400 9061 24409 9095
rect 24409 9061 24443 9095
rect 24443 9061 24452 9095
rect 24400 9052 24452 9061
rect 24584 9052 24636 9104
rect 13452 8780 13504 8832
rect 16856 8780 16908 8832
rect 16948 8780 17000 8832
rect 19156 8780 19208 8832
rect 20628 8780 20680 8832
rect 21272 8848 21324 8900
rect 21548 8780 21600 8832
rect 22100 8780 22152 8832
rect 22284 8823 22336 8832
rect 22284 8789 22293 8823
rect 22293 8789 22327 8823
rect 22327 8789 22336 8823
rect 22284 8780 22336 8789
rect 22468 8823 22520 8832
rect 22468 8789 22477 8823
rect 22477 8789 22511 8823
rect 22511 8789 22520 8823
rect 22468 8780 22520 8789
rect 22652 8848 22704 8900
rect 23848 8916 23900 8968
rect 24860 8984 24912 9036
rect 27160 9052 27212 9104
rect 27252 8984 27304 9036
rect 27804 9027 27856 9036
rect 27804 8993 27813 9027
rect 27813 8993 27847 9027
rect 27847 8993 27856 9027
rect 27804 8984 27856 8993
rect 24492 8780 24544 8832
rect 28080 8916 28132 8968
rect 28724 9052 28776 9104
rect 33048 9027 33100 9036
rect 33048 8993 33057 9027
rect 33057 8993 33091 9027
rect 33091 8993 33100 9027
rect 33048 8984 33100 8993
rect 28172 8891 28224 8900
rect 28172 8857 28181 8891
rect 28181 8857 28215 8891
rect 28215 8857 28224 8891
rect 28172 8848 28224 8857
rect 32772 8959 32824 8968
rect 32772 8925 32781 8959
rect 32781 8925 32815 8959
rect 32815 8925 32824 8959
rect 32772 8916 32824 8925
rect 33140 8848 33192 8900
rect 28356 8780 28408 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 4620 8619 4672 8628
rect 4620 8585 4629 8619
rect 4629 8585 4663 8619
rect 4663 8585 4672 8619
rect 4620 8576 4672 8585
rect 9864 8576 9916 8628
rect 10692 8576 10744 8628
rect 6000 8508 6052 8560
rect 3884 8440 3936 8492
rect 6920 8440 6972 8492
rect 8208 8440 8260 8492
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 10140 8483 10192 8492
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 10876 8576 10928 8628
rect 5264 8372 5316 8424
rect 11336 8372 11388 8424
rect 3976 8304 4028 8356
rect 14372 8576 14424 8628
rect 14464 8576 14516 8628
rect 17408 8576 17460 8628
rect 17500 8576 17552 8628
rect 17776 8619 17828 8628
rect 17776 8585 17785 8619
rect 17785 8585 17819 8619
rect 17819 8585 17828 8619
rect 17776 8576 17828 8585
rect 11520 8372 11572 8424
rect 12348 8440 12400 8492
rect 13176 8440 13228 8492
rect 14188 8440 14240 8492
rect 13636 8415 13688 8424
rect 13636 8381 13645 8415
rect 13645 8381 13679 8415
rect 13679 8381 13688 8415
rect 13636 8372 13688 8381
rect 15476 8508 15528 8560
rect 15568 8508 15620 8560
rect 16948 8440 17000 8492
rect 12808 8236 12860 8288
rect 14280 8236 14332 8288
rect 14924 8236 14976 8288
rect 18052 8483 18104 8492
rect 18052 8449 18061 8483
rect 18061 8449 18095 8483
rect 18095 8449 18104 8483
rect 18052 8440 18104 8449
rect 19156 8576 19208 8628
rect 18420 8483 18472 8492
rect 18420 8449 18429 8483
rect 18429 8449 18463 8483
rect 18463 8449 18472 8483
rect 18420 8440 18472 8449
rect 19248 8508 19300 8560
rect 19892 8508 19944 8560
rect 20812 8551 20864 8560
rect 20812 8517 20821 8551
rect 20821 8517 20855 8551
rect 20855 8517 20864 8551
rect 20812 8508 20864 8517
rect 21732 8576 21784 8628
rect 22100 8576 22152 8628
rect 22744 8619 22796 8628
rect 22744 8585 22753 8619
rect 22753 8585 22787 8619
rect 22787 8585 22796 8619
rect 22744 8576 22796 8585
rect 22836 8619 22888 8628
rect 22836 8585 22845 8619
rect 22845 8585 22879 8619
rect 22879 8585 22888 8619
rect 22836 8576 22888 8585
rect 23112 8619 23164 8628
rect 23112 8585 23121 8619
rect 23121 8585 23155 8619
rect 23155 8585 23164 8619
rect 23112 8576 23164 8585
rect 23388 8576 23440 8628
rect 26792 8576 26844 8628
rect 28080 8576 28132 8628
rect 28172 8576 28224 8628
rect 20628 8483 20680 8492
rect 20628 8449 20635 8483
rect 20635 8449 20680 8483
rect 18604 8347 18656 8356
rect 18604 8313 18613 8347
rect 18613 8313 18647 8347
rect 18647 8313 18656 8347
rect 18604 8304 18656 8313
rect 19984 8372 20036 8424
rect 20628 8440 20680 8449
rect 20720 8483 20772 8492
rect 20720 8449 20729 8483
rect 20729 8449 20763 8483
rect 20763 8449 20772 8483
rect 20720 8440 20772 8449
rect 21548 8440 21600 8492
rect 21916 8440 21968 8492
rect 27436 8508 27488 8560
rect 27804 8508 27856 8560
rect 33140 8508 33192 8560
rect 34796 8551 34848 8560
rect 34796 8517 34805 8551
rect 34805 8517 34839 8551
rect 34839 8517 34848 8551
rect 34796 8508 34848 8517
rect 22560 8440 22612 8492
rect 23112 8440 23164 8492
rect 23388 8440 23440 8492
rect 23480 8483 23532 8492
rect 23480 8449 23489 8483
rect 23489 8449 23523 8483
rect 23523 8449 23532 8483
rect 23480 8440 23532 8449
rect 26884 8440 26936 8492
rect 21088 8372 21140 8424
rect 21180 8372 21232 8424
rect 22192 8372 22244 8424
rect 22928 8372 22980 8424
rect 30380 8440 30432 8492
rect 31300 8440 31352 8492
rect 34244 8440 34296 8492
rect 19248 8304 19300 8356
rect 21548 8304 21600 8356
rect 21916 8304 21968 8356
rect 23756 8304 23808 8356
rect 29644 8372 29696 8424
rect 31116 8372 31168 8424
rect 19616 8236 19668 8288
rect 21364 8236 21416 8288
rect 23296 8279 23348 8288
rect 23296 8245 23305 8279
rect 23305 8245 23339 8279
rect 23339 8245 23348 8279
rect 23296 8236 23348 8245
rect 23388 8236 23440 8288
rect 25136 8236 25188 8288
rect 28356 8347 28408 8356
rect 28356 8313 28365 8347
rect 28365 8313 28399 8347
rect 28399 8313 28408 8347
rect 28356 8304 28408 8313
rect 29828 8236 29880 8288
rect 32404 8415 32456 8424
rect 32404 8381 32413 8415
rect 32413 8381 32447 8415
rect 32447 8381 32456 8415
rect 32404 8372 32456 8381
rect 32496 8372 32548 8424
rect 32772 8236 32824 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 7748 7939 7800 7948
rect 7748 7905 7757 7939
rect 7757 7905 7791 7939
rect 7791 7905 7800 7939
rect 7748 7896 7800 7905
rect 6920 7871 6972 7880
rect 6920 7837 6929 7871
rect 6929 7837 6963 7871
rect 6963 7837 6972 7871
rect 6920 7828 6972 7837
rect 8024 7828 8076 7880
rect 13544 8032 13596 8084
rect 12348 8007 12400 8016
rect 12348 7973 12357 8007
rect 12357 7973 12391 8007
rect 12391 7973 12400 8007
rect 12348 7964 12400 7973
rect 18052 8032 18104 8084
rect 19984 8075 20036 8084
rect 19984 8041 19993 8075
rect 19993 8041 20027 8075
rect 20027 8041 20036 8075
rect 19984 8032 20036 8041
rect 20260 8075 20312 8084
rect 20260 8041 20269 8075
rect 20269 8041 20303 8075
rect 20303 8041 20312 8075
rect 20260 8032 20312 8041
rect 19616 7964 19668 8016
rect 19708 7964 19760 8016
rect 12808 7939 12860 7948
rect 12808 7905 12817 7939
rect 12817 7905 12851 7939
rect 12851 7905 12860 7939
rect 12808 7896 12860 7905
rect 13452 7896 13504 7948
rect 9864 7828 9916 7880
rect 15108 7896 15160 7948
rect 13636 7828 13688 7880
rect 14004 7828 14056 7880
rect 14740 7828 14792 7880
rect 15016 7828 15068 7880
rect 17500 7896 17552 7948
rect 17684 7896 17736 7948
rect 16948 7828 17000 7880
rect 17316 7871 17368 7880
rect 17316 7837 17325 7871
rect 17325 7837 17359 7871
rect 17359 7837 17368 7871
rect 17316 7828 17368 7837
rect 17408 7871 17460 7880
rect 17408 7837 17418 7871
rect 17418 7837 17452 7871
rect 17452 7837 17460 7871
rect 17408 7828 17460 7837
rect 17868 7828 17920 7880
rect 15936 7760 15988 7812
rect 17592 7803 17644 7812
rect 17592 7769 17601 7803
rect 17601 7769 17635 7803
rect 17635 7769 17644 7803
rect 17592 7760 17644 7769
rect 19984 7896 20036 7948
rect 20444 7896 20496 7948
rect 21272 7939 21324 7948
rect 21272 7905 21281 7939
rect 21281 7905 21315 7939
rect 21315 7905 21324 7939
rect 21272 7896 21324 7905
rect 21916 8007 21968 8016
rect 21916 7973 21925 8007
rect 21925 7973 21959 8007
rect 21959 7973 21968 8007
rect 21916 7964 21968 7973
rect 22192 8075 22244 8084
rect 22192 8041 22201 8075
rect 22201 8041 22235 8075
rect 22235 8041 22244 8075
rect 22192 8032 22244 8041
rect 22928 8032 22980 8084
rect 23296 8032 23348 8084
rect 27436 8032 27488 8084
rect 20260 7828 20312 7880
rect 20352 7828 20404 7880
rect 7288 7735 7340 7744
rect 7288 7701 7297 7735
rect 7297 7701 7331 7735
rect 7331 7701 7340 7735
rect 7288 7692 7340 7701
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 8944 7692 8996 7701
rect 9588 7692 9640 7744
rect 13820 7692 13872 7744
rect 16488 7735 16540 7744
rect 16488 7701 16497 7735
rect 16497 7701 16531 7735
rect 16531 7701 16540 7735
rect 16488 7692 16540 7701
rect 17316 7692 17368 7744
rect 20720 7760 20772 7812
rect 19616 7692 19668 7744
rect 20812 7735 20864 7744
rect 20812 7701 20821 7735
rect 20821 7701 20855 7735
rect 20855 7701 20864 7735
rect 20812 7692 20864 7701
rect 28724 8032 28776 8084
rect 31300 8075 31352 8084
rect 31300 8041 31309 8075
rect 31309 8041 31343 8075
rect 31343 8041 31352 8075
rect 31300 8032 31352 8041
rect 32404 8032 32456 8084
rect 29920 7896 29972 7948
rect 31024 7896 31076 7948
rect 31116 7896 31168 7948
rect 22928 7828 22980 7880
rect 23020 7871 23072 7880
rect 23020 7837 23029 7871
rect 23029 7837 23063 7871
rect 23063 7837 23072 7871
rect 23020 7828 23072 7837
rect 23756 7828 23808 7880
rect 23848 7871 23900 7880
rect 23848 7837 23857 7871
rect 23857 7837 23891 7871
rect 23891 7837 23900 7871
rect 23848 7828 23900 7837
rect 27252 7828 27304 7880
rect 28356 7828 28408 7880
rect 33140 7896 33192 7948
rect 32496 7828 32548 7880
rect 34336 7828 34388 7880
rect 21824 7692 21876 7744
rect 22192 7692 22244 7744
rect 22468 7760 22520 7812
rect 23388 7692 23440 7744
rect 27160 7692 27212 7744
rect 29828 7803 29880 7812
rect 29828 7769 29837 7803
rect 29837 7769 29871 7803
rect 29871 7769 29880 7803
rect 29828 7760 29880 7769
rect 32588 7760 32640 7812
rect 34704 7760 34756 7812
rect 31576 7692 31628 7744
rect 32680 7735 32732 7744
rect 32680 7701 32689 7735
rect 32689 7701 32723 7735
rect 32723 7701 32732 7735
rect 32680 7692 32732 7701
rect 33048 7692 33100 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 8024 7488 8076 7540
rect 9864 7488 9916 7540
rect 10140 7488 10192 7540
rect 12716 7488 12768 7540
rect 13452 7488 13504 7540
rect 14004 7531 14056 7540
rect 14004 7497 14013 7531
rect 14013 7497 14047 7531
rect 14047 7497 14056 7531
rect 14004 7488 14056 7497
rect 14188 7531 14240 7540
rect 14188 7497 14197 7531
rect 14197 7497 14231 7531
rect 14231 7497 14240 7531
rect 14188 7488 14240 7497
rect 14464 7488 14516 7540
rect 15108 7531 15160 7540
rect 15108 7497 15117 7531
rect 15117 7497 15151 7531
rect 15151 7497 15160 7531
rect 15108 7488 15160 7497
rect 18420 7488 18472 7540
rect 1308 7352 1360 7404
rect 6920 7420 6972 7472
rect 7288 7352 7340 7404
rect 8944 7352 8996 7404
rect 13820 7420 13872 7472
rect 20628 7488 20680 7540
rect 21824 7531 21876 7540
rect 21824 7497 21833 7531
rect 21833 7497 21867 7531
rect 21867 7497 21876 7531
rect 21824 7488 21876 7497
rect 21916 7488 21968 7540
rect 22744 7488 22796 7540
rect 22928 7488 22980 7540
rect 23388 7488 23440 7540
rect 23664 7488 23716 7540
rect 10048 7352 10100 7404
rect 11520 7395 11572 7404
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 11612 7352 11664 7404
rect 14556 7352 14608 7404
rect 17684 7395 17736 7404
rect 17684 7361 17718 7395
rect 17718 7361 17736 7395
rect 17684 7352 17736 7361
rect 18880 7395 18932 7404
rect 18880 7361 18889 7395
rect 18889 7361 18923 7395
rect 18923 7361 18932 7395
rect 18880 7352 18932 7361
rect 20352 7352 20404 7404
rect 21548 7352 21600 7404
rect 23020 7420 23072 7472
rect 23848 7488 23900 7540
rect 24768 7488 24820 7540
rect 15108 7284 15160 7336
rect 15936 7284 15988 7336
rect 20444 7284 20496 7336
rect 22652 7284 22704 7336
rect 23112 7352 23164 7404
rect 24308 7352 24360 7404
rect 24492 7395 24544 7404
rect 24492 7361 24501 7395
rect 24501 7361 24535 7395
rect 24535 7361 24544 7395
rect 24492 7352 24544 7361
rect 24768 7395 24820 7404
rect 24768 7361 24777 7395
rect 24777 7361 24811 7395
rect 24811 7361 24820 7395
rect 24768 7352 24820 7361
rect 25228 7420 25280 7472
rect 25320 7395 25372 7404
rect 25320 7361 25329 7395
rect 25329 7361 25363 7395
rect 25363 7361 25372 7395
rect 25320 7352 25372 7361
rect 25412 7395 25464 7404
rect 25412 7361 25421 7395
rect 25421 7361 25455 7395
rect 25455 7361 25464 7395
rect 25412 7352 25464 7361
rect 25504 7395 25556 7404
rect 25504 7361 25513 7395
rect 25513 7361 25547 7395
rect 25547 7361 25556 7395
rect 25504 7352 25556 7361
rect 31576 7531 31628 7540
rect 31576 7497 31585 7531
rect 31585 7497 31619 7531
rect 31619 7497 31628 7531
rect 31576 7488 31628 7497
rect 31944 7531 31996 7540
rect 31944 7497 31953 7531
rect 31953 7497 31987 7531
rect 31987 7497 31996 7531
rect 31944 7488 31996 7497
rect 26056 7395 26108 7404
rect 26056 7361 26065 7395
rect 26065 7361 26099 7395
rect 26099 7361 26108 7395
rect 26056 7352 26108 7361
rect 26148 7395 26200 7404
rect 26148 7361 26157 7395
rect 26157 7361 26191 7395
rect 26191 7361 26200 7395
rect 26148 7352 26200 7361
rect 28724 7395 28776 7404
rect 28724 7361 28733 7395
rect 28733 7361 28767 7395
rect 28767 7361 28776 7395
rect 28724 7352 28776 7361
rect 1860 7216 1912 7268
rect 20628 7216 20680 7268
rect 25136 7327 25188 7336
rect 25136 7293 25145 7327
rect 25145 7293 25179 7327
rect 25179 7293 25188 7327
rect 25136 7284 25188 7293
rect 25320 7216 25372 7268
rect 30472 7352 30524 7404
rect 31300 7420 31352 7472
rect 32220 7395 32272 7404
rect 32220 7361 32229 7395
rect 32229 7361 32263 7395
rect 32263 7361 32272 7395
rect 32220 7352 32272 7361
rect 32588 7488 32640 7540
rect 32864 7488 32916 7540
rect 33140 7488 33192 7540
rect 32680 7352 32732 7404
rect 33140 7352 33192 7404
rect 31300 7327 31352 7336
rect 31300 7293 31309 7327
rect 31309 7293 31343 7327
rect 31343 7293 31352 7327
rect 31300 7284 31352 7293
rect 32772 7284 32824 7336
rect 33508 7327 33560 7336
rect 33508 7293 33517 7327
rect 33517 7293 33551 7327
rect 33551 7293 33560 7327
rect 33508 7284 33560 7293
rect 31852 7216 31904 7268
rect 21548 7191 21600 7200
rect 21548 7157 21557 7191
rect 21557 7157 21591 7191
rect 21591 7157 21600 7191
rect 21548 7148 21600 7157
rect 25228 7148 25280 7200
rect 29368 7191 29420 7200
rect 29368 7157 29377 7191
rect 29377 7157 29411 7191
rect 29411 7157 29420 7191
rect 29368 7148 29420 7157
rect 31116 7148 31168 7200
rect 33048 7148 33100 7200
rect 34244 7148 34296 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 10048 6987 10100 6996
rect 10048 6953 10057 6987
rect 10057 6953 10091 6987
rect 10091 6953 10100 6987
rect 10048 6944 10100 6953
rect 11612 6944 11664 6996
rect 17316 6987 17368 6996
rect 17316 6953 17325 6987
rect 17325 6953 17359 6987
rect 17359 6953 17368 6987
rect 17316 6944 17368 6953
rect 17684 6944 17736 6996
rect 20352 6944 20404 6996
rect 21272 6944 21324 6996
rect 22744 6944 22796 6996
rect 23664 6944 23716 6996
rect 25228 6944 25280 6996
rect 26056 6987 26108 6996
rect 26056 6953 26065 6987
rect 26065 6953 26099 6987
rect 26099 6953 26108 6987
rect 26056 6944 26108 6953
rect 26148 6944 26200 6996
rect 31852 6944 31904 6996
rect 25044 6876 25096 6928
rect 25320 6876 25372 6928
rect 9680 6808 9732 6860
rect 10140 6740 10192 6792
rect 11980 6851 12032 6860
rect 11980 6817 11989 6851
rect 11989 6817 12023 6851
rect 12023 6817 12032 6851
rect 11980 6808 12032 6817
rect 12440 6851 12492 6860
rect 12440 6817 12449 6851
rect 12449 6817 12483 6851
rect 12483 6817 12492 6851
rect 12440 6808 12492 6817
rect 15936 6851 15988 6860
rect 15936 6817 15945 6851
rect 15945 6817 15979 6851
rect 15979 6817 15988 6851
rect 15936 6808 15988 6817
rect 12716 6740 12768 6792
rect 16488 6740 16540 6792
rect 16948 6740 17000 6792
rect 18880 6808 18932 6860
rect 19708 6740 19760 6792
rect 23204 6808 23256 6860
rect 27804 6876 27856 6928
rect 28724 6876 28776 6928
rect 22284 6740 22336 6792
rect 22836 6740 22888 6792
rect 23388 6783 23440 6792
rect 23388 6749 23397 6783
rect 23397 6749 23431 6783
rect 23431 6749 23440 6783
rect 23388 6740 23440 6749
rect 23664 6783 23716 6792
rect 23664 6749 23673 6783
rect 23673 6749 23707 6783
rect 23707 6749 23716 6783
rect 23664 6740 23716 6749
rect 12440 6672 12492 6724
rect 14188 6672 14240 6724
rect 18420 6672 18472 6724
rect 20812 6672 20864 6724
rect 23480 6672 23532 6724
rect 24400 6783 24452 6792
rect 24400 6749 24409 6783
rect 24409 6749 24443 6783
rect 24443 6749 24452 6783
rect 24400 6740 24452 6749
rect 24768 6783 24820 6792
rect 24768 6749 24777 6783
rect 24777 6749 24811 6783
rect 24811 6749 24820 6783
rect 24768 6740 24820 6749
rect 25228 6740 25280 6792
rect 25964 6808 26016 6860
rect 27896 6808 27948 6860
rect 28816 6808 28868 6860
rect 30196 6808 30248 6860
rect 31668 6876 31720 6928
rect 31760 6876 31812 6928
rect 32404 6876 32456 6928
rect 33508 6944 33560 6996
rect 33048 6876 33100 6928
rect 31576 6808 31628 6860
rect 14648 6604 14700 6656
rect 21088 6604 21140 6656
rect 24584 6672 24636 6724
rect 24952 6672 25004 6724
rect 24492 6604 24544 6656
rect 26056 6672 26108 6724
rect 29000 6783 29052 6792
rect 29000 6749 29009 6783
rect 29009 6749 29043 6783
rect 29043 6749 29052 6783
rect 29000 6740 29052 6749
rect 29920 6783 29972 6792
rect 29920 6749 29929 6783
rect 29929 6749 29963 6783
rect 29963 6749 29972 6783
rect 29920 6740 29972 6749
rect 31116 6740 31168 6792
rect 31760 6740 31812 6792
rect 31852 6783 31904 6792
rect 31852 6749 31861 6783
rect 31861 6749 31895 6783
rect 31895 6749 31904 6783
rect 31852 6740 31904 6749
rect 31944 6783 31996 6792
rect 31944 6749 31953 6783
rect 31953 6749 31987 6783
rect 31987 6749 31996 6783
rect 33416 6808 33468 6860
rect 31944 6740 31996 6749
rect 32588 6783 32640 6792
rect 32588 6749 32597 6783
rect 32597 6749 32631 6783
rect 32631 6749 32640 6783
rect 32588 6740 32640 6749
rect 25320 6647 25372 6656
rect 25320 6613 25329 6647
rect 25329 6613 25363 6647
rect 25363 6613 25372 6647
rect 25320 6604 25372 6613
rect 25688 6647 25740 6656
rect 25688 6613 25697 6647
rect 25697 6613 25731 6647
rect 25731 6613 25740 6647
rect 25688 6604 25740 6613
rect 26884 6604 26936 6656
rect 27344 6604 27396 6656
rect 27896 6604 27948 6656
rect 30840 6604 30892 6656
rect 31392 6604 31444 6656
rect 31576 6604 31628 6656
rect 31944 6604 31996 6656
rect 32312 6672 32364 6724
rect 32404 6715 32456 6724
rect 32404 6681 32413 6715
rect 32413 6681 32447 6715
rect 32447 6681 32456 6715
rect 32404 6672 32456 6681
rect 32864 6740 32916 6792
rect 34060 6783 34112 6792
rect 34060 6749 34069 6783
rect 34069 6749 34103 6783
rect 34103 6749 34112 6783
rect 34060 6740 34112 6749
rect 34244 6783 34296 6792
rect 34244 6749 34253 6783
rect 34253 6749 34287 6783
rect 34287 6749 34296 6783
rect 34244 6740 34296 6749
rect 33416 6715 33468 6724
rect 33416 6681 33425 6715
rect 33425 6681 33459 6715
rect 33459 6681 33468 6715
rect 33416 6672 33468 6681
rect 34428 6740 34480 6792
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 14188 6443 14240 6452
rect 14188 6409 14197 6443
rect 14197 6409 14231 6443
rect 14231 6409 14240 6443
rect 14188 6400 14240 6409
rect 14556 6443 14608 6452
rect 14556 6409 14565 6443
rect 14565 6409 14599 6443
rect 14599 6409 14608 6443
rect 14556 6400 14608 6409
rect 14648 6443 14700 6452
rect 14648 6409 14657 6443
rect 14657 6409 14691 6443
rect 14691 6409 14700 6443
rect 14648 6400 14700 6409
rect 15016 6443 15068 6452
rect 15016 6409 15025 6443
rect 15025 6409 15059 6443
rect 15059 6409 15068 6443
rect 15016 6400 15068 6409
rect 23112 6400 23164 6452
rect 23756 6400 23808 6452
rect 24584 6400 24636 6452
rect 25320 6400 25372 6452
rect 26148 6400 26200 6452
rect 26240 6400 26292 6452
rect 28816 6443 28868 6452
rect 28816 6409 28825 6443
rect 28825 6409 28859 6443
rect 28859 6409 28868 6443
rect 28816 6400 28868 6409
rect 29460 6400 29512 6452
rect 31208 6400 31260 6452
rect 31300 6443 31352 6452
rect 31300 6409 31309 6443
rect 31309 6409 31343 6443
rect 31343 6409 31352 6443
rect 31300 6400 31352 6409
rect 32220 6400 32272 6452
rect 32312 6400 32364 6452
rect 33416 6443 33468 6452
rect 33416 6409 33425 6443
rect 33425 6409 33459 6443
rect 33459 6409 33468 6443
rect 33416 6400 33468 6409
rect 21088 6307 21140 6316
rect 21088 6273 21097 6307
rect 21097 6273 21131 6307
rect 21131 6273 21140 6307
rect 21088 6264 21140 6273
rect 15016 6196 15068 6248
rect 22284 6307 22336 6316
rect 22284 6273 22293 6307
rect 22293 6273 22327 6307
rect 22327 6273 22336 6307
rect 22284 6264 22336 6273
rect 23664 6264 23716 6316
rect 24492 6264 24544 6316
rect 24584 6307 24636 6316
rect 24584 6273 24593 6307
rect 24593 6273 24627 6307
rect 24627 6273 24636 6307
rect 24584 6264 24636 6273
rect 22468 6060 22520 6112
rect 23388 6239 23440 6248
rect 23388 6205 23397 6239
rect 23397 6205 23431 6239
rect 23431 6205 23440 6239
rect 23388 6196 23440 6205
rect 23848 6196 23900 6248
rect 25044 6264 25096 6316
rect 25136 6264 25188 6316
rect 24952 6196 25004 6248
rect 25688 6196 25740 6248
rect 25228 6128 25280 6180
rect 27804 6128 27856 6180
rect 29092 6332 29144 6384
rect 28816 6264 28868 6316
rect 29000 6264 29052 6316
rect 30012 6264 30064 6316
rect 29368 6196 29420 6248
rect 29736 6196 29788 6248
rect 29920 6239 29972 6248
rect 29920 6205 29929 6239
rect 29929 6205 29963 6239
rect 29963 6205 29972 6239
rect 29920 6196 29972 6205
rect 30748 6264 30800 6316
rect 31116 6264 31168 6316
rect 31484 6307 31536 6316
rect 31484 6273 31493 6307
rect 31493 6273 31527 6307
rect 31527 6273 31536 6307
rect 31484 6264 31536 6273
rect 31668 6307 31720 6316
rect 31668 6273 31677 6307
rect 31677 6273 31711 6307
rect 31711 6273 31720 6307
rect 31668 6264 31720 6273
rect 33048 6332 33100 6384
rect 30472 6239 30524 6248
rect 30472 6205 30481 6239
rect 30481 6205 30515 6239
rect 30515 6205 30524 6239
rect 30472 6196 30524 6205
rect 23664 6060 23716 6112
rect 23756 6060 23808 6112
rect 25044 6103 25096 6112
rect 25044 6069 25053 6103
rect 25053 6069 25087 6103
rect 25087 6069 25096 6103
rect 25044 6060 25096 6069
rect 26240 6060 26292 6112
rect 27436 6060 27488 6112
rect 29828 6128 29880 6180
rect 32864 6307 32916 6316
rect 32864 6273 32873 6307
rect 32873 6273 32907 6307
rect 32907 6273 32916 6307
rect 32864 6264 32916 6273
rect 34428 6264 34480 6316
rect 33048 6239 33100 6248
rect 33048 6205 33053 6239
rect 33053 6205 33087 6239
rect 33087 6205 33100 6239
rect 33048 6196 33100 6205
rect 31300 6060 31352 6112
rect 32496 6103 32548 6112
rect 32496 6069 32505 6103
rect 32505 6069 32539 6103
rect 32539 6069 32548 6103
rect 32496 6060 32548 6069
rect 33140 6171 33192 6180
rect 33140 6137 33149 6171
rect 33149 6137 33183 6171
rect 33183 6137 33192 6171
rect 33140 6128 33192 6137
rect 33232 6103 33284 6112
rect 33232 6069 33241 6103
rect 33241 6069 33275 6103
rect 33275 6069 33284 6103
rect 33232 6060 33284 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1860 5720 1912 5772
rect 23480 5856 23532 5908
rect 24400 5856 24452 5908
rect 25412 5856 25464 5908
rect 22192 5720 22244 5772
rect 22468 5720 22520 5772
rect 23388 5720 23440 5772
rect 23940 5763 23992 5772
rect 23940 5729 23949 5763
rect 23949 5729 23983 5763
rect 23983 5729 23992 5763
rect 23940 5720 23992 5729
rect 25044 5720 25096 5772
rect 23756 5695 23808 5704
rect 23756 5661 23765 5695
rect 23765 5661 23799 5695
rect 23799 5661 23808 5695
rect 23756 5652 23808 5661
rect 23112 5627 23164 5636
rect 23112 5593 23121 5627
rect 23121 5593 23155 5627
rect 23155 5593 23164 5627
rect 23112 5584 23164 5593
rect 23204 5584 23256 5636
rect 25228 5652 25280 5704
rect 27344 5720 27396 5772
rect 28816 5899 28868 5908
rect 28816 5865 28825 5899
rect 28825 5865 28859 5899
rect 28859 5865 28868 5899
rect 28816 5856 28868 5865
rect 29092 5899 29144 5908
rect 29092 5865 29101 5899
rect 29101 5865 29135 5899
rect 29135 5865 29144 5899
rect 29092 5856 29144 5865
rect 31392 5856 31444 5908
rect 32864 5856 32916 5908
rect 30288 5788 30340 5840
rect 30656 5788 30708 5840
rect 32036 5788 32088 5840
rect 33232 5788 33284 5840
rect 34152 5788 34204 5840
rect 29644 5652 29696 5704
rect 30748 5720 30800 5772
rect 30196 5695 30248 5704
rect 30196 5661 30205 5695
rect 30205 5661 30239 5695
rect 30239 5661 30248 5695
rect 30196 5652 30248 5661
rect 30380 5695 30432 5704
rect 30380 5661 30389 5695
rect 30389 5661 30423 5695
rect 30423 5661 30432 5695
rect 30380 5652 30432 5661
rect 27436 5584 27488 5636
rect 28724 5584 28776 5636
rect 29828 5627 29880 5636
rect 29828 5593 29837 5627
rect 29837 5593 29871 5627
rect 29871 5593 29880 5627
rect 29828 5584 29880 5593
rect 30012 5627 30064 5636
rect 30012 5593 30047 5627
rect 30047 5593 30064 5627
rect 30012 5584 30064 5593
rect 30196 5516 30248 5568
rect 30656 5695 30708 5704
rect 30656 5661 30665 5695
rect 30665 5661 30699 5695
rect 30699 5661 30708 5695
rect 30656 5652 30708 5661
rect 31024 5763 31076 5772
rect 31024 5729 31033 5763
rect 31033 5729 31067 5763
rect 31067 5729 31076 5763
rect 31024 5720 31076 5729
rect 31668 5720 31720 5772
rect 32588 5720 32640 5772
rect 31484 5652 31536 5704
rect 31300 5584 31352 5636
rect 32496 5516 32548 5568
rect 33140 5627 33192 5636
rect 33140 5593 33149 5627
rect 33149 5593 33183 5627
rect 33183 5593 33192 5627
rect 33140 5584 33192 5593
rect 33968 5584 34020 5636
rect 34428 5695 34480 5704
rect 34428 5661 34437 5695
rect 34437 5661 34471 5695
rect 34471 5661 34480 5695
rect 34428 5652 34480 5661
rect 34612 5516 34664 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 24032 5312 24084 5364
rect 24768 5312 24820 5364
rect 30380 5312 30432 5364
rect 33140 5312 33192 5364
rect 22284 5244 22336 5296
rect 1308 5176 1360 5228
rect 23572 5219 23624 5228
rect 23572 5185 23581 5219
rect 23581 5185 23615 5219
rect 23615 5185 23624 5219
rect 23572 5176 23624 5185
rect 24032 5219 24084 5228
rect 24032 5185 24041 5219
rect 24041 5185 24075 5219
rect 24075 5185 24084 5219
rect 24032 5176 24084 5185
rect 24860 5244 24912 5296
rect 26056 5244 26108 5296
rect 30472 5176 30524 5228
rect 33968 5219 34020 5228
rect 33968 5185 33977 5219
rect 33977 5185 34011 5219
rect 34011 5185 34020 5219
rect 33968 5176 34020 5185
rect 34152 5219 34204 5228
rect 34152 5185 34161 5219
rect 34161 5185 34195 5219
rect 34195 5185 34204 5219
rect 34152 5176 34204 5185
rect 34428 5219 34480 5228
rect 34428 5185 34437 5219
rect 34437 5185 34471 5219
rect 34471 5185 34480 5219
rect 34428 5176 34480 5185
rect 23296 5151 23348 5160
rect 23296 5117 23305 5151
rect 23305 5117 23339 5151
rect 23339 5117 23348 5151
rect 23296 5108 23348 5117
rect 23848 5108 23900 5160
rect 23940 5151 23992 5160
rect 23940 5117 23949 5151
rect 23949 5117 23983 5151
rect 23983 5117 23992 5151
rect 23940 5108 23992 5117
rect 30840 5108 30892 5160
rect 31024 5108 31076 5160
rect 35348 5108 35400 5160
rect 1860 5015 1912 5024
rect 1860 4981 1869 5015
rect 1869 4981 1903 5015
rect 1903 4981 1912 5015
rect 1860 4972 1912 4981
rect 30748 4972 30800 5024
rect 34060 4972 34112 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1860 4768 1912 4820
rect 33140 4768 33192 4820
rect 22284 4632 22336 4684
rect 23480 4632 23532 4684
rect 22744 4539 22796 4548
rect 22744 4505 22753 4539
rect 22753 4505 22787 4539
rect 22787 4505 22796 4539
rect 22744 4496 22796 4505
rect 29000 4632 29052 4684
rect 30288 4675 30340 4684
rect 30288 4641 30297 4675
rect 30297 4641 30331 4675
rect 30331 4641 30340 4675
rect 30288 4632 30340 4641
rect 30472 4632 30524 4684
rect 32404 4743 32456 4752
rect 32404 4709 32413 4743
rect 32413 4709 32447 4743
rect 32447 4709 32456 4743
rect 32404 4700 32456 4709
rect 30840 4564 30892 4616
rect 31392 4607 31444 4616
rect 31392 4573 31401 4607
rect 31401 4573 31435 4607
rect 31435 4573 31444 4607
rect 31392 4564 31444 4573
rect 32036 4607 32088 4616
rect 32036 4573 32045 4607
rect 32045 4573 32079 4607
rect 32079 4573 32088 4607
rect 32036 4564 32088 4573
rect 24400 4496 24452 4548
rect 29092 4496 29144 4548
rect 29920 4496 29972 4548
rect 33232 4496 33284 4548
rect 23572 4428 23624 4480
rect 31116 4428 31168 4480
rect 34428 4471 34480 4480
rect 34428 4437 34437 4471
rect 34437 4437 34471 4471
rect 34471 4437 34480 4471
rect 34428 4428 34480 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 22744 4224 22796 4276
rect 31116 4224 31168 4276
rect 32404 4224 32456 4276
rect 33232 4267 33284 4276
rect 33232 4233 33241 4267
rect 33241 4233 33275 4267
rect 33275 4233 33284 4267
rect 33232 4224 33284 4233
rect 23296 4088 23348 4140
rect 29000 4088 29052 4140
rect 29092 4131 29144 4140
rect 29092 4097 29101 4131
rect 29101 4097 29135 4131
rect 29135 4097 29144 4131
rect 29092 4088 29144 4097
rect 31300 4156 31352 4208
rect 31392 4156 31444 4208
rect 34428 4156 34480 4208
rect 23204 4020 23256 4072
rect 28724 4063 28776 4072
rect 28724 4029 28733 4063
rect 28733 4029 28767 4063
rect 28767 4029 28776 4063
rect 28724 4020 28776 4029
rect 29828 4020 29880 4072
rect 30104 4020 30156 4072
rect 29000 3927 29052 3936
rect 29000 3893 29009 3927
rect 29009 3893 29043 3927
rect 29043 3893 29052 3927
rect 29000 3884 29052 3893
rect 30840 3927 30892 3936
rect 30840 3893 30849 3927
rect 30849 3893 30883 3927
rect 30883 3893 30892 3927
rect 30840 3884 30892 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 29828 3723 29880 3732
rect 29828 3689 29837 3723
rect 29837 3689 29871 3723
rect 29871 3689 29880 3723
rect 29828 3680 29880 3689
rect 30104 3612 30156 3664
rect 29000 3544 29052 3596
rect 1308 3476 1360 3528
rect 30840 3476 30892 3528
rect 34060 3519 34112 3528
rect 34060 3485 34069 3519
rect 34069 3485 34103 3519
rect 34103 3485 34112 3519
rect 34060 3476 34112 3485
rect 34336 3451 34388 3460
rect 34336 3417 34345 3451
rect 34345 3417 34379 3451
rect 34379 3417 34388 3451
rect 34336 3408 34388 3417
rect 21548 3340 21600 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 1214 37360 1270 37369
rect 1214 37295 1270 37304
rect 1228 35766 1256 37295
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 1216 35760 1268 35766
rect 1216 35702 1268 35708
rect 19708 35760 19760 35766
rect 19708 35702 19760 35708
rect 1308 35692 1360 35698
rect 1308 35634 1360 35640
rect 10968 35692 11020 35698
rect 10968 35634 11020 35640
rect 1320 35465 1348 35634
rect 3608 35556 3660 35562
rect 3608 35498 3660 35504
rect 1306 35456 1362 35465
rect 1306 35391 1362 35400
rect 1320 35290 1348 35391
rect 1308 35284 1360 35290
rect 1308 35226 1360 35232
rect 3620 33998 3648 35498
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 9036 35284 9088 35290
rect 9036 35226 9088 35232
rect 7104 35080 7156 35086
rect 7104 35022 7156 35028
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4804 34060 4856 34066
rect 4804 34002 4856 34008
rect 1308 33992 1360 33998
rect 1308 33934 1360 33940
rect 3608 33992 3660 33998
rect 3608 33934 3660 33940
rect 1320 33561 1348 33934
rect 4068 33856 4120 33862
rect 4068 33798 4120 33804
rect 1306 33552 1362 33561
rect 1306 33487 1362 33496
rect 3976 32428 4028 32434
rect 3976 32370 4028 32376
rect 3424 32360 3476 32366
rect 3424 32302 3476 32308
rect 1400 31816 1452 31822
rect 1400 31758 1452 31764
rect 1412 31657 1440 31758
rect 1398 31648 1454 31657
rect 1398 31583 1454 31592
rect 1412 31482 1440 31583
rect 1400 31476 1452 31482
rect 1400 31418 1452 31424
rect 3436 31414 3464 32302
rect 3424 31408 3476 31414
rect 3424 31350 3476 31356
rect 3988 30938 4016 32370
rect 4080 31346 4108 33798
rect 4816 33454 4844 34002
rect 7116 33998 7144 35022
rect 8116 35012 8168 35018
rect 8116 34954 8168 34960
rect 8128 34746 8156 34954
rect 8760 34944 8812 34950
rect 8760 34886 8812 34892
rect 8116 34740 8168 34746
rect 8116 34682 8168 34688
rect 8772 34610 8800 34886
rect 9048 34746 9076 35226
rect 9588 35012 9640 35018
rect 9588 34954 9640 34960
rect 9600 34746 9628 34954
rect 10980 34950 11008 35634
rect 12072 35624 12124 35630
rect 12072 35566 12124 35572
rect 19064 35624 19116 35630
rect 19064 35566 19116 35572
rect 11336 35488 11388 35494
rect 11336 35430 11388 35436
rect 11348 35018 11376 35430
rect 11888 35080 11940 35086
rect 11888 35022 11940 35028
rect 11336 35012 11388 35018
rect 11336 34954 11388 34960
rect 11520 35012 11572 35018
rect 11520 34954 11572 34960
rect 10876 34944 10928 34950
rect 10876 34886 10928 34892
rect 10968 34944 11020 34950
rect 10968 34886 11020 34892
rect 10888 34746 10916 34886
rect 9036 34740 9088 34746
rect 9036 34682 9088 34688
rect 9588 34740 9640 34746
rect 9588 34682 9640 34688
rect 10600 34740 10652 34746
rect 10600 34682 10652 34688
rect 10876 34740 10928 34746
rect 10876 34682 10928 34688
rect 8760 34604 8812 34610
rect 8760 34546 8812 34552
rect 9048 34542 9076 34682
rect 10416 34672 10468 34678
rect 10416 34614 10468 34620
rect 9680 34604 9732 34610
rect 9680 34546 9732 34552
rect 9036 34536 9088 34542
rect 9036 34478 9088 34484
rect 9404 34536 9456 34542
rect 9404 34478 9456 34484
rect 5908 33992 5960 33998
rect 5908 33934 5960 33940
rect 7104 33992 7156 33998
rect 7104 33934 7156 33940
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 5448 33516 5500 33522
rect 5448 33458 5500 33464
rect 4804 33448 4856 33454
rect 4804 33390 4856 33396
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4816 32910 4844 33390
rect 5460 33114 5488 33458
rect 5448 33108 5500 33114
rect 5448 33050 5500 33056
rect 4804 32904 4856 32910
rect 4804 32846 4856 32852
rect 4816 32502 4844 32846
rect 5920 32774 5948 33934
rect 6368 33856 6420 33862
rect 6368 33798 6420 33804
rect 6380 33522 6408 33798
rect 7116 33590 7144 33934
rect 7380 33924 7432 33930
rect 7380 33866 7432 33872
rect 9036 33924 9088 33930
rect 9036 33866 9088 33872
rect 9220 33924 9272 33930
rect 9220 33866 9272 33872
rect 7392 33658 7420 33866
rect 7656 33856 7708 33862
rect 7656 33798 7708 33804
rect 7668 33658 7696 33798
rect 7380 33652 7432 33658
rect 7380 33594 7432 33600
rect 7656 33652 7708 33658
rect 7656 33594 7708 33600
rect 7104 33584 7156 33590
rect 7104 33526 7156 33532
rect 6368 33516 6420 33522
rect 6368 33458 6420 33464
rect 6184 33312 6236 33318
rect 6184 33254 6236 33260
rect 6196 32842 6224 33254
rect 6184 32836 6236 32842
rect 6184 32778 6236 32784
rect 5908 32768 5960 32774
rect 5908 32710 5960 32716
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 4804 32496 4856 32502
rect 4804 32438 4856 32444
rect 5920 32434 5948 32710
rect 5908 32428 5960 32434
rect 5908 32370 5960 32376
rect 4804 32224 4856 32230
rect 4804 32166 4856 32172
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4712 31884 4764 31890
rect 4712 31826 4764 31832
rect 4620 31816 4672 31822
rect 4620 31758 4672 31764
rect 4632 31346 4660 31758
rect 4068 31340 4120 31346
rect 4068 31282 4120 31288
rect 4620 31340 4672 31346
rect 4620 31282 4672 31288
rect 4632 31142 4660 31282
rect 4724 31278 4752 31826
rect 4712 31272 4764 31278
rect 4712 31214 4764 31220
rect 4620 31136 4672 31142
rect 4620 31078 4672 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 3976 30932 4028 30938
rect 3976 30874 4028 30880
rect 4620 30796 4672 30802
rect 4620 30738 4672 30744
rect 4632 30394 4660 30738
rect 4724 30734 4752 31214
rect 4816 30818 4844 32166
rect 5264 31816 5316 31822
rect 5264 31758 5316 31764
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 5172 31476 5224 31482
rect 5172 31418 5224 31424
rect 4816 30790 4936 30818
rect 4908 30734 4936 30790
rect 5184 30734 5212 31418
rect 4712 30728 4764 30734
rect 4712 30670 4764 30676
rect 4804 30728 4856 30734
rect 4804 30670 4856 30676
rect 4896 30728 4948 30734
rect 4896 30670 4948 30676
rect 5172 30728 5224 30734
rect 5172 30670 5224 30676
rect 4620 30388 4672 30394
rect 4620 30330 4672 30336
rect 1308 30252 1360 30258
rect 1308 30194 1360 30200
rect 3608 30252 3660 30258
rect 3608 30194 3660 30200
rect 1320 29753 1348 30194
rect 2872 30048 2924 30054
rect 2872 29990 2924 29996
rect 1306 29744 1362 29753
rect 1306 29679 1362 29688
rect 2228 29640 2280 29646
rect 2228 29582 2280 29588
rect 1308 28076 1360 28082
rect 1308 28018 1360 28024
rect 1320 27849 1348 28018
rect 1306 27840 1362 27849
rect 1306 27775 1362 27784
rect 2240 27538 2268 29582
rect 2884 28150 2912 29990
rect 3620 29850 3648 30194
rect 4620 30116 4672 30122
rect 4620 30058 4672 30064
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 3608 29844 3660 29850
rect 3608 29786 3660 29792
rect 3056 29572 3108 29578
rect 3056 29514 3108 29520
rect 3068 29306 3096 29514
rect 3620 29306 3648 29786
rect 4252 29572 4304 29578
rect 4252 29514 4304 29520
rect 4528 29572 4580 29578
rect 4528 29514 4580 29520
rect 4264 29306 4292 29514
rect 3056 29300 3108 29306
rect 3056 29242 3108 29248
rect 3608 29300 3660 29306
rect 3608 29242 3660 29248
rect 4252 29300 4304 29306
rect 4252 29242 4304 29248
rect 3700 29096 3752 29102
rect 3700 29038 3752 29044
rect 4540 29050 4568 29514
rect 4632 29510 4660 30058
rect 4620 29504 4672 29510
rect 4620 29446 4672 29452
rect 4632 29306 4660 29446
rect 4724 29306 4752 30670
rect 4816 30394 4844 30670
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 4804 30388 4856 30394
rect 4804 30330 4856 30336
rect 4896 30320 4948 30326
rect 4896 30262 4948 30268
rect 4804 30048 4856 30054
rect 4804 29990 4856 29996
rect 4620 29300 4672 29306
rect 4620 29242 4672 29248
rect 4712 29300 4764 29306
rect 4712 29242 4764 29248
rect 3712 28994 3740 29038
rect 3792 29028 3844 29034
rect 3712 28976 3792 28994
rect 4540 29022 4660 29050
rect 3712 28970 3844 28976
rect 3712 28966 3832 28970
rect 3424 28416 3476 28422
rect 3424 28358 3476 28364
rect 2872 28144 2924 28150
rect 2872 28086 2924 28092
rect 3436 28082 3464 28358
rect 3424 28076 3476 28082
rect 3424 28018 3476 28024
rect 2228 27532 2280 27538
rect 2228 27474 2280 27480
rect 2596 27396 2648 27402
rect 2596 27338 2648 27344
rect 3056 27396 3108 27402
rect 3056 27338 3108 27344
rect 2608 27130 2636 27338
rect 2596 27124 2648 27130
rect 2596 27066 2648 27072
rect 3068 26926 3096 27338
rect 3056 26920 3108 26926
rect 3056 26862 3108 26868
rect 3424 26920 3476 26926
rect 3424 26862 3476 26868
rect 1308 26376 1360 26382
rect 1308 26318 1360 26324
rect 1858 26344 1914 26353
rect 1320 25945 1348 26318
rect 1858 26279 1860 26288
rect 1912 26279 1914 26288
rect 1860 26250 1912 26256
rect 3068 26246 3096 26862
rect 3056 26240 3108 26246
rect 3056 26182 3108 26188
rect 1306 25936 1362 25945
rect 1306 25871 1362 25880
rect 3436 25362 3464 26862
rect 3712 26790 3740 28966
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4158 28112 4214 28121
rect 4158 28047 4160 28056
rect 4212 28047 4214 28056
rect 4252 28076 4304 28082
rect 4160 28018 4212 28024
rect 4252 28018 4304 28024
rect 3792 28008 3844 28014
rect 4264 27962 4292 28018
rect 3792 27950 3844 27956
rect 3804 26874 3832 27950
rect 4080 27934 4292 27962
rect 4080 27606 4108 27934
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4068 27600 4120 27606
rect 4120 27548 4200 27554
rect 4068 27542 4200 27548
rect 4080 27526 4200 27542
rect 3884 27328 3936 27334
rect 3884 27270 3936 27276
rect 3896 27062 3924 27270
rect 4172 27130 4200 27526
rect 4252 27532 4304 27538
rect 4252 27474 4304 27480
rect 4160 27124 4212 27130
rect 4160 27066 4212 27072
rect 4264 27062 4292 27474
rect 4632 27418 4660 29022
rect 4712 28144 4764 28150
rect 4712 28086 4764 28092
rect 4540 27390 4660 27418
rect 4344 27328 4396 27334
rect 4344 27270 4396 27276
rect 4356 27130 4384 27270
rect 4344 27124 4396 27130
rect 4344 27066 4396 27072
rect 3884 27056 3936 27062
rect 3884 26998 3936 27004
rect 4252 27056 4304 27062
rect 4252 26998 4304 27004
rect 3804 26846 3924 26874
rect 3700 26784 3752 26790
rect 3700 26726 3752 26732
rect 3712 26314 3740 26726
rect 3896 26382 3924 26846
rect 4540 26790 4568 27390
rect 4620 27328 4672 27334
rect 4620 27270 4672 27276
rect 4528 26784 4580 26790
rect 4528 26726 4580 26732
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 3884 26376 3936 26382
rect 3884 26318 3936 26324
rect 3700 26308 3752 26314
rect 3700 26250 3752 26256
rect 3608 25696 3660 25702
rect 3608 25638 3660 25644
rect 3424 25356 3476 25362
rect 3424 25298 3476 25304
rect 3436 24886 3464 25298
rect 3424 24880 3476 24886
rect 3424 24822 3476 24828
rect 1216 24200 1268 24206
rect 1216 24142 1268 24148
rect 1228 24041 1256 24142
rect 3436 24138 3464 24822
rect 3620 24818 3648 25638
rect 3608 24812 3660 24818
rect 3608 24754 3660 24760
rect 3424 24132 3476 24138
rect 3424 24074 3476 24080
rect 1214 24032 1270 24041
rect 1214 23967 1270 23976
rect 1308 22636 1360 22642
rect 1308 22578 1360 22584
rect 1320 22137 1348 22578
rect 1858 22536 1914 22545
rect 1858 22471 1860 22480
rect 1912 22471 1914 22480
rect 1860 22442 1912 22448
rect 1306 22128 1362 22137
rect 1306 22063 1362 22072
rect 3148 21888 3200 21894
rect 3148 21830 3200 21836
rect 3160 21622 3188 21830
rect 3148 21616 3200 21622
rect 3148 21558 3200 21564
rect 1308 20460 1360 20466
rect 1308 20402 1360 20408
rect 1320 20233 1348 20402
rect 1306 20224 1362 20233
rect 1306 20159 1362 20168
rect 3516 19440 3568 19446
rect 3516 19382 3568 19388
rect 3528 18766 3556 19382
rect 1308 18760 1360 18766
rect 1308 18702 1360 18708
rect 3516 18760 3568 18766
rect 3516 18702 3568 18708
rect 1320 18329 1348 18702
rect 1768 18624 1820 18630
rect 1768 18566 1820 18572
rect 1306 18320 1362 18329
rect 1306 18255 1362 18264
rect 1780 17882 1808 18566
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 3528 17134 3556 18702
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 1400 16584 1452 16590
rect 1400 16526 1452 16532
rect 1412 16425 1440 16526
rect 3528 16522 3556 17070
rect 2780 16516 2832 16522
rect 2780 16458 2832 16464
rect 3516 16516 3568 16522
rect 3516 16458 3568 16464
rect 1584 16448 1636 16454
rect 1398 16416 1454 16425
rect 1584 16390 1636 16396
rect 1398 16351 1454 16360
rect 1596 16114 1624 16390
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 2792 15502 2820 16458
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 1308 15020 1360 15026
rect 1308 14962 1360 14968
rect 1320 14521 1348 14962
rect 1306 14512 1362 14521
rect 1306 14447 1362 14456
rect 2792 13326 2820 15438
rect 2872 15428 2924 15434
rect 2872 15370 2924 15376
rect 2884 15162 2912 15370
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3252 15162 3280 15302
rect 3712 15162 3740 26250
rect 3896 24682 3924 26318
rect 4252 26240 4304 26246
rect 4252 26182 4304 26188
rect 4068 25968 4120 25974
rect 4068 25910 4120 25916
rect 4080 25378 4108 25910
rect 4264 25770 4292 26182
rect 4252 25764 4304 25770
rect 4252 25706 4304 25712
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4080 25350 4200 25378
rect 4172 24954 4200 25350
rect 4528 25220 4580 25226
rect 4528 25162 4580 25168
rect 4540 24954 4568 25162
rect 4160 24948 4212 24954
rect 4160 24890 4212 24896
rect 4528 24948 4580 24954
rect 4528 24890 4580 24896
rect 3884 24676 3936 24682
rect 3884 24618 3936 24624
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3884 24132 3936 24138
rect 3884 24074 3936 24080
rect 3896 23730 3924 24074
rect 3792 23724 3844 23730
rect 3792 23666 3844 23672
rect 3884 23724 3936 23730
rect 3936 23684 4108 23712
rect 3884 23666 3936 23672
rect 3804 22778 3832 23666
rect 4080 23304 4108 23684
rect 4632 23610 4660 27270
rect 4724 27130 4752 28086
rect 4816 28014 4844 29990
rect 4908 29578 4936 30262
rect 5276 29714 5304 31758
rect 6276 31340 6328 31346
rect 6276 31282 6328 31288
rect 5356 31272 5408 31278
rect 5356 31214 5408 31220
rect 5368 30326 5396 31214
rect 6288 30938 6316 31282
rect 6276 30932 6328 30938
rect 6276 30874 6328 30880
rect 5816 30592 5868 30598
rect 5816 30534 5868 30540
rect 5356 30320 5408 30326
rect 5356 30262 5408 30268
rect 5448 30252 5500 30258
rect 5448 30194 5500 30200
rect 5264 29708 5316 29714
rect 5264 29650 5316 29656
rect 4896 29572 4948 29578
rect 4896 29514 4948 29520
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 5276 29102 5304 29650
rect 5264 29096 5316 29102
rect 5264 29038 5316 29044
rect 5264 28416 5316 28422
rect 5264 28358 5316 28364
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 5276 28150 5304 28358
rect 5264 28144 5316 28150
rect 5264 28086 5316 28092
rect 4896 28076 4948 28082
rect 4896 28018 4948 28024
rect 4804 28008 4856 28014
rect 4804 27950 4856 27956
rect 4804 27872 4856 27878
rect 4804 27814 4856 27820
rect 4712 27124 4764 27130
rect 4712 27066 4764 27072
rect 4712 26784 4764 26790
rect 4712 26726 4764 26732
rect 4724 26042 4752 26726
rect 4712 26036 4764 26042
rect 4712 25978 4764 25984
rect 4724 25838 4752 25978
rect 4816 25906 4844 27814
rect 4908 27334 4936 28018
rect 5356 27872 5408 27878
rect 5356 27814 5408 27820
rect 4896 27328 4948 27334
rect 4896 27270 4948 27276
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4988 27056 5040 27062
rect 4988 26998 5040 27004
rect 5000 26790 5028 26998
rect 4988 26784 5040 26790
rect 4988 26726 5040 26732
rect 5000 26518 5028 26726
rect 4988 26512 5040 26518
rect 4988 26454 5040 26460
rect 5264 26512 5316 26518
rect 5264 26454 5316 26460
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 5276 26024 5304 26454
rect 4908 25996 5304 26024
rect 4804 25900 4856 25906
rect 4804 25842 4856 25848
rect 4712 25832 4764 25838
rect 4712 25774 4764 25780
rect 4908 25242 4936 25996
rect 5172 25900 5224 25906
rect 5172 25842 5224 25848
rect 5184 25498 5212 25842
rect 5172 25492 5224 25498
rect 5172 25434 5224 25440
rect 4816 25214 4936 25242
rect 5184 25242 5212 25434
rect 5184 25214 5304 25242
rect 4632 23582 4752 23610
rect 4620 23520 4672 23526
rect 4620 23462 4672 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4080 23276 4200 23304
rect 4172 23186 4200 23276
rect 4632 23202 4660 23462
rect 4160 23180 4212 23186
rect 4160 23122 4212 23128
rect 4540 23174 4660 23202
rect 4540 22778 4568 23174
rect 4620 23044 4672 23050
rect 4620 22986 4672 22992
rect 3792 22772 3844 22778
rect 3792 22714 3844 22720
rect 4528 22772 4580 22778
rect 4528 22714 4580 22720
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4528 22092 4580 22098
rect 4448 22052 4528 22080
rect 4160 21888 4212 21894
rect 4160 21830 4212 21836
rect 4172 21690 4200 21830
rect 4160 21684 4212 21690
rect 4160 21626 4212 21632
rect 4068 21548 4120 21554
rect 4068 21490 4120 21496
rect 4080 21146 4108 21490
rect 4448 21350 4476 22052
rect 4528 22034 4580 22040
rect 4528 21888 4580 21894
rect 4528 21830 4580 21836
rect 4540 21434 4568 21830
rect 4632 21622 4660 22986
rect 4724 22778 4752 23582
rect 4712 22772 4764 22778
rect 4712 22714 4764 22720
rect 4712 22568 4764 22574
rect 4712 22510 4764 22516
rect 4724 22030 4752 22510
rect 4816 22438 4844 25214
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 5276 24954 5304 25214
rect 5264 24948 5316 24954
rect 5264 24890 5316 24896
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 5276 23526 5304 23666
rect 5264 23520 5316 23526
rect 5264 23462 5316 23468
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5276 22710 5304 23462
rect 5264 22704 5316 22710
rect 5264 22646 5316 22652
rect 4804 22432 4856 22438
rect 4804 22374 4856 22380
rect 5264 22432 5316 22438
rect 5264 22374 5316 22380
rect 5172 22160 5224 22166
rect 5172 22102 5224 22108
rect 4712 22024 4764 22030
rect 5184 22012 5212 22102
rect 5276 22094 5304 22374
rect 5368 22234 5396 27814
rect 5460 26586 5488 30194
rect 5632 29164 5684 29170
rect 5632 29106 5684 29112
rect 5540 29096 5592 29102
rect 5540 29038 5592 29044
rect 5552 28558 5580 29038
rect 5540 28552 5592 28558
rect 5540 28494 5592 28500
rect 5448 26580 5500 26586
rect 5448 26522 5500 26528
rect 5460 25906 5488 26522
rect 5540 25968 5592 25974
rect 5540 25910 5592 25916
rect 5448 25900 5500 25906
rect 5448 25842 5500 25848
rect 5552 25786 5580 25910
rect 5460 25770 5580 25786
rect 5448 25764 5580 25770
rect 5500 25758 5580 25764
rect 5448 25706 5500 25712
rect 5460 24818 5488 25706
rect 5644 25702 5672 29106
rect 5722 26616 5778 26625
rect 5722 26551 5724 26560
rect 5776 26551 5778 26560
rect 5724 26522 5776 26528
rect 5736 26382 5764 26522
rect 5724 26376 5776 26382
rect 5724 26318 5776 26324
rect 5828 25838 5856 30534
rect 6276 29572 6328 29578
rect 6276 29514 6328 29520
rect 6184 29096 6236 29102
rect 6184 29038 6236 29044
rect 6196 28694 6224 29038
rect 6288 29034 6316 29514
rect 6380 29238 6408 33458
rect 7668 32978 7696 33594
rect 7840 33448 7892 33454
rect 7840 33390 7892 33396
rect 7012 32972 7064 32978
rect 7012 32914 7064 32920
rect 7656 32972 7708 32978
rect 7656 32914 7708 32920
rect 7748 32972 7800 32978
rect 7748 32914 7800 32920
rect 7024 32774 7052 32914
rect 7380 32904 7432 32910
rect 7760 32858 7788 32914
rect 7380 32846 7432 32852
rect 7012 32768 7064 32774
rect 7012 32710 7064 32716
rect 6736 32224 6788 32230
rect 6736 32166 6788 32172
rect 6748 30802 6776 32166
rect 6920 31476 6972 31482
rect 6920 31418 6972 31424
rect 6736 30796 6788 30802
rect 6788 30756 6868 30784
rect 6736 30738 6788 30744
rect 6736 29504 6788 29510
rect 6736 29446 6788 29452
rect 6748 29306 6776 29446
rect 6840 29306 6868 30756
rect 6932 30734 6960 31418
rect 6920 30728 6972 30734
rect 6920 30670 6972 30676
rect 6736 29300 6788 29306
rect 6736 29242 6788 29248
rect 6828 29300 6880 29306
rect 6828 29242 6880 29248
rect 6368 29232 6420 29238
rect 6368 29174 6420 29180
rect 6276 29028 6328 29034
rect 6276 28970 6328 28976
rect 6380 28762 6408 29174
rect 6368 28756 6420 28762
rect 6368 28698 6420 28704
rect 6184 28688 6236 28694
rect 6184 28630 6236 28636
rect 6092 28076 6144 28082
rect 6092 28018 6144 28024
rect 6104 27674 6132 28018
rect 6276 27872 6328 27878
rect 6276 27814 6328 27820
rect 6092 27668 6144 27674
rect 6092 27610 6144 27616
rect 6184 27464 6236 27470
rect 6184 27406 6236 27412
rect 6196 27062 6224 27406
rect 6288 27402 6316 27814
rect 6276 27396 6328 27402
rect 6276 27338 6328 27344
rect 6828 27396 6880 27402
rect 6828 27338 6880 27344
rect 6840 27130 6868 27338
rect 6828 27124 6880 27130
rect 6828 27066 6880 27072
rect 6184 27056 6236 27062
rect 6184 26998 6236 27004
rect 6552 26240 6604 26246
rect 6552 26182 6604 26188
rect 6564 25838 6592 26182
rect 5816 25832 5868 25838
rect 5816 25774 5868 25780
rect 6552 25832 6604 25838
rect 6552 25774 6604 25780
rect 5632 25696 5684 25702
rect 5632 25638 5684 25644
rect 6184 25696 6236 25702
rect 6184 25638 6236 25644
rect 5448 24812 5500 24818
rect 5448 24754 5500 24760
rect 5644 24750 5672 25638
rect 5632 24744 5684 24750
rect 5632 24686 5684 24692
rect 5448 24336 5500 24342
rect 5448 24278 5500 24284
rect 5460 23866 5488 24278
rect 6092 24064 6144 24070
rect 6092 24006 6144 24012
rect 5448 23860 5500 23866
rect 5448 23802 5500 23808
rect 5460 22574 5488 23802
rect 6104 23118 6132 24006
rect 6092 23112 6144 23118
rect 6092 23054 6144 23060
rect 5724 22636 5776 22642
rect 5724 22578 5776 22584
rect 5448 22568 5500 22574
rect 5448 22510 5500 22516
rect 5540 22568 5592 22574
rect 5540 22510 5592 22516
rect 5552 22250 5580 22510
rect 5736 22438 5764 22578
rect 5724 22432 5776 22438
rect 5724 22374 5776 22380
rect 5356 22228 5408 22234
rect 5356 22170 5408 22176
rect 5543 22222 5580 22250
rect 5632 22228 5684 22234
rect 5543 22094 5571 22222
rect 5632 22170 5684 22176
rect 5276 22066 5396 22094
rect 5543 22066 5580 22094
rect 5184 21984 5304 22012
rect 4712 21966 4764 21972
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4724 21690 4752 21830
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4712 21684 4764 21690
rect 4764 21644 4936 21672
rect 4712 21626 4764 21632
rect 4620 21616 4672 21622
rect 4672 21564 4844 21570
rect 4620 21558 4844 21564
rect 4632 21542 4844 21558
rect 4816 21486 4844 21542
rect 4804 21480 4856 21486
rect 4540 21406 4660 21434
rect 4804 21422 4856 21428
rect 4436 21344 4488 21350
rect 4436 21286 4488 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4068 21140 4120 21146
rect 4068 21082 4120 21088
rect 4632 20874 4660 21406
rect 4712 21344 4764 21350
rect 4712 21286 4764 21292
rect 4620 20868 4672 20874
rect 4620 20810 4672 20816
rect 3792 20256 3844 20262
rect 3792 20198 3844 20204
rect 3804 19854 3832 20198
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4160 19984 4212 19990
rect 4160 19926 4212 19932
rect 3792 19848 3844 19854
rect 3792 19790 3844 19796
rect 4172 19446 4200 19926
rect 4436 19848 4488 19854
rect 4436 19790 4488 19796
rect 4160 19440 4212 19446
rect 4160 19382 4212 19388
rect 4448 19310 4476 19790
rect 4724 19334 4752 21286
rect 4816 19922 4844 21422
rect 4908 20942 4936 21644
rect 4896 20936 4948 20942
rect 4896 20878 4948 20884
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4804 19916 4856 19922
rect 4804 19858 4856 19864
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4816 19468 5028 19496
rect 4816 19334 4844 19468
rect 5000 19378 5028 19468
rect 4436 19304 4488 19310
rect 4724 19306 4844 19334
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 4988 19372 5040 19378
rect 4988 19314 5040 19320
rect 4436 19246 4488 19252
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3884 18692 3936 18698
rect 3884 18634 3936 18640
rect 3896 18426 3924 18634
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 4172 18426 4200 18566
rect 3884 18420 3936 18426
rect 3884 18362 3936 18368
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 4080 16250 4108 17138
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16250 4660 17206
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4724 16046 4752 18158
rect 4816 17218 4844 19306
rect 4908 18630 4936 19314
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 5276 18222 5304 21984
rect 5368 21622 5396 22066
rect 5552 21962 5580 22066
rect 5540 21956 5592 21962
rect 5540 21898 5592 21904
rect 5644 21842 5672 22170
rect 5552 21814 5672 21842
rect 5356 21616 5408 21622
rect 5356 21558 5408 21564
rect 5368 19938 5396 21558
rect 5552 20262 5580 21814
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 5368 19910 5488 19938
rect 5460 19854 5488 19910
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5356 19780 5408 19786
rect 5356 19722 5408 19728
rect 5368 19514 5396 19722
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5460 19310 5488 19450
rect 5448 19304 5500 19310
rect 5448 19246 5500 19252
rect 5356 19236 5408 19242
rect 5356 19178 5408 19184
rect 5368 18630 5396 19178
rect 5460 18970 5488 19246
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5000 17218 5028 17274
rect 4816 17190 5028 17218
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 3700 15156 3752 15162
rect 3700 15098 3752 15104
rect 3712 14958 3740 15098
rect 4080 15094 4108 15846
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4160 15428 4212 15434
rect 4160 15370 4212 15376
rect 4172 15162 4200 15370
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4632 15162 4660 15302
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 3712 14822 3740 14894
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3436 13938 3464 14554
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2884 12986 2912 13874
rect 3700 13728 3752 13734
rect 4172 13716 4200 13874
rect 3700 13670 3752 13676
rect 4080 13688 4200 13716
rect 2964 13252 3016 13258
rect 2964 13194 3016 13200
rect 2976 12986 3004 13194
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 3712 12850 3740 13670
rect 4080 13530 4108 13688
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4068 13524 4120 13530
rect 4120 13484 4200 13512
rect 4068 13466 4120 13472
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 4080 12986 4108 13194
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 4172 12918 4200 13484
rect 4632 13190 4660 13874
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4356 12986 4384 13126
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 1308 12844 1360 12850
rect 1308 12786 1360 12792
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 1320 12617 1348 12786
rect 4724 12782 4752 15982
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4816 12628 4844 14758
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5276 13938 5304 17274
rect 5368 16794 5396 18566
rect 5460 18426 5488 18906
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5552 16946 5580 20198
rect 5736 17066 5764 22374
rect 6196 22234 6224 25638
rect 6368 25220 6420 25226
rect 6368 25162 6420 25168
rect 6380 24954 6408 25162
rect 6368 24948 6420 24954
rect 6368 24890 6420 24896
rect 6460 24064 6512 24070
rect 6460 24006 6512 24012
rect 6472 23254 6500 24006
rect 6460 23248 6512 23254
rect 6460 23190 6512 23196
rect 6184 22228 6236 22234
rect 6184 22170 6236 22176
rect 6460 21616 6512 21622
rect 6460 21558 6512 21564
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 5828 21146 5856 21490
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 5816 21140 5868 21146
rect 5816 21082 5868 21088
rect 6196 20942 6224 21286
rect 6472 21078 6500 21558
rect 6460 21072 6512 21078
rect 6460 21014 6512 21020
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 6184 20936 6236 20942
rect 6184 20878 6236 20884
rect 6380 20806 6408 20946
rect 6368 20800 6420 20806
rect 6288 20748 6368 20754
rect 6288 20742 6420 20748
rect 6288 20726 6408 20742
rect 6000 19780 6052 19786
rect 6000 19722 6052 19728
rect 6012 19310 6040 19722
rect 6184 19712 6236 19718
rect 6184 19654 6236 19660
rect 6196 19446 6224 19654
rect 6184 19440 6236 19446
rect 6184 19382 6236 19388
rect 6000 19304 6052 19310
rect 6000 19246 6052 19252
rect 6012 18358 6040 19246
rect 6000 18352 6052 18358
rect 6000 18294 6052 18300
rect 5724 17060 5776 17066
rect 5724 17002 5776 17008
rect 5460 16918 5580 16946
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5368 16114 5396 16594
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5460 15994 5488 16918
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5368 15966 5488 15994
rect 5368 15434 5396 15966
rect 5552 15858 5580 16730
rect 5460 15830 5580 15858
rect 5460 15570 5488 15830
rect 6288 15570 6316 20726
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 6380 16590 6408 16934
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 5356 15428 5408 15434
rect 5356 15370 5408 15376
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 5368 14822 5396 14894
rect 5460 14822 5488 15506
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5552 15366 5580 15438
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 5276 12866 5304 13874
rect 1306 12608 1362 12617
rect 1306 12543 1362 12552
rect 4724 12600 4844 12628
rect 5092 12838 5304 12866
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3240 11824 3292 11830
rect 3240 11766 3292 11772
rect 1308 11144 1360 11150
rect 1308 11086 1360 11092
rect 1320 10713 1348 11086
rect 3148 11076 3200 11082
rect 3148 11018 3200 11024
rect 3160 10713 3188 11018
rect 1306 10704 1362 10713
rect 1306 10639 1362 10648
rect 3146 10704 3202 10713
rect 3252 10674 3280 11766
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 3712 11354 3740 11698
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4264 10810 4292 11154
rect 4632 11150 4660 11494
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 3146 10639 3202 10648
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3620 10266 3648 10746
rect 4356 10690 4384 10950
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4264 10662 4384 10690
rect 4172 10554 4200 10610
rect 4264 10606 4292 10662
rect 4632 10606 4660 11086
rect 4080 10526 4200 10554
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 4080 10146 4108 10526
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4724 10198 4752 12600
rect 5092 12434 5120 12838
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 4816 12406 5120 12434
rect 4816 10538 4844 12406
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4908 11354 4936 11698
rect 5276 11642 5304 12718
rect 5368 12646 5396 14758
rect 5460 14006 5488 14758
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5448 14000 5500 14006
rect 5448 13942 5500 13948
rect 5552 13394 5580 14214
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5184 11614 5304 11642
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 5080 11280 5132 11286
rect 5080 11222 5132 11228
rect 5092 11121 5120 11222
rect 5078 11112 5134 11121
rect 5078 11047 5080 11056
rect 5132 11047 5134 11056
rect 5080 11018 5132 11024
rect 5184 11014 5212 11614
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 5276 11150 5304 11494
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4712 10192 4764 10198
rect 4080 10118 4200 10146
rect 4712 10134 4764 10140
rect 4172 10010 4200 10118
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4252 10056 4304 10062
rect 4172 10004 4252 10010
rect 4172 9998 4304 10004
rect 4172 9982 4292 9998
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3804 9654 3832 9862
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3896 8974 3924 9454
rect 3988 9382 4016 9522
rect 4264 9518 4292 9982
rect 4356 9722 4384 10066
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 1308 8968 1360 8974
rect 1308 8910 1360 8916
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 1320 8809 1348 8910
rect 1306 8800 1362 8809
rect 1306 8735 1362 8744
rect 3896 8498 3924 8910
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3988 8362 4016 9318
rect 4080 8974 4108 9386
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4632 8634 4660 9522
rect 4724 9178 4752 9998
rect 4816 9994 4844 10474
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4908 10266 4936 10406
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 5092 10062 5120 10746
rect 5276 10742 5304 11086
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5368 10554 5396 12582
rect 5552 12238 5580 13330
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 11830 5580 12174
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5276 10526 5396 10554
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4804 9988 4856 9994
rect 4804 9930 4856 9936
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 5276 8430 5304 10526
rect 5460 10010 5488 10950
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5368 9982 5488 10010
rect 5368 9625 5396 9982
rect 5552 9738 5580 10406
rect 5644 10266 5672 15302
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6380 14550 6408 14758
rect 6368 14544 6420 14550
rect 6368 14486 6420 14492
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 6380 14074 6408 14282
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6288 12918 6316 14010
rect 6368 13252 6420 13258
rect 6368 13194 6420 13200
rect 6380 12986 6408 13194
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 6472 12714 6500 16390
rect 6460 12708 6512 12714
rect 6460 12650 6512 12656
rect 6472 12170 6500 12650
rect 6564 12434 6592 25774
rect 6736 25152 6788 25158
rect 6736 25094 6788 25100
rect 6748 24954 6776 25094
rect 6736 24948 6788 24954
rect 6736 24890 6788 24896
rect 6644 24064 6696 24070
rect 6644 24006 6696 24012
rect 6656 23866 6684 24006
rect 6644 23860 6696 23866
rect 6644 23802 6696 23808
rect 7024 22094 7052 32710
rect 7196 32224 7248 32230
rect 7196 32166 7248 32172
rect 7104 32020 7156 32026
rect 7104 31962 7156 31968
rect 7116 31754 7144 31962
rect 7208 31822 7236 32166
rect 7392 32026 7420 32846
rect 7668 32842 7788 32858
rect 7656 32836 7788 32842
rect 7708 32830 7788 32836
rect 7656 32778 7708 32784
rect 7380 32020 7432 32026
rect 7380 31962 7432 31968
rect 7288 31884 7340 31890
rect 7288 31826 7340 31832
rect 7196 31816 7248 31822
rect 7196 31758 7248 31764
rect 7104 31748 7156 31754
rect 7104 31690 7156 31696
rect 7300 31414 7328 31826
rect 7472 31816 7524 31822
rect 7472 31758 7524 31764
rect 7288 31408 7340 31414
rect 7288 31350 7340 31356
rect 7196 27940 7248 27946
rect 7196 27882 7248 27888
rect 7208 27538 7236 27882
rect 7196 27532 7248 27538
rect 7196 27474 7248 27480
rect 7208 26994 7236 27474
rect 7196 26988 7248 26994
rect 7196 26930 7248 26936
rect 7300 26976 7328 31350
rect 7484 30666 7512 31758
rect 7564 31680 7616 31686
rect 7564 31622 7616 31628
rect 7576 30938 7604 31622
rect 7564 30932 7616 30938
rect 7564 30874 7616 30880
rect 7472 30660 7524 30666
rect 7472 30602 7524 30608
rect 7380 29572 7432 29578
rect 7380 29514 7432 29520
rect 7392 29306 7420 29514
rect 7380 29300 7432 29306
rect 7380 29242 7432 29248
rect 7484 28994 7512 30602
rect 7484 28966 7604 28994
rect 7576 28082 7604 28966
rect 7472 28076 7524 28082
rect 7472 28018 7524 28024
rect 7564 28076 7616 28082
rect 7564 28018 7616 28024
rect 7484 27674 7512 28018
rect 7472 27668 7524 27674
rect 7472 27610 7524 27616
rect 7484 27130 7512 27610
rect 7472 27124 7524 27130
rect 7472 27066 7524 27072
rect 7380 26988 7432 26994
rect 7300 26948 7380 26976
rect 7300 25906 7328 26948
rect 7380 26930 7432 26936
rect 7576 25922 7604 28018
rect 7668 27554 7696 32778
rect 7852 32774 7880 33390
rect 7840 32768 7892 32774
rect 7840 32710 7892 32716
rect 7852 32570 7880 32710
rect 7840 32564 7892 32570
rect 7840 32506 7892 32512
rect 9048 32502 9076 33866
rect 9232 33658 9260 33866
rect 9220 33652 9272 33658
rect 9220 33594 9272 33600
rect 9220 33380 9272 33386
rect 9220 33322 9272 33328
rect 9128 32564 9180 32570
rect 9128 32506 9180 32512
rect 8208 32496 8260 32502
rect 8208 32438 8260 32444
rect 9036 32496 9088 32502
rect 9036 32438 9088 32444
rect 8220 31890 8248 32438
rect 8852 32020 8904 32026
rect 8852 31962 8904 31968
rect 8208 31884 8260 31890
rect 8208 31826 8260 31832
rect 8116 31816 8168 31822
rect 8116 31758 8168 31764
rect 8128 31482 8156 31758
rect 8116 31476 8168 31482
rect 8116 31418 8168 31424
rect 8220 31346 8248 31826
rect 8760 31816 8812 31822
rect 8760 31758 8812 31764
rect 8208 31340 8260 31346
rect 8208 31282 8260 31288
rect 7748 29504 7800 29510
rect 7748 29446 7800 29452
rect 7760 29306 7788 29446
rect 7748 29300 7800 29306
rect 7748 29242 7800 29248
rect 8220 29238 8248 31282
rect 8772 29850 8800 31758
rect 8760 29844 8812 29850
rect 8760 29786 8812 29792
rect 8576 29640 8628 29646
rect 8576 29582 8628 29588
rect 8208 29232 8260 29238
rect 8208 29174 8260 29180
rect 8208 28552 8260 28558
rect 8208 28494 8260 28500
rect 7668 27526 7788 27554
rect 8220 27538 8248 28494
rect 8300 27872 8352 27878
rect 8588 27826 8616 29582
rect 8668 28960 8720 28966
rect 8668 28902 8720 28908
rect 8300 27814 8352 27820
rect 7760 26246 7788 27526
rect 8208 27532 8260 27538
rect 8208 27474 8260 27480
rect 8312 27470 8340 27814
rect 8496 27798 8616 27826
rect 8300 27464 8352 27470
rect 8300 27406 8352 27412
rect 8024 27328 8076 27334
rect 8024 27270 8076 27276
rect 8036 26994 8064 27270
rect 8024 26988 8076 26994
rect 8024 26930 8076 26936
rect 7748 26240 7800 26246
rect 7748 26182 7800 26188
rect 7288 25900 7340 25906
rect 7576 25894 7696 25922
rect 7288 25842 7340 25848
rect 7300 24750 7328 25842
rect 7668 25702 7696 25894
rect 8208 25900 8260 25906
rect 8208 25842 8260 25848
rect 7564 25696 7616 25702
rect 7564 25638 7616 25644
rect 7656 25696 7708 25702
rect 7656 25638 7708 25644
rect 7576 25294 7604 25638
rect 8220 25498 8248 25842
rect 8312 25838 8340 27406
rect 8300 25832 8352 25838
rect 8300 25774 8352 25780
rect 8208 25492 8260 25498
rect 8208 25434 8260 25440
rect 7564 25288 7616 25294
rect 7564 25230 7616 25236
rect 8312 25158 8340 25774
rect 8300 25152 8352 25158
rect 8300 25094 8352 25100
rect 7288 24744 7340 24750
rect 7288 24686 7340 24692
rect 8300 24132 8352 24138
rect 8300 24074 8352 24080
rect 8312 23730 8340 24074
rect 7196 23724 7248 23730
rect 7196 23666 7248 23672
rect 8300 23724 8352 23730
rect 8300 23666 8352 23672
rect 7208 23254 7236 23666
rect 7656 23588 7708 23594
rect 7656 23530 7708 23536
rect 8208 23588 8260 23594
rect 8208 23530 8260 23536
rect 7196 23248 7248 23254
rect 7196 23190 7248 23196
rect 7668 23186 7696 23530
rect 8024 23520 8076 23526
rect 8024 23462 8076 23468
rect 8036 23254 8064 23462
rect 8024 23248 8076 23254
rect 8024 23190 8076 23196
rect 8116 23248 8168 23254
rect 8116 23190 8168 23196
rect 7656 23180 7708 23186
rect 7656 23122 7708 23128
rect 7748 23180 7800 23186
rect 7748 23122 7800 23128
rect 7760 22778 7788 23122
rect 7840 23112 7892 23118
rect 7840 23054 7892 23060
rect 7748 22772 7800 22778
rect 7748 22714 7800 22720
rect 7024 22066 7144 22094
rect 6644 19712 6696 19718
rect 6644 19654 6696 19660
rect 6656 19446 6684 19654
rect 6644 19440 6696 19446
rect 6644 19382 6696 19388
rect 7012 19440 7064 19446
rect 7012 19382 7064 19388
rect 7024 18970 7052 19382
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 7024 18766 7052 18906
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 7116 18426 7144 22066
rect 7472 21344 7524 21350
rect 7472 21286 7524 21292
rect 7196 21140 7248 21146
rect 7196 21082 7248 21088
rect 7104 18420 7156 18426
rect 7104 18362 7156 18368
rect 7208 17814 7236 21082
rect 7484 20942 7512 21286
rect 7852 21146 7880 23054
rect 8128 22642 8156 23190
rect 8220 23066 8248 23530
rect 8220 23038 8340 23066
rect 8312 22642 8340 23038
rect 8116 22636 8168 22642
rect 8116 22578 8168 22584
rect 8300 22636 8352 22642
rect 8300 22578 8352 22584
rect 8312 21690 8340 22578
rect 8496 22094 8524 27798
rect 8576 26240 8628 26246
rect 8576 26182 8628 26188
rect 8588 25906 8616 26182
rect 8576 25900 8628 25906
rect 8576 25842 8628 25848
rect 8404 22066 8524 22094
rect 8680 22094 8708 28902
rect 8864 27878 8892 31962
rect 9140 31822 9168 32506
rect 9128 31816 9180 31822
rect 9128 31758 9180 31764
rect 9232 30326 9260 33322
rect 9416 32434 9444 34478
rect 9692 33522 9720 34546
rect 10428 34542 10456 34614
rect 10416 34536 10468 34542
rect 10416 34478 10468 34484
rect 10324 34468 10376 34474
rect 10324 34410 10376 34416
rect 10232 33992 10284 33998
rect 9770 33960 9826 33969
rect 10232 33934 10284 33940
rect 9770 33895 9826 33904
rect 9680 33516 9732 33522
rect 9680 33458 9732 33464
rect 9784 33454 9812 33895
rect 9956 33856 10008 33862
rect 9956 33798 10008 33804
rect 9862 33688 9918 33697
rect 9862 33623 9918 33632
rect 9876 33590 9904 33623
rect 9968 33590 9996 33798
rect 10244 33658 10272 33934
rect 10232 33652 10284 33658
rect 10232 33594 10284 33600
rect 9864 33584 9916 33590
rect 9864 33526 9916 33532
rect 9956 33584 10008 33590
rect 9956 33526 10008 33532
rect 9772 33448 9824 33454
rect 9772 33390 9824 33396
rect 9588 33108 9640 33114
rect 9588 33050 9640 33056
rect 9404 32428 9456 32434
rect 9324 32388 9404 32416
rect 9324 32026 9352 32388
rect 9404 32370 9456 32376
rect 9496 32360 9548 32366
rect 9496 32302 9548 32308
rect 9312 32020 9364 32026
rect 9312 31962 9364 31968
rect 9508 31958 9536 32302
rect 9600 32026 9628 33050
rect 9784 32978 9812 33390
rect 9772 32972 9824 32978
rect 9772 32914 9824 32920
rect 9772 32836 9824 32842
rect 9772 32778 9824 32784
rect 9784 32570 9812 32778
rect 9772 32564 9824 32570
rect 9772 32506 9824 32512
rect 9876 32026 9904 33526
rect 9968 33386 9996 33526
rect 10048 33516 10100 33522
rect 10048 33458 10100 33464
rect 10060 33386 10088 33458
rect 9956 33380 10008 33386
rect 9956 33322 10008 33328
rect 10048 33380 10100 33386
rect 10048 33322 10100 33328
rect 9956 32972 10008 32978
rect 9956 32914 10008 32920
rect 9588 32020 9640 32026
rect 9588 31962 9640 31968
rect 9864 32020 9916 32026
rect 9864 31962 9916 31968
rect 9496 31952 9548 31958
rect 9496 31894 9548 31900
rect 9312 31816 9364 31822
rect 9312 31758 9364 31764
rect 9404 31816 9456 31822
rect 9404 31758 9456 31764
rect 9508 31770 9536 31894
rect 9876 31822 9904 31962
rect 9864 31816 9916 31822
rect 9324 31482 9352 31758
rect 9312 31476 9364 31482
rect 9312 31418 9364 31424
rect 9324 31346 9352 31418
rect 9312 31340 9364 31346
rect 9312 31282 9364 31288
rect 9220 30320 9272 30326
rect 9220 30262 9272 30268
rect 9312 30184 9364 30190
rect 9416 30172 9444 31758
rect 9508 31754 9674 31770
rect 9864 31758 9916 31764
rect 9508 31742 9720 31754
rect 9646 31726 9720 31742
rect 9692 31482 9720 31726
rect 9680 31476 9732 31482
rect 9680 31418 9732 31424
rect 9680 31204 9732 31210
rect 9680 31146 9732 31152
rect 9364 30144 9444 30172
rect 9588 30184 9640 30190
rect 9312 30126 9364 30132
rect 9588 30126 9640 30132
rect 9036 30116 9088 30122
rect 9036 30058 9088 30064
rect 8944 30048 8996 30054
rect 8944 29990 8996 29996
rect 8956 29170 8984 29990
rect 9048 29646 9076 30058
rect 9600 30054 9628 30126
rect 9588 30048 9640 30054
rect 9588 29990 9640 29996
rect 9600 29730 9628 29990
rect 9508 29702 9628 29730
rect 9036 29640 9088 29646
rect 9036 29582 9088 29588
rect 8944 29164 8996 29170
rect 8944 29106 8996 29112
rect 8942 28112 8998 28121
rect 8942 28047 8998 28056
rect 8852 27872 8904 27878
rect 8852 27814 8904 27820
rect 8956 26926 8984 28047
rect 9036 27940 9088 27946
rect 9036 27882 9088 27888
rect 9048 27470 9076 27882
rect 9128 27532 9180 27538
rect 9128 27474 9180 27480
rect 9036 27464 9088 27470
rect 9036 27406 9088 27412
rect 9036 26988 9088 26994
rect 9036 26930 9088 26936
rect 8944 26920 8996 26926
rect 8944 26862 8996 26868
rect 8760 25696 8812 25702
rect 8760 25638 8812 25644
rect 8852 25696 8904 25702
rect 8852 25638 8904 25644
rect 8772 25362 8800 25638
rect 8760 25356 8812 25362
rect 8760 25298 8812 25304
rect 8864 24886 8892 25638
rect 8852 24880 8904 24886
rect 8852 24822 8904 24828
rect 9048 24698 9076 26930
rect 9140 26858 9168 27474
rect 9220 27464 9272 27470
rect 9220 27406 9272 27412
rect 9232 27130 9260 27406
rect 9220 27124 9272 27130
rect 9220 27066 9272 27072
rect 9128 26852 9180 26858
rect 9128 26794 9180 26800
rect 9508 26518 9536 29702
rect 9588 29640 9640 29646
rect 9588 29582 9640 29588
rect 9600 29238 9628 29582
rect 9692 29306 9720 31146
rect 9772 30252 9824 30258
rect 9772 30194 9824 30200
rect 9784 29306 9812 30194
rect 9680 29300 9732 29306
rect 9680 29242 9732 29248
rect 9772 29300 9824 29306
rect 9772 29242 9824 29248
rect 9588 29232 9640 29238
rect 9588 29174 9640 29180
rect 9588 27464 9640 27470
rect 9588 27406 9640 27412
rect 9600 27062 9628 27406
rect 9772 27328 9824 27334
rect 9876 27316 9904 31758
rect 9968 28014 9996 32914
rect 10060 28218 10088 33322
rect 10336 30682 10364 34410
rect 10428 31142 10456 34478
rect 10612 33998 10640 34682
rect 10600 33992 10652 33998
rect 10980 33946 11008 34886
rect 11532 34542 11560 34954
rect 11520 34536 11572 34542
rect 11520 34478 11572 34484
rect 11610 34504 11666 34513
rect 10600 33934 10652 33940
rect 10888 33930 11008 33946
rect 10876 33924 11008 33930
rect 10928 33918 11008 33924
rect 10876 33866 10928 33872
rect 11152 33856 11204 33862
rect 11152 33798 11204 33804
rect 10506 33688 10562 33697
rect 10506 33623 10508 33632
rect 10560 33623 10562 33632
rect 10508 33594 10560 33600
rect 10508 32904 10560 32910
rect 10508 32846 10560 32852
rect 10520 32434 10548 32846
rect 10784 32564 10836 32570
rect 10784 32506 10836 32512
rect 10508 32428 10560 32434
rect 10508 32370 10560 32376
rect 10692 31680 10744 31686
rect 10692 31622 10744 31628
rect 10416 31136 10468 31142
rect 10416 31078 10468 31084
rect 10244 30654 10364 30682
rect 10244 30308 10272 30654
rect 10428 30598 10456 31078
rect 10324 30592 10376 30598
rect 10324 30534 10376 30540
rect 10416 30592 10468 30598
rect 10416 30534 10468 30540
rect 10336 30410 10364 30534
rect 10336 30382 10456 30410
rect 10244 30280 10364 30308
rect 10232 30184 10284 30190
rect 10232 30126 10284 30132
rect 10140 29572 10192 29578
rect 10140 29514 10192 29520
rect 10152 29306 10180 29514
rect 10140 29300 10192 29306
rect 10140 29242 10192 29248
rect 10244 28422 10272 30126
rect 10232 28416 10284 28422
rect 10232 28358 10284 28364
rect 10048 28212 10100 28218
rect 10048 28154 10100 28160
rect 9956 28008 10008 28014
rect 9956 27950 10008 27956
rect 9824 27288 9904 27316
rect 9772 27270 9824 27276
rect 9588 27056 9640 27062
rect 9588 26998 9640 27004
rect 9784 26790 9812 27270
rect 9772 26784 9824 26790
rect 9824 26732 9904 26738
rect 9772 26726 9904 26732
rect 9784 26710 9904 26726
rect 9772 26580 9824 26586
rect 9772 26522 9824 26528
rect 9496 26512 9548 26518
rect 9496 26454 9548 26460
rect 9404 26240 9456 26246
rect 9404 26182 9456 26188
rect 9128 25696 9180 25702
rect 9128 25638 9180 25644
rect 9140 25226 9168 25638
rect 9416 25430 9444 26182
rect 9680 25968 9732 25974
rect 9680 25910 9732 25916
rect 9496 25900 9548 25906
rect 9496 25842 9548 25848
rect 9508 25498 9536 25842
rect 9496 25492 9548 25498
rect 9496 25434 9548 25440
rect 9404 25424 9456 25430
rect 9404 25366 9456 25372
rect 9128 25220 9180 25226
rect 9128 25162 9180 25168
rect 8864 24670 9076 24698
rect 8864 23118 8892 24670
rect 9036 23724 9088 23730
rect 9036 23666 9088 23672
rect 8852 23112 8904 23118
rect 8852 23054 8904 23060
rect 8760 23044 8812 23050
rect 8760 22986 8812 22992
rect 8772 22778 8800 22986
rect 8864 22778 8892 23054
rect 8944 22976 8996 22982
rect 8944 22918 8996 22924
rect 8760 22772 8812 22778
rect 8760 22714 8812 22720
rect 8852 22772 8904 22778
rect 8852 22714 8904 22720
rect 8956 22438 8984 22918
rect 9048 22778 9076 23666
rect 9036 22772 9088 22778
rect 9036 22714 9088 22720
rect 8944 22432 8996 22438
rect 8944 22374 8996 22380
rect 8956 22166 8984 22374
rect 8944 22160 8996 22166
rect 8944 22102 8996 22108
rect 9416 22094 9444 25366
rect 9692 24954 9720 25910
rect 9784 25838 9812 26522
rect 9772 25832 9824 25838
rect 9772 25774 9824 25780
rect 9876 25702 9904 26710
rect 9968 26586 9996 27950
rect 9956 26580 10008 26586
rect 9956 26522 10008 26528
rect 10060 25922 10088 28154
rect 10140 27396 10192 27402
rect 10140 27338 10192 27344
rect 10152 27130 10180 27338
rect 10140 27124 10192 27130
rect 10140 27066 10192 27072
rect 10336 26081 10364 30280
rect 10428 29102 10456 30382
rect 10704 30258 10732 31622
rect 10600 30252 10652 30258
rect 10600 30194 10652 30200
rect 10692 30252 10744 30258
rect 10692 30194 10744 30200
rect 10612 29850 10640 30194
rect 10600 29844 10652 29850
rect 10600 29786 10652 29792
rect 10508 29504 10560 29510
rect 10508 29446 10560 29452
rect 10416 29096 10468 29102
rect 10416 29038 10468 29044
rect 10428 26926 10456 29038
rect 10416 26920 10468 26926
rect 10520 26897 10548 29446
rect 10612 29306 10640 29786
rect 10600 29300 10652 29306
rect 10600 29242 10652 29248
rect 10692 27532 10744 27538
rect 10692 27474 10744 27480
rect 10598 27024 10654 27033
rect 10598 26959 10600 26968
rect 10652 26959 10654 26968
rect 10600 26930 10652 26936
rect 10416 26862 10468 26868
rect 10506 26888 10562 26897
rect 10506 26823 10562 26832
rect 10508 26784 10560 26790
rect 10508 26726 10560 26732
rect 10416 26240 10468 26246
rect 10416 26182 10468 26188
rect 10322 26072 10378 26081
rect 10244 26030 10322 26058
rect 10060 25906 10180 25922
rect 10060 25900 10192 25906
rect 10060 25894 10140 25900
rect 10140 25842 10192 25848
rect 9864 25696 9916 25702
rect 9864 25638 9916 25644
rect 9772 25288 9824 25294
rect 9772 25230 9824 25236
rect 9680 24948 9732 24954
rect 9680 24890 9732 24896
rect 9784 24614 9812 25230
rect 10140 25220 10192 25226
rect 10140 25162 10192 25168
rect 10152 24954 10180 25162
rect 10140 24948 10192 24954
rect 10140 24890 10192 24896
rect 10048 24676 10100 24682
rect 10048 24618 10100 24624
rect 9772 24608 9824 24614
rect 9772 24550 9824 24556
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 9692 22574 9720 24210
rect 9784 24206 9812 24550
rect 10060 24410 10088 24618
rect 10244 24614 10272 26030
rect 10322 26007 10378 26016
rect 10428 25906 10456 26182
rect 10520 25922 10548 26726
rect 10600 26308 10652 26314
rect 10600 26250 10652 26256
rect 10612 26042 10640 26250
rect 10600 26036 10652 26042
rect 10600 25978 10652 25984
rect 10324 25900 10376 25906
rect 10324 25842 10376 25848
rect 10416 25900 10468 25906
rect 10520 25894 10640 25922
rect 10416 25842 10468 25848
rect 10336 25158 10364 25842
rect 10324 25152 10376 25158
rect 10324 25094 10376 25100
rect 10336 24954 10364 25094
rect 10324 24948 10376 24954
rect 10324 24890 10376 24896
rect 10232 24608 10284 24614
rect 10232 24550 10284 24556
rect 10048 24404 10100 24410
rect 10048 24346 10100 24352
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 9784 23730 9812 24142
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 9784 23186 9812 23666
rect 9772 23180 9824 23186
rect 9772 23122 9824 23128
rect 9784 22642 9812 23122
rect 10060 23118 10088 24346
rect 10140 23860 10192 23866
rect 10244 23848 10272 24550
rect 10192 23820 10272 23848
rect 10140 23802 10192 23808
rect 10232 23520 10284 23526
rect 10232 23462 10284 23468
rect 10244 23118 10272 23462
rect 10428 23322 10456 25842
rect 10508 25696 10560 25702
rect 10508 25638 10560 25644
rect 10416 23316 10468 23322
rect 10416 23258 10468 23264
rect 10048 23112 10100 23118
rect 10048 23054 10100 23060
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 9956 22976 10008 22982
rect 9956 22918 10008 22924
rect 9968 22710 9996 22918
rect 10244 22778 10272 23054
rect 10232 22772 10284 22778
rect 10232 22714 10284 22720
rect 10520 22710 10548 25638
rect 10612 25401 10640 25894
rect 10598 25392 10654 25401
rect 10598 25327 10654 25336
rect 10704 23186 10732 27474
rect 10692 23180 10744 23186
rect 10692 23122 10744 23128
rect 9956 22704 10008 22710
rect 9956 22646 10008 22652
rect 10508 22704 10560 22710
rect 10508 22646 10560 22652
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 10416 22636 10468 22642
rect 10416 22578 10468 22584
rect 9680 22568 9732 22574
rect 9680 22510 9732 22516
rect 8680 22066 8892 22094
rect 9416 22066 9536 22094
rect 8300 21684 8352 21690
rect 8300 21626 8352 21632
rect 8116 21616 8168 21622
rect 8116 21558 8168 21564
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 8036 21146 8064 21422
rect 7840 21140 7892 21146
rect 7840 21082 7892 21088
rect 8024 21140 8076 21146
rect 8024 21082 8076 21088
rect 7472 20936 7524 20942
rect 7472 20878 7524 20884
rect 8036 20874 8064 21082
rect 7656 20868 7708 20874
rect 7656 20810 7708 20816
rect 8024 20868 8076 20874
rect 8024 20810 8076 20816
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7392 18290 7420 19246
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7196 17808 7248 17814
rect 7196 17750 7248 17756
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6748 16794 6776 17138
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6656 15706 6684 16050
rect 6736 15904 6788 15910
rect 6840 15858 6868 17070
rect 7024 16794 7052 17070
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 6788 15852 6868 15858
rect 6736 15846 6868 15852
rect 6748 15830 6868 15846
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 6840 15434 6868 15830
rect 6828 15428 6880 15434
rect 6828 15370 6880 15376
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6748 14074 6776 14214
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 12850 6868 13670
rect 6932 13530 6960 13942
rect 7024 13870 7052 15302
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7024 13530 7052 13806
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 6932 12986 6960 13466
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 7208 12782 7236 17750
rect 7392 17542 7420 18226
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7392 16658 7420 17478
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7576 15706 7604 16050
rect 7668 15706 7696 20810
rect 8128 20466 8156 21558
rect 8404 21321 8432 22066
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 8390 21312 8446 21321
rect 8390 21247 8446 21256
rect 8404 21146 8432 21247
rect 8392 21140 8444 21146
rect 8392 21082 8444 21088
rect 8404 20942 8432 21082
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 8116 20460 8168 20466
rect 8116 20402 8168 20408
rect 8496 19990 8524 21966
rect 8864 21486 8892 22066
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 9312 20800 9364 20806
rect 9312 20742 9364 20748
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 8956 20534 8984 20742
rect 9324 20602 9352 20742
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 8944 20528 8996 20534
rect 8944 20470 8996 20476
rect 8484 19984 8536 19990
rect 8404 19944 8484 19972
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 7944 18970 7972 19314
rect 8116 19168 8168 19174
rect 8116 19110 8168 19116
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 7932 18964 7984 18970
rect 7932 18906 7984 18912
rect 7932 18828 7984 18834
rect 7932 18770 7984 18776
rect 7944 18086 7972 18770
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7760 17338 7788 17614
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7944 15858 7972 18022
rect 8024 16516 8076 16522
rect 8024 16458 8076 16464
rect 8036 16250 8064 16458
rect 8024 16244 8076 16250
rect 8024 16186 8076 16192
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 7668 15502 7696 15642
rect 7760 15570 7788 15846
rect 7944 15830 8064 15858
rect 7748 15564 7800 15570
rect 7748 15506 7800 15512
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7668 14006 7696 15438
rect 7932 15360 7984 15366
rect 7932 15302 7984 15308
rect 7944 15026 7972 15302
rect 8036 15026 8064 15830
rect 8128 15706 8156 19110
rect 8312 18698 8340 19110
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 8116 15700 8168 15706
rect 8116 15642 8168 15648
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7760 14074 7788 14350
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7656 14000 7708 14006
rect 7656 13942 7708 13948
rect 7668 13870 7696 13942
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 8036 12434 8064 14962
rect 6564 12406 6684 12434
rect 6000 12164 6052 12170
rect 6000 12106 6052 12112
rect 6460 12164 6512 12170
rect 6460 12106 6512 12112
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5736 10606 5764 10746
rect 5906 10704 5962 10713
rect 5906 10639 5908 10648
rect 5960 10639 5962 10648
rect 5908 10610 5960 10616
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5644 9994 5672 10202
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5552 9722 5672 9738
rect 5552 9716 5684 9722
rect 5552 9710 5632 9716
rect 5632 9658 5684 9664
rect 5736 9654 5764 9998
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5540 9648 5592 9654
rect 5354 9616 5410 9625
rect 5540 9590 5592 9596
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 5354 9551 5410 9560
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5460 8906 5488 9318
rect 5552 9178 5580 9590
rect 5920 9518 5948 9862
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 6012 8566 6040 12106
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6104 11286 6132 11494
rect 6092 11280 6144 11286
rect 6092 11222 6144 11228
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6090 9616 6146 9625
rect 6380 9586 6408 9930
rect 6656 9586 6684 12406
rect 7944 12406 8064 12434
rect 7944 12306 7972 12406
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6748 11762 6776 12106
rect 7944 12102 7972 12242
rect 8128 12238 8156 15642
rect 8404 14074 8432 19944
rect 8484 19926 8536 19932
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 9128 19372 9180 19378
rect 9128 19314 9180 19320
rect 9048 19174 9076 19314
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8956 18358 8984 18566
rect 8944 18352 8996 18358
rect 8944 18294 8996 18300
rect 9048 17066 9076 19110
rect 9140 18698 9168 19314
rect 9416 18834 9444 20742
rect 9312 18828 9364 18834
rect 9312 18770 9364 18776
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 9128 18692 9180 18698
rect 9128 18634 9180 18640
rect 9140 18426 9168 18634
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9324 18086 9352 18770
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9312 17536 9364 17542
rect 9416 17524 9444 18634
rect 9364 17496 9444 17524
rect 9312 17478 9364 17484
rect 9324 17202 9352 17478
rect 9508 17338 9536 22066
rect 9692 21962 9720 22510
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9784 21622 9812 22578
rect 9864 22092 9916 22098
rect 9864 22034 9916 22040
rect 9876 21690 9904 22034
rect 10428 21894 10456 22578
rect 10416 21888 10468 21894
rect 10416 21830 10468 21836
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 9772 21616 9824 21622
rect 9772 21558 9824 21564
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9600 18834 9628 21286
rect 9784 21010 9812 21558
rect 9772 21004 9824 21010
rect 9772 20946 9824 20952
rect 9876 20942 9904 21626
rect 10416 21344 10468 21350
rect 10416 21286 10468 21292
rect 9864 20936 9916 20942
rect 9864 20878 9916 20884
rect 10324 20868 10376 20874
rect 10324 20810 10376 20816
rect 10336 20602 10364 20810
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10232 20256 10284 20262
rect 10232 20198 10284 20204
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 9600 18426 9628 18770
rect 9692 18630 9720 19994
rect 10244 19378 10272 20198
rect 10336 19768 10364 20402
rect 10428 20398 10456 21286
rect 10796 20482 10824 32506
rect 11060 32360 11112 32366
rect 11060 32302 11112 32308
rect 11072 32026 11100 32302
rect 11060 32020 11112 32026
rect 11060 31962 11112 31968
rect 10876 31340 10928 31346
rect 10876 31282 10928 31288
rect 11060 31340 11112 31346
rect 11164 31328 11192 33798
rect 11532 33454 11560 34478
rect 11610 34439 11612 34448
rect 11664 34439 11666 34448
rect 11612 34410 11664 34416
rect 11796 33516 11848 33522
rect 11796 33458 11848 33464
rect 11520 33448 11572 33454
rect 11520 33390 11572 33396
rect 11532 32366 11560 33390
rect 11808 33114 11836 33458
rect 11796 33108 11848 33114
rect 11796 33050 11848 33056
rect 11796 32904 11848 32910
rect 11796 32846 11848 32852
rect 11520 32360 11572 32366
rect 11520 32302 11572 32308
rect 11808 31414 11836 32846
rect 11900 32774 11928 35022
rect 12084 34610 12112 35566
rect 14004 35488 14056 35494
rect 14004 35430 14056 35436
rect 18880 35488 18932 35494
rect 18880 35430 18932 35436
rect 14016 35154 14044 35430
rect 17224 35284 17276 35290
rect 17224 35226 17276 35232
rect 14004 35148 14056 35154
rect 14004 35090 14056 35096
rect 13636 34944 13688 34950
rect 13636 34886 13688 34892
rect 13728 34944 13780 34950
rect 13728 34886 13780 34892
rect 12072 34604 12124 34610
rect 12072 34546 12124 34552
rect 13176 34604 13228 34610
rect 13176 34546 13228 34552
rect 12084 32774 12112 34546
rect 13188 34202 13216 34546
rect 13648 34406 13676 34886
rect 13740 34610 13768 34886
rect 13728 34604 13780 34610
rect 13728 34546 13780 34552
rect 13360 34400 13412 34406
rect 13360 34342 13412 34348
rect 13636 34400 13688 34406
rect 13636 34342 13688 34348
rect 13176 34196 13228 34202
rect 13176 34138 13228 34144
rect 13372 33998 13400 34342
rect 13452 34196 13504 34202
rect 13452 34138 13504 34144
rect 13360 33992 13412 33998
rect 13360 33934 13412 33940
rect 13464 33930 13492 34138
rect 13452 33924 13504 33930
rect 13452 33866 13504 33872
rect 13648 33862 13676 34342
rect 13728 34060 13780 34066
rect 13728 34002 13780 34008
rect 13740 33969 13768 34002
rect 13726 33960 13782 33969
rect 13726 33895 13782 33904
rect 13636 33856 13688 33862
rect 13636 33798 13688 33804
rect 12164 33312 12216 33318
rect 12164 33254 12216 33260
rect 12176 32910 12204 33254
rect 12164 32904 12216 32910
rect 12164 32846 12216 32852
rect 12992 32904 13044 32910
rect 12992 32846 13044 32852
rect 13176 32904 13228 32910
rect 13176 32846 13228 32852
rect 11888 32768 11940 32774
rect 12072 32768 12124 32774
rect 11888 32710 11940 32716
rect 12070 32736 12072 32745
rect 12124 32736 12126 32745
rect 11900 31754 11928 32710
rect 12070 32671 12126 32680
rect 12084 31822 12112 32671
rect 13004 32570 13032 32846
rect 12992 32564 13044 32570
rect 12992 32506 13044 32512
rect 12716 32496 12768 32502
rect 12900 32496 12952 32502
rect 12768 32444 12900 32450
rect 12716 32438 12952 32444
rect 12624 32428 12676 32434
rect 12728 32422 12940 32438
rect 12624 32370 12676 32376
rect 12636 32026 12664 32370
rect 12624 32020 12676 32026
rect 12624 31962 12676 31968
rect 12716 31884 12768 31890
rect 12716 31826 12768 31832
rect 12072 31816 12124 31822
rect 11992 31776 12072 31804
rect 11888 31748 11940 31754
rect 11888 31690 11940 31696
rect 11796 31408 11848 31414
rect 11796 31350 11848 31356
rect 11112 31300 11192 31328
rect 11244 31340 11296 31346
rect 11060 31282 11112 31288
rect 11244 31282 11296 31288
rect 10888 30870 10916 31282
rect 10876 30864 10928 30870
rect 10876 30806 10928 30812
rect 11060 30320 11112 30326
rect 11058 30288 11060 30297
rect 11112 30288 11114 30297
rect 11058 30223 11114 30232
rect 11256 30122 11284 31282
rect 11336 30728 11388 30734
rect 11336 30670 11388 30676
rect 11244 30116 11296 30122
rect 11244 30058 11296 30064
rect 11060 30048 11112 30054
rect 11060 29990 11112 29996
rect 11072 29850 11100 29990
rect 11060 29844 11112 29850
rect 11060 29786 11112 29792
rect 11348 29714 11376 30670
rect 11888 30252 11940 30258
rect 11888 30194 11940 30200
rect 11336 29708 11388 29714
rect 11336 29650 11388 29656
rect 11796 27872 11848 27878
rect 11796 27814 11848 27820
rect 11808 27470 11836 27814
rect 11900 27520 11928 30194
rect 11992 29170 12020 31776
rect 12072 31758 12124 31764
rect 12728 31754 12756 31826
rect 13004 31822 13032 32506
rect 13084 32224 13136 32230
rect 13084 32166 13136 32172
rect 12992 31816 13044 31822
rect 12992 31758 13044 31764
rect 12728 31726 12940 31754
rect 12072 31680 12124 31686
rect 12072 31622 12124 31628
rect 12084 31346 12112 31622
rect 12348 31476 12400 31482
rect 12348 31418 12400 31424
rect 12072 31340 12124 31346
rect 12072 31282 12124 31288
rect 12360 31142 12388 31418
rect 12716 31408 12768 31414
rect 12716 31350 12768 31356
rect 12532 31340 12584 31346
rect 12532 31282 12584 31288
rect 12544 31142 12572 31282
rect 12728 31142 12756 31350
rect 12348 31136 12400 31142
rect 12348 31078 12400 31084
rect 12532 31136 12584 31142
rect 12532 31078 12584 31084
rect 12716 31136 12768 31142
rect 12716 31078 12768 31084
rect 11980 29164 12032 29170
rect 11980 29106 12032 29112
rect 12164 28076 12216 28082
rect 12164 28018 12216 28024
rect 12176 27606 12204 28018
rect 12164 27600 12216 27606
rect 12164 27542 12216 27548
rect 11980 27532 12032 27538
rect 11900 27492 11980 27520
rect 11980 27474 12032 27480
rect 11796 27464 11848 27470
rect 11796 27406 11848 27412
rect 10968 27328 11020 27334
rect 10968 27270 11020 27276
rect 11612 27328 11664 27334
rect 11612 27270 11664 27276
rect 10980 27130 11008 27270
rect 10968 27124 11020 27130
rect 10968 27066 11020 27072
rect 11624 27062 11652 27270
rect 11808 27062 11836 27406
rect 11992 27062 12020 27474
rect 12360 27130 12388 31078
rect 12544 27878 12572 31078
rect 12728 30258 12756 31078
rect 12912 30734 12940 31726
rect 12900 30728 12952 30734
rect 12900 30670 12952 30676
rect 12808 30660 12860 30666
rect 12808 30602 12860 30608
rect 12820 30394 12848 30602
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 13096 30326 13124 32166
rect 13084 30320 13136 30326
rect 13084 30262 13136 30268
rect 12716 30252 12768 30258
rect 12716 30194 12768 30200
rect 13096 29646 13124 30262
rect 13188 30122 13216 32846
rect 13360 32768 13412 32774
rect 13360 32710 13412 32716
rect 13544 32768 13596 32774
rect 13544 32710 13596 32716
rect 13372 32366 13400 32710
rect 13360 32360 13412 32366
rect 13360 32302 13412 32308
rect 13268 30728 13320 30734
rect 13268 30670 13320 30676
rect 13280 30190 13308 30670
rect 13268 30184 13320 30190
rect 13268 30126 13320 30132
rect 13176 30116 13228 30122
rect 13176 30058 13228 30064
rect 13084 29640 13136 29646
rect 13084 29582 13136 29588
rect 12992 29096 13044 29102
rect 13280 29050 13308 30126
rect 12992 29038 13044 29044
rect 13004 28014 13032 29038
rect 13188 29022 13308 29050
rect 12992 28008 13044 28014
rect 12992 27950 13044 27956
rect 12532 27872 12584 27878
rect 12532 27814 12584 27820
rect 13084 27872 13136 27878
rect 13084 27814 13136 27820
rect 12900 27396 12952 27402
rect 12900 27338 12952 27344
rect 12624 27328 12676 27334
rect 12624 27270 12676 27276
rect 12636 27130 12664 27270
rect 12348 27124 12400 27130
rect 12348 27066 12400 27072
rect 12624 27124 12676 27130
rect 12624 27066 12676 27072
rect 11612 27056 11664 27062
rect 11612 26998 11664 27004
rect 11796 27056 11848 27062
rect 11796 26998 11848 27004
rect 11980 27056 12032 27062
rect 11980 26998 12032 27004
rect 12808 27056 12860 27062
rect 12808 26998 12860 27004
rect 12716 26988 12768 26994
rect 12716 26930 12768 26936
rect 11794 26888 11850 26897
rect 11794 26823 11850 26832
rect 11152 26784 11204 26790
rect 11152 26726 11204 26732
rect 11520 26784 11572 26790
rect 11520 26726 11572 26732
rect 10968 25832 11020 25838
rect 10966 25800 10968 25809
rect 11020 25800 11022 25809
rect 10966 25735 11022 25744
rect 10874 25392 10930 25401
rect 10874 25327 10930 25336
rect 10888 23322 10916 25327
rect 10968 25220 11020 25226
rect 10968 25162 11020 25168
rect 10980 24886 11008 25162
rect 11060 24948 11112 24954
rect 11060 24890 11112 24896
rect 10968 24880 11020 24886
rect 10968 24822 11020 24828
rect 11072 24750 11100 24890
rect 11060 24744 11112 24750
rect 11060 24686 11112 24692
rect 11072 24274 11100 24686
rect 11164 24342 11192 26726
rect 11336 26444 11388 26450
rect 11336 26386 11388 26392
rect 11348 25974 11376 26386
rect 11532 26382 11560 26726
rect 11704 26512 11756 26518
rect 11702 26480 11704 26489
rect 11756 26480 11758 26489
rect 11702 26415 11758 26424
rect 11520 26376 11572 26382
rect 11520 26318 11572 26324
rect 11336 25968 11388 25974
rect 11336 25910 11388 25916
rect 11704 25764 11756 25770
rect 11704 25706 11756 25712
rect 11716 25294 11744 25706
rect 11704 25288 11756 25294
rect 11704 25230 11756 25236
rect 11704 24608 11756 24614
rect 11704 24550 11756 24556
rect 11152 24336 11204 24342
rect 11152 24278 11204 24284
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 11336 23588 11388 23594
rect 11336 23530 11388 23536
rect 10876 23316 10928 23322
rect 10876 23258 10928 23264
rect 10888 23118 10916 23258
rect 10968 23180 11020 23186
rect 10968 23122 11020 23128
rect 10876 23112 10928 23118
rect 10876 23054 10928 23060
rect 10980 21690 11008 23122
rect 11348 23118 11376 23530
rect 11152 23112 11204 23118
rect 11336 23112 11388 23118
rect 11204 23060 11284 23066
rect 11152 23054 11284 23060
rect 11336 23054 11388 23060
rect 11164 23038 11284 23054
rect 11256 22438 11284 23038
rect 11244 22432 11296 22438
rect 11244 22374 11296 22380
rect 11256 22030 11284 22374
rect 11244 22024 11296 22030
rect 11244 21966 11296 21972
rect 10968 21684 11020 21690
rect 10968 21626 11020 21632
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 11164 20602 11192 20742
rect 11152 20596 11204 20602
rect 11152 20538 11204 20544
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 10704 20454 10824 20482
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10428 19922 10456 20334
rect 10416 19916 10468 19922
rect 10416 19858 10468 19864
rect 10416 19780 10468 19786
rect 10336 19740 10416 19768
rect 10416 19722 10468 19728
rect 10428 19689 10456 19722
rect 10414 19680 10470 19689
rect 10414 19615 10470 19624
rect 10704 19446 10732 20454
rect 11624 19718 11652 20538
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 10692 19440 10744 19446
rect 10692 19382 10744 19388
rect 10782 19408 10838 19417
rect 10232 19372 10284 19378
rect 10782 19343 10838 19352
rect 11244 19372 11296 19378
rect 10232 19314 10284 19320
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 10692 19304 10744 19310
rect 10692 19246 10744 19252
rect 9876 19174 9904 19246
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9876 18154 9904 19110
rect 10324 18692 10376 18698
rect 10324 18634 10376 18640
rect 10336 18426 10364 18634
rect 10704 18630 10732 19246
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10704 18426 10732 18566
rect 10796 18426 10824 19343
rect 11244 19314 11296 19320
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10416 18352 10468 18358
rect 10416 18294 10468 18300
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9600 17898 9628 18022
rect 9600 17870 9720 17898
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 8484 17060 8536 17066
rect 8484 17002 8536 17008
rect 9036 17060 9088 17066
rect 9036 17002 9088 17008
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6748 11150 6776 11698
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6748 9586 6776 11086
rect 7024 11082 7052 12038
rect 7392 11354 7420 12038
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7484 11218 7512 12038
rect 7944 11898 7972 12038
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7668 11354 7696 11698
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 8220 11218 8248 12718
rect 8496 12374 8524 17002
rect 9324 16658 9352 17138
rect 9692 16794 9720 17870
rect 10336 17746 10364 18226
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9876 17270 9904 17478
rect 9864 17264 9916 17270
rect 9864 17206 9916 17212
rect 10336 16998 10364 17682
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8956 16114 8984 16390
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 9048 15366 9076 15982
rect 9128 15564 9180 15570
rect 9128 15506 9180 15512
rect 9036 15360 9088 15366
rect 9034 15328 9036 15337
rect 9088 15328 9090 15337
rect 9034 15263 9090 15272
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8772 12238 8800 14010
rect 9140 13394 9168 15506
rect 9232 15434 9260 16050
rect 9324 15570 9352 16594
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9232 15162 9260 15370
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9324 15094 9352 15506
rect 9312 15088 9364 15094
rect 9312 15030 9364 15036
rect 9324 13938 9352 15030
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9324 13326 9352 13874
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 8852 13184 8904 13190
rect 9036 13184 9088 13190
rect 8904 13132 9036 13138
rect 8852 13126 9088 13132
rect 8864 13110 9076 13126
rect 8864 12850 8892 13110
rect 9416 12918 9444 16050
rect 9496 14340 9548 14346
rect 9496 14282 9548 14288
rect 9508 13734 9536 14282
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9508 13258 9536 13670
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9496 13252 9548 13258
rect 9496 13194 9548 13200
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 9416 12170 9444 12854
rect 9600 12434 9628 13330
rect 9692 12850 9720 16730
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9508 12406 9628 12434
rect 9784 12434 9812 15846
rect 9956 15428 10008 15434
rect 9956 15370 10008 15376
rect 9968 15162 9996 15370
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9876 14006 9904 14214
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 9784 12406 9904 12434
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8404 11558 8432 12038
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 6090 9551 6146 9560
rect 6368 9580 6420 9586
rect 6104 9518 6132 9551
rect 6368 9522 6420 9528
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6380 9178 6408 9522
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6656 9042 6684 9522
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6748 8838 6776 9522
rect 7392 9178 7420 9522
rect 7484 9382 7512 11154
rect 8404 11150 8432 11494
rect 9324 11354 9352 11698
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8680 10266 8708 10950
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 8772 10266 8800 10746
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8680 10062 8708 10202
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 7852 9722 7880 9998
rect 9416 9994 9444 12106
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 9404 9988 9456 9994
rect 9404 9930 9456 9936
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 6828 8968 6880 8974
rect 6826 8936 6828 8945
rect 6880 8936 6882 8945
rect 6826 8871 6882 8880
rect 7484 8838 7512 9318
rect 7852 8974 7880 9658
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 6932 7886 6960 8434
rect 7760 7954 7788 8774
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 8036 7886 8064 9930
rect 9508 9874 9536 12406
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9692 10962 9720 11154
rect 9784 11150 9812 11494
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9600 10934 9720 10962
rect 9600 9926 9628 10934
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9784 10033 9812 10066
rect 9770 10024 9826 10033
rect 9770 9959 9826 9968
rect 9416 9846 9536 9874
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8220 8498 8248 9454
rect 8956 9178 8984 9522
rect 9416 9450 9444 9846
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 9416 9110 9444 9386
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9600 8838 9628 9862
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9692 8838 9720 8978
rect 9784 8974 9812 9658
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 6932 7478 6960 7822
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 7300 7410 7328 7686
rect 8036 7546 8064 7822
rect 9600 7750 9628 8774
rect 9876 8634 9904 12406
rect 10060 11218 10088 12786
rect 10336 12374 10364 16934
rect 10428 14482 10456 18294
rect 10692 17604 10744 17610
rect 10692 17546 10744 17552
rect 10704 17338 10732 17546
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10888 16114 10916 17478
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10796 15162 10824 15302
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10888 15094 10916 16050
rect 10876 15088 10928 15094
rect 10876 15030 10928 15036
rect 11072 14482 11100 19110
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 11164 17338 11192 17546
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 11164 16250 11192 16458
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11164 16114 11192 16186
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11256 15026 11284 19314
rect 11624 17542 11652 19654
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 11612 17536 11664 17542
rect 11612 17478 11664 17484
rect 11336 15972 11388 15978
rect 11336 15914 11388 15920
rect 11348 15094 11376 15914
rect 11336 15088 11388 15094
rect 11336 15030 11388 15036
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11256 14822 11284 14962
rect 11440 14958 11468 17478
rect 11520 17128 11572 17134
rect 11520 17070 11572 17076
rect 11532 16658 11560 17070
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11428 14952 11480 14958
rect 11428 14894 11480 14900
rect 11532 14822 11560 15302
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 10416 14476 10468 14482
rect 10416 14418 10468 14424
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 10428 14006 10456 14418
rect 10692 14340 10744 14346
rect 10692 14282 10744 14288
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 10704 14074 10732 14282
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10416 14000 10468 14006
rect 10416 13942 10468 13948
rect 10140 12368 10192 12374
rect 10140 12310 10192 12316
rect 10324 12368 10376 12374
rect 10324 12310 10376 12316
rect 10152 11218 10180 12310
rect 10336 11558 10364 12310
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10060 10810 10088 11154
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10060 10606 10088 10746
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9968 8956 9996 10134
rect 10060 10062 10088 10406
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 10060 9178 10088 9862
rect 10152 9382 10180 9930
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10152 8974 10180 9318
rect 10244 9042 10272 11086
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 10048 8968 10100 8974
rect 9968 8928 10048 8956
rect 10048 8910 10100 8916
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10336 8838 10364 11494
rect 10428 11354 10456 13942
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10704 11150 10732 12038
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10428 10810 10456 11086
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10796 10470 10824 14214
rect 11164 14074 11192 14282
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11152 12912 11204 12918
rect 11256 12900 11284 14758
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11532 13326 11560 13670
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11204 12872 11284 12900
rect 11152 12854 11204 12860
rect 11164 11830 11192 12854
rect 11624 12434 11652 17478
rect 11716 15994 11744 24550
rect 11808 23322 11836 26823
rect 12348 26784 12400 26790
rect 12348 26726 12400 26732
rect 12360 26586 12388 26726
rect 12728 26586 12756 26930
rect 12348 26580 12400 26586
rect 12348 26522 12400 26528
rect 12716 26580 12768 26586
rect 12716 26522 12768 26528
rect 12532 26308 12584 26314
rect 12532 26250 12584 26256
rect 12544 26042 12572 26250
rect 12728 26042 12756 26522
rect 12532 26036 12584 26042
rect 12532 25978 12584 25984
rect 12716 26036 12768 26042
rect 12716 25978 12768 25984
rect 12714 25528 12770 25537
rect 12714 25463 12716 25472
rect 12768 25463 12770 25472
rect 12716 25434 12768 25440
rect 12164 25220 12216 25226
rect 12164 25162 12216 25168
rect 12176 24410 12204 25162
rect 12532 24812 12584 24818
rect 12532 24754 12584 24760
rect 12164 24404 12216 24410
rect 12164 24346 12216 24352
rect 12256 24336 12308 24342
rect 12256 24278 12308 24284
rect 11796 23316 11848 23322
rect 11796 23258 11848 23264
rect 12164 23112 12216 23118
rect 12164 23054 12216 23060
rect 12070 22400 12126 22409
rect 12070 22335 12126 22344
rect 12084 22234 12112 22335
rect 12072 22228 12124 22234
rect 12072 22170 12124 22176
rect 12176 22030 12204 23054
rect 12268 22438 12296 24278
rect 12544 24206 12572 24754
rect 12716 24268 12768 24274
rect 12716 24210 12768 24216
rect 12532 24200 12584 24206
rect 12532 24142 12584 24148
rect 12440 24064 12492 24070
rect 12440 24006 12492 24012
rect 12452 23730 12480 24006
rect 12728 23866 12756 24210
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12440 23724 12492 23730
rect 12440 23666 12492 23672
rect 12728 23662 12756 23802
rect 12716 23656 12768 23662
rect 12716 23598 12768 23604
rect 12820 23322 12848 26998
rect 12912 25974 12940 27338
rect 13096 26994 13124 27814
rect 12992 26988 13044 26994
rect 12992 26930 13044 26936
rect 13084 26988 13136 26994
rect 13084 26930 13136 26936
rect 12900 25968 12952 25974
rect 12900 25910 12952 25916
rect 12912 24818 12940 25910
rect 13004 25498 13032 26930
rect 13096 26246 13124 26930
rect 13084 26240 13136 26246
rect 13084 26182 13136 26188
rect 12992 25492 13044 25498
rect 12992 25434 13044 25440
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 12900 24268 12952 24274
rect 12900 24210 12952 24216
rect 12808 23316 12860 23322
rect 12808 23258 12860 23264
rect 12716 23044 12768 23050
rect 12716 22986 12768 22992
rect 12728 22778 12756 22986
rect 12716 22772 12768 22778
rect 12716 22714 12768 22720
rect 12256 22432 12308 22438
rect 12256 22374 12308 22380
rect 12912 22234 12940 24210
rect 13004 24206 13032 25434
rect 13188 24342 13216 29022
rect 13372 28994 13400 32302
rect 13556 31346 13584 32710
rect 13648 32230 13676 33798
rect 13912 32972 13964 32978
rect 13912 32914 13964 32920
rect 13924 32570 13952 32914
rect 13912 32564 13964 32570
rect 13912 32506 13964 32512
rect 13636 32224 13688 32230
rect 13636 32166 13688 32172
rect 13544 31340 13596 31346
rect 13544 31282 13596 31288
rect 13636 30592 13688 30598
rect 13636 30534 13688 30540
rect 13648 30326 13676 30534
rect 13636 30320 13688 30326
rect 13636 30262 13688 30268
rect 13450 29064 13506 29073
rect 13450 28999 13506 29008
rect 13280 28966 13400 28994
rect 13280 26042 13308 28966
rect 13464 27062 13492 28999
rect 13544 27600 13596 27606
rect 13544 27542 13596 27548
rect 13452 27056 13504 27062
rect 13452 26998 13504 27004
rect 13360 26920 13412 26926
rect 13360 26862 13412 26868
rect 13372 26382 13400 26862
rect 13360 26376 13412 26382
rect 13360 26318 13412 26324
rect 13268 26036 13320 26042
rect 13268 25978 13320 25984
rect 13280 25838 13308 25978
rect 13268 25832 13320 25838
rect 13320 25792 13400 25820
rect 13268 25774 13320 25780
rect 13268 24880 13320 24886
rect 13268 24822 13320 24828
rect 13176 24336 13228 24342
rect 13176 24278 13228 24284
rect 12992 24200 13044 24206
rect 12992 24142 13044 24148
rect 13280 23866 13308 24822
rect 13372 24721 13400 25792
rect 13358 24712 13414 24721
rect 13358 24647 13414 24656
rect 13268 23860 13320 23866
rect 13268 23802 13320 23808
rect 13176 23724 13228 23730
rect 13176 23666 13228 23672
rect 13188 22574 13216 23666
rect 13280 22574 13308 23802
rect 13176 22568 13228 22574
rect 13176 22510 13228 22516
rect 13268 22568 13320 22574
rect 13268 22510 13320 22516
rect 12900 22228 12952 22234
rect 12900 22170 12952 22176
rect 12164 22024 12216 22030
rect 12164 21966 12216 21972
rect 12176 20942 12204 21966
rect 13188 21962 13216 22510
rect 13280 22234 13308 22510
rect 13268 22228 13320 22234
rect 13268 22170 13320 22176
rect 12808 21956 12860 21962
rect 12808 21898 12860 21904
rect 13176 21956 13228 21962
rect 13176 21898 13228 21904
rect 12820 21690 12848 21898
rect 13188 21690 13216 21898
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 13176 21684 13228 21690
rect 13176 21626 13228 21632
rect 13372 21486 13400 24647
rect 13556 24274 13584 27542
rect 14016 27520 14044 35090
rect 15108 35080 15160 35086
rect 15108 35022 15160 35028
rect 14464 34944 14516 34950
rect 14464 34886 14516 34892
rect 14476 34746 14504 34886
rect 14464 34740 14516 34746
rect 14464 34682 14516 34688
rect 14096 34672 14148 34678
rect 14096 34614 14148 34620
rect 14108 33114 14136 34614
rect 14476 33998 14504 34682
rect 15120 34678 15148 35022
rect 15568 35012 15620 35018
rect 15568 34954 15620 34960
rect 15580 34746 15608 34954
rect 16028 34944 16080 34950
rect 16028 34886 16080 34892
rect 16040 34746 16068 34886
rect 15568 34740 15620 34746
rect 15568 34682 15620 34688
rect 16028 34740 16080 34746
rect 16028 34682 16080 34688
rect 15108 34672 15160 34678
rect 15108 34614 15160 34620
rect 14740 34196 14792 34202
rect 14740 34138 14792 34144
rect 14752 33998 14780 34138
rect 14464 33992 14516 33998
rect 14464 33934 14516 33940
rect 14740 33992 14792 33998
rect 14740 33934 14792 33940
rect 15292 33992 15344 33998
rect 15292 33934 15344 33940
rect 14556 33924 14608 33930
rect 14556 33866 14608 33872
rect 14568 33658 14596 33866
rect 14924 33856 14976 33862
rect 14924 33798 14976 33804
rect 14556 33652 14608 33658
rect 14556 33594 14608 33600
rect 14936 33522 14964 33798
rect 14924 33516 14976 33522
rect 14924 33458 14976 33464
rect 15108 33516 15160 33522
rect 15108 33458 15160 33464
rect 14096 33108 14148 33114
rect 14096 33050 14148 33056
rect 14108 32978 14136 33050
rect 14096 32972 14148 32978
rect 14096 32914 14148 32920
rect 14188 32904 14240 32910
rect 14188 32846 14240 32852
rect 14200 32502 14228 32846
rect 14464 32836 14516 32842
rect 14464 32778 14516 32784
rect 14476 32570 14504 32778
rect 15120 32774 15148 33458
rect 14832 32768 14884 32774
rect 14832 32710 14884 32716
rect 15108 32768 15160 32774
rect 15108 32710 15160 32716
rect 14844 32570 14872 32710
rect 14372 32564 14424 32570
rect 14372 32506 14424 32512
rect 14464 32564 14516 32570
rect 14464 32506 14516 32512
rect 14832 32564 14884 32570
rect 14832 32506 14884 32512
rect 14188 32496 14240 32502
rect 14188 32438 14240 32444
rect 14096 30252 14148 30258
rect 14096 30194 14148 30200
rect 14108 29646 14136 30194
rect 14096 29640 14148 29646
rect 14096 29582 14148 29588
rect 14200 28218 14228 32438
rect 14384 32314 14412 32506
rect 15108 32496 15160 32502
rect 15108 32438 15160 32444
rect 15120 32366 15148 32438
rect 15108 32360 15160 32366
rect 14384 32286 14504 32314
rect 15108 32302 15160 32308
rect 14476 32230 14504 32286
rect 14556 32292 14608 32298
rect 14556 32234 14608 32240
rect 14464 32224 14516 32230
rect 14464 32166 14516 32172
rect 14568 31754 14596 32234
rect 14476 31726 14596 31754
rect 14476 30394 14504 31726
rect 15304 30734 15332 33934
rect 15660 33924 15712 33930
rect 15660 33866 15712 33872
rect 15384 33856 15436 33862
rect 15384 33798 15436 33804
rect 15396 33454 15424 33798
rect 15672 33522 15700 33866
rect 16040 33590 16068 34682
rect 17236 34678 17264 35226
rect 17408 35080 17460 35086
rect 17408 35022 17460 35028
rect 17224 34672 17276 34678
rect 17224 34614 17276 34620
rect 16212 34536 16264 34542
rect 16212 34478 16264 34484
rect 16120 34400 16172 34406
rect 16120 34342 16172 34348
rect 16132 33590 16160 34342
rect 16028 33584 16080 33590
rect 16028 33526 16080 33532
rect 16120 33584 16172 33590
rect 16120 33526 16172 33532
rect 15660 33516 15712 33522
rect 15660 33458 15712 33464
rect 15384 33448 15436 33454
rect 15384 33390 15436 33396
rect 15108 30728 15160 30734
rect 15108 30670 15160 30676
rect 15292 30728 15344 30734
rect 15292 30670 15344 30676
rect 14556 30660 14608 30666
rect 14556 30602 14608 30608
rect 14568 30394 14596 30602
rect 14464 30388 14516 30394
rect 14464 30330 14516 30336
rect 14556 30388 14608 30394
rect 14556 30330 14608 30336
rect 14280 30320 14332 30326
rect 14278 30288 14280 30297
rect 14332 30288 14334 30297
rect 14334 30246 14412 30274
rect 14278 30223 14334 30232
rect 14280 30048 14332 30054
rect 14280 29990 14332 29996
rect 14292 29714 14320 29990
rect 14384 29850 14412 30246
rect 14372 29844 14424 29850
rect 14372 29786 14424 29792
rect 14280 29708 14332 29714
rect 14280 29650 14332 29656
rect 14188 28212 14240 28218
rect 14188 28154 14240 28160
rect 14096 27532 14148 27538
rect 14016 27492 14096 27520
rect 14096 27474 14148 27480
rect 14108 27334 14136 27474
rect 13912 27328 13964 27334
rect 13912 27270 13964 27276
rect 14096 27328 14148 27334
rect 14096 27270 14148 27276
rect 13924 27062 13952 27270
rect 13912 27056 13964 27062
rect 13912 26998 13964 27004
rect 13728 26376 13780 26382
rect 13728 26318 13780 26324
rect 13636 26240 13688 26246
rect 13636 26182 13688 26188
rect 13648 25401 13676 26182
rect 13740 25906 13768 26318
rect 14108 26246 14136 27270
rect 14096 26240 14148 26246
rect 14096 26182 14148 26188
rect 13728 25900 13780 25906
rect 13728 25842 13780 25848
rect 13634 25392 13690 25401
rect 13634 25327 13690 25336
rect 13740 24818 13768 25842
rect 14004 25288 14056 25294
rect 14004 25230 14056 25236
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13728 24812 13780 24818
rect 13728 24754 13780 24760
rect 13544 24268 13596 24274
rect 13544 24210 13596 24216
rect 13452 24132 13504 24138
rect 13452 24074 13504 24080
rect 13464 22574 13492 24074
rect 13648 24070 13676 24754
rect 13636 24064 13688 24070
rect 13636 24006 13688 24012
rect 13544 22976 13596 22982
rect 13544 22918 13596 22924
rect 13556 22642 13584 22918
rect 13544 22636 13596 22642
rect 13544 22578 13596 22584
rect 13452 22568 13504 22574
rect 13452 22510 13504 22516
rect 13360 21480 13412 21486
rect 13360 21422 13412 21428
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 12348 20936 12400 20942
rect 12348 20878 12400 20884
rect 12360 20534 12388 20878
rect 12440 20868 12492 20874
rect 12440 20810 12492 20816
rect 12348 20528 12400 20534
rect 12348 20470 12400 20476
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 12084 18766 12112 19110
rect 12360 18766 12388 20334
rect 12452 20330 12480 20810
rect 13452 20800 13504 20806
rect 13452 20742 13504 20748
rect 13464 20466 13492 20742
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 12900 20392 12952 20398
rect 12900 20334 12952 20340
rect 12992 20392 13044 20398
rect 12992 20334 13044 20340
rect 12440 20324 12492 20330
rect 12440 20266 12492 20272
rect 12912 19990 12940 20334
rect 12532 19984 12584 19990
rect 12532 19926 12584 19932
rect 12900 19984 12952 19990
rect 12900 19926 12952 19932
rect 12438 19408 12494 19417
rect 12544 19360 12572 19926
rect 12808 19780 12860 19786
rect 12808 19722 12860 19728
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12494 19352 12572 19360
rect 12438 19343 12440 19352
rect 12492 19332 12572 19352
rect 12440 19314 12492 19320
rect 12728 19310 12756 19654
rect 12820 19514 12848 19722
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 13004 19334 13032 20334
rect 13464 19378 13492 20402
rect 13452 19372 13504 19378
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12728 18426 12756 19246
rect 12912 18970 12940 19314
rect 13004 19306 13216 19334
rect 13452 19314 13504 19320
rect 13648 19310 13676 24006
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 13832 21894 13860 22578
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13832 21622 13860 21830
rect 13820 21616 13872 21622
rect 13820 21558 13872 21564
rect 13912 19916 13964 19922
rect 13912 19858 13964 19864
rect 13924 19446 13952 19858
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13912 19440 13964 19446
rect 13912 19382 13964 19388
rect 12992 19236 13044 19242
rect 12992 19178 13044 19184
rect 12900 18964 12952 18970
rect 12900 18906 12952 18912
rect 13004 18698 13032 19178
rect 12992 18692 13044 18698
rect 12992 18634 13044 18640
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11808 16250 11836 17138
rect 11900 16658 11928 17750
rect 12084 17202 12112 18158
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12072 17196 12124 17202
rect 12072 17138 12124 17144
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 12268 16250 12296 17274
rect 12452 16794 12480 17478
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12728 16250 12756 18362
rect 13004 17542 13032 18634
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12728 16046 12756 16186
rect 12716 16040 12768 16046
rect 11716 15966 11836 15994
rect 12716 15982 12768 15988
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11716 15502 11744 15846
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11808 13433 11836 15966
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 11992 14618 12204 14634
rect 11992 14612 12216 14618
rect 11992 14606 12164 14612
rect 11992 14550 12020 14606
rect 12164 14554 12216 14560
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 12268 14482 12296 15438
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12452 14940 12480 15302
rect 12636 15162 12664 15370
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12624 14952 12676 14958
rect 12452 14912 12624 14940
rect 12624 14894 12676 14900
rect 12728 14482 12756 15982
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 12912 15366 12940 15642
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12820 14958 12848 15098
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 12268 14362 12296 14418
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11900 13530 11928 14010
rect 11992 13938 12020 14350
rect 12268 14334 12388 14362
rect 12360 14278 12388 14334
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11794 13424 11850 13433
rect 11794 13359 11850 13368
rect 11532 12406 11652 12434
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11348 11898 11376 12174
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10980 11354 11008 11698
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 10428 10062 10456 10202
rect 10888 10130 10916 11290
rect 11164 11150 11192 11766
rect 11256 11218 11284 11834
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11348 11150 11376 11834
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11164 10810 11192 11086
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11532 10266 11560 12406
rect 11808 10266 11836 13359
rect 11992 13258 12020 13874
rect 12268 13530 12296 14214
rect 12440 13932 12492 13938
rect 12624 13932 12676 13938
rect 12492 13892 12572 13920
rect 12440 13874 12492 13880
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 11980 13252 12032 13258
rect 11980 13194 12032 13200
rect 12268 12986 12296 13262
rect 12440 13252 12492 13258
rect 12440 13194 12492 13200
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12360 11354 12388 11698
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 11978 11112 12034 11121
rect 12452 11082 12480 13194
rect 12544 12782 12572 13892
rect 12624 13874 12676 13880
rect 12636 13530 12664 13874
rect 12728 13734 12756 14418
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12636 13025 12664 13126
rect 12622 13016 12678 13025
rect 12622 12951 12678 12960
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12544 11830 12572 12718
rect 12728 12646 12756 13398
rect 12912 13190 12940 15302
rect 13004 14260 13032 17478
rect 13096 17270 13124 18158
rect 13084 17264 13136 17270
rect 13084 17206 13136 17212
rect 13096 17066 13124 17206
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 13096 16114 13124 17002
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 13096 15570 13124 16050
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 13188 15337 13216 19306
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13372 18358 13400 19110
rect 13360 18352 13412 18358
rect 13360 18294 13412 18300
rect 13648 16726 13676 19246
rect 13740 18630 13768 19382
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13636 16720 13688 16726
rect 13636 16662 13688 16668
rect 13648 16590 13676 16662
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13740 16114 13768 18566
rect 14016 18358 14044 25230
rect 14096 24608 14148 24614
rect 14200 24562 14228 28154
rect 14280 27464 14332 27470
rect 14280 27406 14332 27412
rect 14292 27334 14320 27406
rect 14280 27328 14332 27334
rect 14280 27270 14332 27276
rect 14278 26616 14334 26625
rect 14278 26551 14334 26560
rect 14148 24556 14228 24562
rect 14096 24550 14228 24556
rect 14108 24534 14228 24550
rect 14108 23322 14136 24534
rect 14200 24410 14228 24534
rect 14188 24404 14240 24410
rect 14188 24346 14240 24352
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 14108 21146 14136 23258
rect 14292 22094 14320 26551
rect 14476 26466 14504 30330
rect 14556 30048 14608 30054
rect 14556 29990 14608 29996
rect 14568 29073 14596 29990
rect 15120 29646 15148 30670
rect 15292 30388 15344 30394
rect 15292 30330 15344 30336
rect 15200 30252 15252 30258
rect 15200 30194 15252 30200
rect 15212 29850 15240 30194
rect 15200 29844 15252 29850
rect 15200 29786 15252 29792
rect 14648 29640 14700 29646
rect 14648 29582 14700 29588
rect 15108 29640 15160 29646
rect 15108 29582 15160 29588
rect 14660 29170 14688 29582
rect 14648 29164 14700 29170
rect 14648 29106 14700 29112
rect 14554 29064 14610 29073
rect 14554 28999 14610 29008
rect 15016 28552 15068 28558
rect 15016 28494 15068 28500
rect 14556 28008 14608 28014
rect 14556 27950 14608 27956
rect 14568 27470 14596 27950
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14922 27432 14978 27441
rect 14568 26994 14596 27406
rect 14922 27367 14978 27376
rect 14556 26988 14608 26994
rect 14556 26930 14608 26936
rect 14832 26988 14884 26994
rect 14832 26930 14884 26936
rect 14740 26852 14792 26858
rect 14740 26794 14792 26800
rect 14384 26438 14504 26466
rect 14384 24614 14412 26438
rect 14464 26308 14516 26314
rect 14464 26250 14516 26256
rect 14372 24608 14424 24614
rect 14372 24550 14424 24556
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14384 22778 14412 23054
rect 14372 22772 14424 22778
rect 14372 22714 14424 22720
rect 14476 22094 14504 26250
rect 14648 25900 14700 25906
rect 14648 25842 14700 25848
rect 14660 25498 14688 25842
rect 14648 25492 14700 25498
rect 14648 25434 14700 25440
rect 14200 22066 14320 22094
rect 14384 22066 14504 22094
rect 14096 21140 14148 21146
rect 14096 21082 14148 21088
rect 14108 20942 14136 21082
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 14108 19718 14136 20402
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14004 18352 14056 18358
rect 14004 18294 14056 18300
rect 14096 18148 14148 18154
rect 14096 18090 14148 18096
rect 14004 18080 14056 18086
rect 14004 18022 14056 18028
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13832 16658 13860 17070
rect 14016 16794 14044 18022
rect 14108 17134 14136 18090
rect 14200 17270 14228 22066
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 14292 18970 14320 19450
rect 14384 19310 14412 22066
rect 14556 21344 14608 21350
rect 14556 21286 14608 21292
rect 14568 20874 14596 21286
rect 14556 20868 14608 20874
rect 14556 20810 14608 20816
rect 14568 20534 14596 20810
rect 14556 20528 14608 20534
rect 14556 20470 14608 20476
rect 14568 19854 14596 20470
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14660 19718 14688 20198
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14752 19446 14780 26794
rect 14844 25974 14872 26930
rect 14936 26625 14964 27367
rect 15028 27334 15056 28494
rect 15120 28014 15148 29582
rect 15304 29306 15332 30330
rect 15292 29300 15344 29306
rect 15292 29242 15344 29248
rect 15108 28008 15160 28014
rect 15108 27950 15160 27956
rect 15108 27396 15160 27402
rect 15108 27338 15160 27344
rect 15016 27328 15068 27334
rect 15016 27270 15068 27276
rect 14922 26616 14978 26625
rect 14922 26551 14978 26560
rect 15028 26314 15056 27270
rect 15120 26586 15148 27338
rect 15396 26586 15424 33390
rect 15568 32224 15620 32230
rect 15568 32166 15620 32172
rect 15580 31754 15608 32166
rect 15568 31748 15620 31754
rect 15568 31690 15620 31696
rect 15672 31482 15700 33458
rect 15844 33380 15896 33386
rect 15844 33322 15896 33328
rect 15856 31754 15884 33322
rect 16224 32570 16252 34478
rect 16500 34156 17080 34184
rect 16304 34128 16356 34134
rect 16304 34070 16356 34076
rect 16316 33930 16344 34070
rect 16500 33998 16528 34156
rect 16488 33992 16540 33998
rect 16488 33934 16540 33940
rect 16672 33992 16724 33998
rect 16672 33934 16724 33940
rect 16304 33924 16356 33930
rect 16304 33866 16356 33872
rect 16580 33856 16632 33862
rect 16580 33798 16632 33804
rect 16304 33652 16356 33658
rect 16304 33594 16356 33600
rect 16212 32564 16264 32570
rect 16212 32506 16264 32512
rect 16120 32292 16172 32298
rect 16120 32234 16172 32240
rect 15856 31726 16068 31754
rect 15660 31476 15712 31482
rect 15660 31418 15712 31424
rect 15660 30864 15712 30870
rect 15660 30806 15712 30812
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 15488 28150 15516 30670
rect 15568 30592 15620 30598
rect 15568 30534 15620 30540
rect 15580 30258 15608 30534
rect 15568 30252 15620 30258
rect 15568 30194 15620 30200
rect 15672 30190 15700 30806
rect 15752 30592 15804 30598
rect 15752 30534 15804 30540
rect 15764 30394 15792 30534
rect 15752 30388 15804 30394
rect 15752 30330 15804 30336
rect 15844 30252 15896 30258
rect 15844 30194 15896 30200
rect 15660 30184 15712 30190
rect 15660 30126 15712 30132
rect 15476 28144 15528 28150
rect 15476 28086 15528 28092
rect 15672 27606 15700 30126
rect 15752 29572 15804 29578
rect 15752 29514 15804 29520
rect 15764 29306 15792 29514
rect 15856 29510 15884 30194
rect 15844 29504 15896 29510
rect 15844 29446 15896 29452
rect 15856 29306 15884 29446
rect 15752 29300 15804 29306
rect 15752 29242 15804 29248
rect 15844 29300 15896 29306
rect 15844 29242 15896 29248
rect 16040 29102 16068 31726
rect 16132 31686 16160 32234
rect 16120 31680 16172 31686
rect 16120 31622 16172 31628
rect 16132 30870 16160 31622
rect 16120 30864 16172 30870
rect 16120 30806 16172 30812
rect 16316 30394 16344 33594
rect 16592 33386 16620 33798
rect 16684 33454 16712 33934
rect 17052 33590 17080 34156
rect 17224 34060 17276 34066
rect 17224 34002 17276 34008
rect 17040 33584 17092 33590
rect 17040 33526 17092 33532
rect 16672 33448 16724 33454
rect 16672 33390 16724 33396
rect 16580 33380 16632 33386
rect 16580 33322 16632 33328
rect 16684 32910 16712 33390
rect 16672 32904 16724 32910
rect 16672 32846 16724 32852
rect 16580 32564 16632 32570
rect 16580 32506 16632 32512
rect 16592 32366 16620 32506
rect 16580 32360 16632 32366
rect 16580 32302 16632 32308
rect 16488 31476 16540 31482
rect 16488 31418 16540 31424
rect 16304 30388 16356 30394
rect 16304 30330 16356 30336
rect 16212 30252 16264 30258
rect 16212 30194 16264 30200
rect 16224 30138 16252 30194
rect 16224 30110 16344 30138
rect 16316 30054 16344 30110
rect 16304 30048 16356 30054
rect 16304 29990 16356 29996
rect 16028 29096 16080 29102
rect 16028 29038 16080 29044
rect 16040 28994 16068 29038
rect 16040 28966 16160 28994
rect 15844 27668 15896 27674
rect 15844 27610 15896 27616
rect 15660 27600 15712 27606
rect 15712 27560 15792 27588
rect 15660 27542 15712 27548
rect 15108 26580 15160 26586
rect 15108 26522 15160 26528
rect 15384 26580 15436 26586
rect 15384 26522 15436 26528
rect 15016 26308 15068 26314
rect 15016 26250 15068 26256
rect 14832 25968 14884 25974
rect 14832 25910 14884 25916
rect 14924 25152 14976 25158
rect 15028 25140 15056 26250
rect 15108 26240 15160 26246
rect 15108 26182 15160 26188
rect 15120 25838 15148 26182
rect 15396 26042 15424 26522
rect 15384 26036 15436 26042
rect 15384 25978 15436 25984
rect 15660 26036 15712 26042
rect 15660 25978 15712 25984
rect 15108 25832 15160 25838
rect 15108 25774 15160 25780
rect 15568 25696 15620 25702
rect 15568 25638 15620 25644
rect 15200 25356 15252 25362
rect 15200 25298 15252 25304
rect 15108 25288 15160 25294
rect 15108 25230 15160 25236
rect 14976 25112 15056 25140
rect 14924 25094 14976 25100
rect 14924 24948 14976 24954
rect 14924 24890 14976 24896
rect 14936 24732 14964 24890
rect 15028 24886 15056 25112
rect 15120 24954 15148 25230
rect 15108 24948 15160 24954
rect 15108 24890 15160 24896
rect 15016 24880 15068 24886
rect 15016 24822 15068 24828
rect 15212 24732 15240 25298
rect 15580 25294 15608 25638
rect 15568 25288 15620 25294
rect 15568 25230 15620 25236
rect 15672 25226 15700 25978
rect 15660 25220 15712 25226
rect 15660 25162 15712 25168
rect 14936 24704 15240 24732
rect 15476 24608 15528 24614
rect 15672 24562 15700 25162
rect 15476 24550 15528 24556
rect 14832 23044 14884 23050
rect 14832 22986 14884 22992
rect 14844 22778 14872 22986
rect 14832 22772 14884 22778
rect 14832 22714 14884 22720
rect 15488 22166 15516 24550
rect 15580 24534 15700 24562
rect 15476 22160 15528 22166
rect 15476 22102 15528 22108
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 14844 21622 14872 21830
rect 15212 21690 15240 21830
rect 15200 21684 15252 21690
rect 15200 21626 15252 21632
rect 14832 21616 14884 21622
rect 14832 21558 14884 21564
rect 15580 20602 15608 24534
rect 15764 23798 15792 27560
rect 15856 26314 15884 27610
rect 16028 27464 16080 27470
rect 16028 27406 16080 27412
rect 15936 27328 15988 27334
rect 15936 27270 15988 27276
rect 15948 26382 15976 27270
rect 16040 27130 16068 27406
rect 16028 27124 16080 27130
rect 16028 27066 16080 27072
rect 15936 26376 15988 26382
rect 15936 26318 15988 26324
rect 16028 26376 16080 26382
rect 16028 26318 16080 26324
rect 15844 26308 15896 26314
rect 15844 26250 15896 26256
rect 16040 25498 16068 26318
rect 16132 25702 16160 28966
rect 16212 28212 16264 28218
rect 16212 28154 16264 28160
rect 16224 27470 16252 28154
rect 16212 27464 16264 27470
rect 16212 27406 16264 27412
rect 16224 27062 16252 27406
rect 16212 27056 16264 27062
rect 16212 26998 16264 27004
rect 16316 25809 16344 29990
rect 16396 27464 16448 27470
rect 16396 27406 16448 27412
rect 16408 26858 16436 27406
rect 16396 26852 16448 26858
rect 16396 26794 16448 26800
rect 16500 26586 16528 31418
rect 16592 30190 16620 32302
rect 16684 31822 16712 32846
rect 16764 32836 16816 32842
rect 16764 32778 16816 32784
rect 16672 31816 16724 31822
rect 16672 31758 16724 31764
rect 16580 30184 16632 30190
rect 16580 30126 16632 30132
rect 16684 29714 16712 31758
rect 16776 31414 16804 32778
rect 17038 32736 17094 32745
rect 17038 32671 17094 32680
rect 17052 32434 17080 32671
rect 17040 32428 17092 32434
rect 17040 32370 17092 32376
rect 17132 32360 17184 32366
rect 17132 32302 17184 32308
rect 17144 32026 17172 32302
rect 17132 32020 17184 32026
rect 17132 31962 17184 31968
rect 16764 31408 16816 31414
rect 16764 31350 16816 31356
rect 17144 31346 17172 31962
rect 16856 31340 16908 31346
rect 16856 31282 16908 31288
rect 17132 31340 17184 31346
rect 17236 31328 17264 34002
rect 17420 33998 17448 35022
rect 18328 34604 18380 34610
rect 18328 34546 18380 34552
rect 17684 34400 17736 34406
rect 17684 34342 17736 34348
rect 17696 33998 17724 34342
rect 18340 34202 18368 34546
rect 18892 34542 18920 35430
rect 19076 35290 19104 35566
rect 19156 35488 19208 35494
rect 19156 35430 19208 35436
rect 19248 35488 19300 35494
rect 19248 35430 19300 35436
rect 19168 35290 19196 35430
rect 19064 35284 19116 35290
rect 19064 35226 19116 35232
rect 19156 35284 19208 35290
rect 19156 35226 19208 35232
rect 18420 34536 18472 34542
rect 18420 34478 18472 34484
rect 18880 34536 18932 34542
rect 18880 34478 18932 34484
rect 18328 34196 18380 34202
rect 18328 34138 18380 34144
rect 18432 34134 18460 34478
rect 18788 34196 18840 34202
rect 18788 34138 18840 34144
rect 18420 34128 18472 34134
rect 18420 34070 18472 34076
rect 17408 33992 17460 33998
rect 17408 33934 17460 33940
rect 17684 33992 17736 33998
rect 17684 33934 17736 33940
rect 17592 33924 17644 33930
rect 17592 33866 17644 33872
rect 17316 33856 17368 33862
rect 17316 33798 17368 33804
rect 17328 32366 17356 33798
rect 17604 33697 17632 33866
rect 17590 33688 17646 33697
rect 17590 33623 17646 33632
rect 18800 33522 18828 34138
rect 18892 33998 18920 34478
rect 18880 33992 18932 33998
rect 18880 33934 18932 33940
rect 19076 33590 19104 35226
rect 19260 35086 19288 35430
rect 19248 35080 19300 35086
rect 19248 35022 19300 35028
rect 19720 34542 19748 35702
rect 25688 35692 25740 35698
rect 25688 35634 25740 35640
rect 28724 35692 28776 35698
rect 28724 35634 28776 35640
rect 34520 35692 34572 35698
rect 34520 35634 34572 35640
rect 25596 35624 25648 35630
rect 25596 35566 25648 35572
rect 25608 35290 25636 35566
rect 25596 35284 25648 35290
rect 25596 35226 25648 35232
rect 22192 35080 22244 35086
rect 22192 35022 22244 35028
rect 20168 35012 20220 35018
rect 20168 34954 20220 34960
rect 20180 34746 20208 34954
rect 20996 34944 21048 34950
rect 20996 34886 21048 34892
rect 21008 34746 21036 34886
rect 20168 34740 20220 34746
rect 20168 34682 20220 34688
rect 20720 34740 20772 34746
rect 20720 34682 20772 34688
rect 20996 34740 21048 34746
rect 20996 34682 21048 34688
rect 19708 34536 19760 34542
rect 19708 34478 19760 34484
rect 19248 34128 19300 34134
rect 19248 34070 19300 34076
rect 19064 33584 19116 33590
rect 19064 33526 19116 33532
rect 18696 33516 18748 33522
rect 18696 33458 18748 33464
rect 18788 33516 18840 33522
rect 18788 33458 18840 33464
rect 17776 33380 17828 33386
rect 17776 33322 17828 33328
rect 17408 33312 17460 33318
rect 17408 33254 17460 33260
rect 17420 32910 17448 33254
rect 17788 32910 17816 33322
rect 17408 32904 17460 32910
rect 17408 32846 17460 32852
rect 17776 32904 17828 32910
rect 17776 32846 17828 32852
rect 18604 32904 18656 32910
rect 18604 32846 18656 32852
rect 17684 32768 17736 32774
rect 17684 32710 17736 32716
rect 17316 32360 17368 32366
rect 17316 32302 17368 32308
rect 17328 32230 17356 32302
rect 17316 32224 17368 32230
rect 17316 32166 17368 32172
rect 17408 31680 17460 31686
rect 17408 31622 17460 31628
rect 17420 31482 17448 31622
rect 17408 31476 17460 31482
rect 17408 31418 17460 31424
rect 17592 31408 17644 31414
rect 17592 31350 17644 31356
rect 17316 31340 17368 31346
rect 17236 31300 17316 31328
rect 17132 31282 17184 31288
rect 17316 31282 17368 31288
rect 16868 30122 16896 31282
rect 17604 30598 17632 31350
rect 17696 31278 17724 32710
rect 18236 32496 18288 32502
rect 18236 32438 18288 32444
rect 18248 31958 18276 32438
rect 18236 31952 18288 31958
rect 18236 31894 18288 31900
rect 17776 31748 17828 31754
rect 17776 31690 17828 31696
rect 17788 31482 17816 31690
rect 18144 31680 18196 31686
rect 18144 31622 18196 31628
rect 17776 31476 17828 31482
rect 17776 31418 17828 31424
rect 18156 31346 18184 31622
rect 18616 31346 18644 32846
rect 18144 31340 18196 31346
rect 18144 31282 18196 31288
rect 18604 31340 18656 31346
rect 18604 31282 18656 31288
rect 17684 31272 17736 31278
rect 17684 31214 17736 31220
rect 17868 31136 17920 31142
rect 17868 31078 17920 31084
rect 17592 30592 17644 30598
rect 17592 30534 17644 30540
rect 17040 30184 17092 30190
rect 17040 30126 17092 30132
rect 16856 30116 16908 30122
rect 16856 30058 16908 30064
rect 16672 29708 16724 29714
rect 16672 29650 16724 29656
rect 16684 28082 16712 29650
rect 16672 28076 16724 28082
rect 16672 28018 16724 28024
rect 16764 28076 16816 28082
rect 16764 28018 16816 28024
rect 16776 27674 16804 28018
rect 16764 27668 16816 27674
rect 16764 27610 16816 27616
rect 16948 27532 17000 27538
rect 16948 27474 17000 27480
rect 16580 27328 16632 27334
rect 16580 27270 16632 27276
rect 16764 27328 16816 27334
rect 16764 27270 16816 27276
rect 16592 26994 16620 27270
rect 16580 26988 16632 26994
rect 16580 26930 16632 26936
rect 16776 26790 16804 27270
rect 16764 26784 16816 26790
rect 16764 26726 16816 26732
rect 16488 26580 16540 26586
rect 16488 26522 16540 26528
rect 16396 26240 16448 26246
rect 16396 26182 16448 26188
rect 16408 26042 16436 26182
rect 16396 26036 16448 26042
rect 16396 25978 16448 25984
rect 16408 25906 16436 25978
rect 16488 25968 16540 25974
rect 16488 25910 16540 25916
rect 16396 25900 16448 25906
rect 16396 25842 16448 25848
rect 16302 25800 16358 25809
rect 16302 25735 16358 25744
rect 16120 25696 16172 25702
rect 16120 25638 16172 25644
rect 16028 25492 16080 25498
rect 16028 25434 16080 25440
rect 16028 25356 16080 25362
rect 16132 25344 16160 25638
rect 16316 25498 16344 25735
rect 16304 25492 16356 25498
rect 16304 25434 16356 25440
rect 16080 25316 16160 25344
rect 16028 25298 16080 25304
rect 16132 24954 16160 25316
rect 16316 25158 16344 25434
rect 16304 25152 16356 25158
rect 16304 25094 16356 25100
rect 16120 24948 16172 24954
rect 16120 24890 16172 24896
rect 16316 24857 16344 25094
rect 16302 24848 16358 24857
rect 16302 24783 16358 24792
rect 15936 24200 15988 24206
rect 15936 24142 15988 24148
rect 15752 23792 15804 23798
rect 15752 23734 15804 23740
rect 15764 23526 15792 23734
rect 15948 23730 15976 24142
rect 15936 23724 15988 23730
rect 15936 23666 15988 23672
rect 15844 23656 15896 23662
rect 15842 23624 15844 23633
rect 15896 23624 15898 23633
rect 15842 23559 15898 23568
rect 15752 23520 15804 23526
rect 15752 23462 15804 23468
rect 15660 22976 15712 22982
rect 15660 22918 15712 22924
rect 15672 22778 15700 22918
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15764 22574 15792 23462
rect 15752 22568 15804 22574
rect 15804 22528 15884 22556
rect 15752 22510 15804 22516
rect 15752 22160 15804 22166
rect 15752 22102 15804 22108
rect 15764 21622 15792 22102
rect 15856 21894 15884 22528
rect 15948 22030 15976 23666
rect 16408 23254 16436 25842
rect 16500 25430 16528 25910
rect 16488 25424 16540 25430
rect 16488 25366 16540 25372
rect 16580 25356 16632 25362
rect 16580 25298 16632 25304
rect 16592 25158 16620 25298
rect 16776 25294 16804 26726
rect 16856 26376 16908 26382
rect 16856 26318 16908 26324
rect 16868 26042 16896 26318
rect 16856 26036 16908 26042
rect 16856 25978 16908 25984
rect 16868 25362 16896 25978
rect 16856 25356 16908 25362
rect 16856 25298 16908 25304
rect 16764 25288 16816 25294
rect 16960 25242 16988 27474
rect 17052 27130 17080 30126
rect 17408 29572 17460 29578
rect 17408 29514 17460 29520
rect 17420 29306 17448 29514
rect 17408 29300 17460 29306
rect 17408 29242 17460 29248
rect 17224 28416 17276 28422
rect 17224 28358 17276 28364
rect 17236 27334 17264 28358
rect 17316 27396 17368 27402
rect 17316 27338 17368 27344
rect 17224 27328 17276 27334
rect 17224 27270 17276 27276
rect 17040 27124 17092 27130
rect 17040 27066 17092 27072
rect 17052 26926 17080 27066
rect 17328 26994 17356 27338
rect 17500 27328 17552 27334
rect 17500 27270 17552 27276
rect 17512 27062 17540 27270
rect 17500 27056 17552 27062
rect 17500 26998 17552 27004
rect 17316 26988 17368 26994
rect 17316 26930 17368 26936
rect 17408 26988 17460 26994
rect 17408 26930 17460 26936
rect 17040 26920 17092 26926
rect 17420 26897 17448 26930
rect 17040 26862 17092 26868
rect 17406 26888 17462 26897
rect 16764 25230 16816 25236
rect 16868 25214 16988 25242
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16592 24410 16620 25094
rect 16672 24608 16724 24614
rect 16672 24550 16724 24556
rect 16580 24404 16632 24410
rect 16580 24346 16632 24352
rect 16684 24138 16712 24550
rect 16672 24132 16724 24138
rect 16672 24074 16724 24080
rect 16396 23248 16448 23254
rect 16448 23196 16528 23202
rect 16396 23190 16528 23196
rect 16028 23180 16080 23186
rect 16408 23174 16528 23190
rect 16028 23122 16080 23128
rect 16040 22642 16068 23122
rect 16212 23112 16264 23118
rect 16212 23054 16264 23060
rect 16120 23044 16172 23050
rect 16120 22986 16172 22992
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 15844 21888 15896 21894
rect 15844 21830 15896 21836
rect 15752 21616 15804 21622
rect 15752 21558 15804 21564
rect 15764 21146 15792 21558
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15856 20330 15884 21830
rect 16132 21690 16160 22986
rect 16224 22574 16252 23054
rect 16500 22642 16528 23174
rect 16764 22976 16816 22982
rect 16764 22918 16816 22924
rect 16776 22710 16804 22918
rect 16764 22704 16816 22710
rect 16764 22646 16816 22652
rect 16488 22636 16540 22642
rect 16488 22578 16540 22584
rect 16212 22568 16264 22574
rect 16212 22510 16264 22516
rect 16764 22568 16816 22574
rect 16764 22510 16816 22516
rect 16224 22409 16252 22510
rect 16210 22400 16266 22409
rect 16210 22335 16266 22344
rect 16776 22094 16804 22510
rect 16868 22234 16896 25214
rect 17052 23254 17080 26862
rect 17406 26823 17462 26832
rect 17222 26752 17278 26761
rect 17222 26687 17278 26696
rect 17130 26616 17186 26625
rect 17130 26551 17186 26560
rect 17144 26518 17172 26551
rect 17132 26512 17184 26518
rect 17132 26454 17184 26460
rect 17132 26376 17184 26382
rect 17236 26353 17264 26687
rect 17408 26512 17460 26518
rect 17408 26454 17460 26460
rect 17604 26466 17632 30534
rect 17776 27328 17828 27334
rect 17776 27270 17828 27276
rect 17788 27033 17816 27270
rect 17774 27024 17830 27033
rect 17774 26959 17830 26968
rect 17880 26790 17908 31078
rect 18156 30326 18184 31282
rect 18328 31272 18380 31278
rect 18328 31214 18380 31220
rect 18340 30870 18368 31214
rect 18328 30864 18380 30870
rect 18328 30806 18380 30812
rect 18144 30320 18196 30326
rect 18512 30320 18564 30326
rect 18144 30262 18196 30268
rect 18510 30288 18512 30297
rect 18564 30288 18566 30297
rect 18420 30252 18472 30258
rect 18510 30223 18566 30232
rect 18420 30194 18472 30200
rect 18328 30116 18380 30122
rect 18328 30058 18380 30064
rect 18340 29510 18368 30058
rect 18432 29850 18460 30194
rect 18708 30122 18736 33458
rect 19260 32502 19288 34070
rect 19616 33584 19668 33590
rect 19536 33532 19616 33538
rect 19536 33526 19668 33532
rect 19536 33510 19656 33526
rect 19536 32570 19564 33510
rect 19616 32836 19668 32842
rect 19616 32778 19668 32784
rect 19628 32570 19656 32778
rect 19524 32564 19576 32570
rect 19524 32506 19576 32512
rect 19616 32564 19668 32570
rect 19616 32506 19668 32512
rect 19248 32496 19300 32502
rect 19248 32438 19300 32444
rect 19720 31414 19748 34478
rect 20732 33522 20760 34682
rect 22204 34678 22232 35022
rect 23296 35012 23348 35018
rect 23296 34954 23348 34960
rect 24676 35012 24728 35018
rect 24676 34954 24728 34960
rect 23308 34746 23336 34954
rect 23572 34944 23624 34950
rect 23572 34886 23624 34892
rect 23584 34746 23612 34886
rect 24688 34746 24716 34954
rect 23296 34740 23348 34746
rect 23296 34682 23348 34688
rect 23572 34740 23624 34746
rect 23572 34682 23624 34688
rect 24676 34740 24728 34746
rect 24676 34682 24728 34688
rect 25320 34740 25372 34746
rect 25320 34682 25372 34688
rect 22192 34672 22244 34678
rect 22192 34614 22244 34620
rect 22560 34672 22612 34678
rect 22560 34614 22612 34620
rect 22100 34604 22152 34610
rect 22100 34546 22152 34552
rect 20812 34536 20864 34542
rect 20810 34504 20812 34513
rect 20864 34504 20866 34513
rect 20810 34439 20866 34448
rect 22112 34202 22140 34546
rect 22468 34400 22520 34406
rect 22468 34342 22520 34348
rect 22100 34196 22152 34202
rect 22100 34138 22152 34144
rect 20904 33992 20956 33998
rect 20904 33934 20956 33940
rect 20812 33856 20864 33862
rect 20812 33798 20864 33804
rect 20824 33522 20852 33798
rect 20444 33516 20496 33522
rect 20444 33458 20496 33464
rect 20720 33516 20772 33522
rect 20720 33458 20772 33464
rect 20812 33516 20864 33522
rect 20812 33458 20864 33464
rect 20456 32774 20484 33458
rect 19984 32768 20036 32774
rect 19984 32710 20036 32716
rect 20444 32768 20496 32774
rect 20444 32710 20496 32716
rect 19996 32570 20024 32710
rect 19984 32564 20036 32570
rect 19984 32506 20036 32512
rect 20444 32224 20496 32230
rect 20444 32166 20496 32172
rect 19708 31408 19760 31414
rect 19708 31350 19760 31356
rect 19248 31340 19300 31346
rect 19248 31282 19300 31288
rect 19260 30870 19288 31282
rect 19248 30864 19300 30870
rect 19248 30806 19300 30812
rect 19720 30598 19748 31350
rect 19984 31136 20036 31142
rect 19984 31078 20036 31084
rect 19800 30796 19852 30802
rect 19800 30738 19852 30744
rect 19708 30592 19760 30598
rect 19708 30534 19760 30540
rect 19720 30394 19748 30534
rect 19812 30433 19840 30738
rect 19996 30734 20024 31078
rect 19984 30728 20036 30734
rect 19984 30670 20036 30676
rect 19798 30424 19854 30433
rect 19708 30388 19760 30394
rect 19798 30359 19854 30368
rect 19708 30330 19760 30336
rect 18696 30116 18748 30122
rect 18696 30058 18748 30064
rect 19340 30048 19392 30054
rect 19340 29990 19392 29996
rect 18420 29844 18472 29850
rect 18420 29786 18472 29792
rect 19352 29646 19380 29990
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 19340 29640 19392 29646
rect 19340 29582 19392 29588
rect 18328 29504 18380 29510
rect 18328 29446 18380 29452
rect 18340 29306 18368 29446
rect 18328 29300 18380 29306
rect 18328 29242 18380 29248
rect 19260 29238 19288 29582
rect 19248 29232 19300 29238
rect 19248 29174 19300 29180
rect 19154 29064 19210 29073
rect 19720 29034 19748 30330
rect 19892 29504 19944 29510
rect 19892 29446 19944 29452
rect 19154 28999 19210 29008
rect 19708 29028 19760 29034
rect 19168 28966 19196 28999
rect 19708 28970 19760 28976
rect 19156 28960 19208 28966
rect 19156 28902 19208 28908
rect 18052 27872 18104 27878
rect 18052 27814 18104 27820
rect 18144 27872 18196 27878
rect 18144 27814 18196 27820
rect 17960 27600 18012 27606
rect 17960 27542 18012 27548
rect 17972 26926 18000 27542
rect 18064 27470 18092 27814
rect 18156 27674 18184 27814
rect 18144 27668 18196 27674
rect 18144 27610 18196 27616
rect 18052 27464 18104 27470
rect 18052 27406 18104 27412
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 17960 26920 18012 26926
rect 18064 26897 18092 26930
rect 17960 26862 18012 26868
rect 18050 26888 18106 26897
rect 18050 26823 18106 26832
rect 17776 26784 17828 26790
rect 17696 26744 17776 26772
rect 17696 26586 17724 26744
rect 17776 26726 17828 26732
rect 17868 26784 17920 26790
rect 17868 26726 17920 26732
rect 17684 26580 17736 26586
rect 17684 26522 17736 26528
rect 17776 26512 17828 26518
rect 17604 26460 17776 26466
rect 17604 26454 17828 26460
rect 17420 26364 17448 26454
rect 17604 26438 17816 26454
rect 17592 26376 17644 26382
rect 17132 26318 17184 26324
rect 17222 26344 17278 26353
rect 17144 24818 17172 26318
rect 17420 26336 17592 26364
rect 17592 26318 17644 26324
rect 17222 26279 17278 26288
rect 17224 25900 17276 25906
rect 17224 25842 17276 25848
rect 17236 25498 17264 25842
rect 17224 25492 17276 25498
rect 17224 25434 17276 25440
rect 17500 25152 17552 25158
rect 17500 25094 17552 25100
rect 17314 24848 17370 24857
rect 17132 24812 17184 24818
rect 17314 24783 17370 24792
rect 17132 24754 17184 24760
rect 17144 24410 17172 24754
rect 17328 24750 17356 24783
rect 17224 24744 17276 24750
rect 17222 24712 17224 24721
rect 17316 24744 17368 24750
rect 17276 24712 17278 24721
rect 17316 24686 17368 24692
rect 17222 24647 17278 24656
rect 17132 24404 17184 24410
rect 17132 24346 17184 24352
rect 17512 24274 17540 25094
rect 17590 24712 17646 24721
rect 17590 24647 17646 24656
rect 17604 24614 17632 24647
rect 17592 24608 17644 24614
rect 17592 24550 17644 24556
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 17040 23248 17092 23254
rect 17040 23190 17092 23196
rect 17052 23050 17080 23190
rect 17040 23044 17092 23050
rect 17040 22986 17092 22992
rect 17788 22778 17816 26438
rect 17776 22772 17828 22778
rect 17776 22714 17828 22720
rect 17224 22636 17276 22642
rect 17224 22578 17276 22584
rect 16856 22228 16908 22234
rect 16856 22170 16908 22176
rect 17236 22166 17264 22578
rect 17880 22574 17908 26726
rect 18050 26616 18106 26625
rect 18050 26551 18106 26560
rect 18064 26382 18092 26551
rect 18052 26376 18104 26382
rect 18052 26318 18104 26324
rect 18156 26314 18184 27610
rect 18972 27396 19024 27402
rect 18972 27338 19024 27344
rect 18984 27130 19012 27338
rect 18972 27124 19024 27130
rect 18972 27066 19024 27072
rect 19168 26625 19196 28902
rect 19720 28626 19748 28970
rect 19708 28620 19760 28626
rect 19708 28562 19760 28568
rect 19708 27872 19760 27878
rect 19708 27814 19760 27820
rect 19720 27402 19748 27814
rect 19708 27396 19760 27402
rect 19708 27338 19760 27344
rect 19800 26988 19852 26994
rect 19800 26930 19852 26936
rect 19154 26616 19210 26625
rect 19154 26551 19210 26560
rect 18236 26376 18288 26382
rect 18236 26318 18288 26324
rect 18144 26308 18196 26314
rect 18144 26250 18196 26256
rect 18052 25832 18104 25838
rect 18052 25774 18104 25780
rect 18064 25498 18092 25774
rect 18052 25492 18104 25498
rect 18052 25434 18104 25440
rect 18052 23724 18104 23730
rect 18052 23666 18104 23672
rect 18064 22778 18092 23666
rect 18248 23050 18276 26318
rect 18878 26072 18934 26081
rect 18878 26007 18934 26016
rect 18892 25838 18920 26007
rect 19064 25900 19116 25906
rect 19064 25842 19116 25848
rect 19616 25900 19668 25906
rect 19616 25842 19668 25848
rect 18880 25832 18932 25838
rect 18880 25774 18932 25780
rect 18328 25696 18380 25702
rect 18328 25638 18380 25644
rect 18340 25294 18368 25638
rect 19076 25498 19104 25842
rect 19154 25528 19210 25537
rect 19064 25492 19116 25498
rect 19154 25463 19156 25472
rect 19064 25434 19116 25440
rect 19208 25463 19210 25472
rect 19156 25434 19208 25440
rect 19062 25392 19118 25401
rect 19062 25327 19118 25336
rect 18328 25288 18380 25294
rect 18328 25230 18380 25236
rect 18972 25288 19024 25294
rect 18972 25230 19024 25236
rect 18328 24676 18380 24682
rect 18328 24618 18380 24624
rect 18236 23044 18288 23050
rect 18236 22986 18288 22992
rect 18340 22778 18368 24618
rect 18984 23730 19012 25230
rect 19076 23730 19104 25327
rect 19524 24948 19576 24954
rect 19524 24890 19576 24896
rect 19536 24342 19564 24890
rect 19628 24410 19656 25842
rect 19708 25220 19760 25226
rect 19708 25162 19760 25168
rect 19720 24954 19748 25162
rect 19708 24948 19760 24954
rect 19708 24890 19760 24896
rect 19812 24886 19840 26930
rect 19800 24880 19852 24886
rect 19800 24822 19852 24828
rect 19904 24410 19932 29446
rect 20260 29164 20312 29170
rect 20260 29106 20312 29112
rect 20272 28762 20300 29106
rect 20260 28756 20312 28762
rect 20260 28698 20312 28704
rect 20352 28688 20404 28694
rect 20352 28630 20404 28636
rect 20076 28076 20128 28082
rect 20076 28018 20128 28024
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 19996 26518 20024 26930
rect 19984 26512 20036 26518
rect 19984 26454 20036 26460
rect 20088 26042 20116 28018
rect 20168 28008 20220 28014
rect 20168 27950 20220 27956
rect 20180 27674 20208 27950
rect 20168 27668 20220 27674
rect 20168 27610 20220 27616
rect 20168 26988 20220 26994
rect 20168 26930 20220 26936
rect 20180 26042 20208 26930
rect 20260 26920 20312 26926
rect 20260 26862 20312 26868
rect 20272 26586 20300 26862
rect 20260 26580 20312 26586
rect 20260 26522 20312 26528
rect 20260 26444 20312 26450
rect 20260 26386 20312 26392
rect 20076 26036 20128 26042
rect 20076 25978 20128 25984
rect 20168 26036 20220 26042
rect 20168 25978 20220 25984
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 19996 25158 20024 25842
rect 19984 25152 20036 25158
rect 19984 25094 20036 25100
rect 19996 24954 20024 25094
rect 19984 24948 20036 24954
rect 19984 24890 20036 24896
rect 20088 24818 20116 25978
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 20088 24682 20116 24754
rect 20076 24676 20128 24682
rect 20076 24618 20128 24624
rect 19984 24608 20036 24614
rect 19984 24550 20036 24556
rect 20168 24608 20220 24614
rect 20168 24550 20220 24556
rect 19996 24410 20024 24550
rect 19616 24404 19668 24410
rect 19616 24346 19668 24352
rect 19892 24404 19944 24410
rect 19892 24346 19944 24352
rect 19984 24404 20036 24410
rect 19984 24346 20036 24352
rect 19524 24336 19576 24342
rect 19524 24278 19576 24284
rect 19248 24200 19300 24206
rect 19154 24168 19210 24177
rect 19248 24142 19300 24148
rect 19154 24103 19210 24112
rect 19168 23866 19196 24103
rect 19156 23860 19208 23866
rect 19156 23802 19208 23808
rect 18972 23724 19024 23730
rect 18972 23666 19024 23672
rect 19064 23724 19116 23730
rect 19064 23666 19116 23672
rect 18420 23520 18472 23526
rect 18420 23462 18472 23468
rect 18432 22778 18460 23462
rect 18984 23186 19012 23666
rect 18972 23180 19024 23186
rect 18972 23122 19024 23128
rect 18052 22772 18104 22778
rect 18052 22714 18104 22720
rect 18328 22772 18380 22778
rect 18328 22714 18380 22720
rect 18420 22772 18472 22778
rect 18420 22714 18472 22720
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 17408 22432 17460 22438
rect 17408 22374 17460 22380
rect 17420 22234 17448 22374
rect 17408 22228 17460 22234
rect 17408 22170 17460 22176
rect 18984 22166 19012 23122
rect 17224 22160 17276 22166
rect 17224 22102 17276 22108
rect 18972 22160 19024 22166
rect 18972 22102 19024 22108
rect 16776 22066 16896 22094
rect 16672 21956 16724 21962
rect 16672 21898 16724 21904
rect 16684 21690 16712 21898
rect 16120 21684 16172 21690
rect 16120 21626 16172 21632
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 15936 20392 15988 20398
rect 15936 20334 15988 20340
rect 15844 20324 15896 20330
rect 15844 20266 15896 20272
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 14924 19848 14976 19854
rect 14924 19790 14976 19796
rect 14832 19712 14884 19718
rect 14832 19654 14884 19660
rect 14844 19446 14872 19654
rect 14740 19440 14792 19446
rect 14740 19382 14792 19388
rect 14832 19440 14884 19446
rect 14832 19382 14884 19388
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14384 18970 14412 19246
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14384 18154 14412 18906
rect 14476 18426 14504 19314
rect 14660 19258 14688 19314
rect 14752 19310 14780 19382
rect 14568 19230 14688 19258
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14372 18148 14424 18154
rect 14372 18090 14424 18096
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14292 17338 14320 17478
rect 14280 17332 14332 17338
rect 14280 17274 14332 17280
rect 14188 17264 14240 17270
rect 14568 17218 14596 19230
rect 14648 17604 14700 17610
rect 14648 17546 14700 17552
rect 14660 17338 14688 17546
rect 14752 17338 14780 19246
rect 14936 18834 14964 19790
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 14936 17678 14964 18770
rect 14924 17672 14976 17678
rect 14924 17614 14976 17620
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14188 17206 14240 17212
rect 14292 17190 14596 17218
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 14004 16788 14056 16794
rect 13924 16748 14004 16776
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13174 15328 13230 15337
rect 13174 15263 13230 15272
rect 13084 14272 13136 14278
rect 13004 14232 13084 14260
rect 13084 14214 13136 14220
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 13004 12442 13032 13874
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12544 11558 12572 11766
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 11978 11047 12034 11056
rect 12440 11076 12492 11082
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 10876 10124 10928 10130
rect 10796 10084 10876 10112
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10520 9722 10548 9998
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10520 8838 10548 8978
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10704 8634 10732 9998
rect 10796 8838 10824 10084
rect 10876 10066 10928 10072
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11716 9654 11744 9862
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11072 9178 11100 9522
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 10876 8900 10928 8906
rect 10876 8842 10928 8848
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10888 8634 10916 8842
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 9876 7886 9904 8434
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 9588 7744 9640 7750
rect 9640 7692 9720 7698
rect 9588 7686 9720 7692
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8956 7410 8984 7686
rect 9600 7670 9720 7686
rect 1308 7404 1360 7410
rect 1308 7346 1360 7352
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 1320 6905 1348 7346
rect 1860 7268 1912 7274
rect 1860 7210 1912 7216
rect 1306 6896 1362 6905
rect 1306 6831 1362 6840
rect 1872 5778 1900 7210
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 9692 6866 9720 7670
rect 9876 7546 9904 7822
rect 10152 7546 10180 8434
rect 11348 8430 11376 8774
rect 11532 8430 11560 9454
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 10060 7002 10088 7346
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 10152 6798 10180 7482
rect 11532 7410 11560 8366
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11624 7002 11652 7346
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11992 6866 12020 11047
rect 12440 11018 12492 11024
rect 12440 10736 12492 10742
rect 12438 10704 12440 10713
rect 12492 10704 12494 10713
rect 12438 10639 12494 10648
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12176 10130 12204 10406
rect 12268 10130 12296 10542
rect 12544 10130 12572 11494
rect 12728 11286 12756 11494
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12820 10810 12848 11154
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 13096 9178 13124 14214
rect 13188 13462 13216 15263
rect 13740 14890 13768 15506
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 13280 13394 13308 14010
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13188 12306 13216 13126
rect 13556 12356 13584 13670
rect 13636 13456 13688 13462
rect 13636 13398 13688 13404
rect 13464 12328 13584 12356
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13176 12164 13228 12170
rect 13176 12106 13228 12112
rect 13188 11898 13216 12106
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13188 11150 13216 11834
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13372 9926 13400 11086
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13372 9722 13400 9862
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 13096 8974 13124 9114
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12360 8022 12388 8434
rect 12348 8016 12400 8022
rect 12348 7958 12400 7964
rect 12728 7546 12756 8910
rect 12820 8294 12848 8910
rect 13464 8838 13492 12328
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13556 11558 13584 11834
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13556 11150 13584 11494
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13648 10962 13676 13398
rect 13740 13326 13768 13670
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13924 12442 13952 16748
rect 14004 16730 14056 16736
rect 14200 16726 14228 17070
rect 14188 16720 14240 16726
rect 14188 16662 14240 16668
rect 14096 16108 14148 16114
rect 14096 16050 14148 16056
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 14016 14006 14044 14758
rect 14004 14000 14056 14006
rect 14004 13942 14056 13948
rect 14108 13938 14136 16050
rect 14292 15910 14320 17190
rect 14568 17134 14596 17190
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 14660 16794 14688 17138
rect 14752 16833 14780 17138
rect 14738 16824 14794 16833
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14648 16788 14700 16794
rect 14738 16759 14794 16768
rect 14648 16730 14700 16736
rect 14568 16674 14596 16730
rect 14568 16646 14688 16674
rect 14660 16590 14688 16646
rect 14740 16652 14792 16658
rect 14740 16594 14792 16600
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14568 16114 14596 16526
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14292 13938 14320 15846
rect 14752 15434 14780 16594
rect 14844 16590 14872 17478
rect 15028 16810 15056 19858
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 15658 19680 15714 19689
rect 15120 19378 15148 19654
rect 15658 19615 15714 19624
rect 15108 19372 15160 19378
rect 15108 19314 15160 19320
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15488 18766 15516 19110
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 15120 17814 15148 18158
rect 15108 17808 15160 17814
rect 15108 17750 15160 17756
rect 15108 17332 15160 17338
rect 15108 17274 15160 17280
rect 14936 16782 15056 16810
rect 14832 16584 14884 16590
rect 14832 16526 14884 16532
rect 14740 15428 14792 15434
rect 14740 15370 14792 15376
rect 14648 15020 14700 15026
rect 14648 14962 14700 14968
rect 14660 14618 14688 14962
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14568 14074 14596 14418
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14200 13394 14228 13874
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14108 12918 14136 13126
rect 14200 12986 14228 13330
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 14096 12912 14148 12918
rect 14096 12854 14148 12860
rect 14660 12753 14688 13806
rect 14646 12744 14702 12753
rect 14646 12679 14702 12688
rect 13912 12436 13964 12442
rect 13964 12406 14044 12434
rect 13912 12378 13964 12384
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13740 11150 13768 12242
rect 14016 12238 14044 12406
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13924 11354 13952 11630
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 13556 10934 13676 10962
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13188 8498 13216 8774
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12820 7954 12848 8230
rect 13464 7954 13492 8774
rect 13556 8090 13584 10934
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13832 10130 13860 10406
rect 13924 10266 13952 11018
rect 14016 11014 14044 12174
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13648 9178 13676 9998
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13464 7546 13492 7890
rect 13648 7886 13676 8366
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13832 7750 13860 10066
rect 14016 8906 14044 10950
rect 14004 8900 14056 8906
rect 14004 8842 14056 8848
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 12438 6896 12494 6905
rect 11980 6860 12032 6866
rect 12438 6831 12440 6840
rect 11980 6802 12032 6808
rect 12492 6831 12494 6840
rect 12440 6802 12492 6808
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 12452 6730 12480 6802
rect 12728 6798 12756 7482
rect 13832 7478 13860 7686
rect 14016 7546 14044 7822
rect 14200 7546 14228 8434
rect 14292 8294 14320 12174
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14660 11558 14688 11698
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14752 10742 14780 15370
rect 14936 15162 14964 16782
rect 15016 16720 15068 16726
rect 15016 16662 15068 16668
rect 15028 16046 15056 16662
rect 15120 16590 15148 17274
rect 15292 16720 15344 16726
rect 15290 16688 15292 16697
rect 15344 16688 15346 16697
rect 15290 16623 15346 16632
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15120 16250 15148 16526
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15212 16114 15240 16390
rect 15672 16250 15700 19615
rect 15948 19446 15976 20334
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 15936 19440 15988 19446
rect 15936 19382 15988 19388
rect 16304 19372 16356 19378
rect 16304 19314 16356 19320
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 16040 19174 16068 19246
rect 16028 19168 16080 19174
rect 16028 19110 16080 19116
rect 16040 18902 16068 19110
rect 16224 18970 16252 19246
rect 16316 18970 16344 19314
rect 16212 18964 16264 18970
rect 16212 18906 16264 18912
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16028 18896 16080 18902
rect 16028 18838 16080 18844
rect 15844 18624 15896 18630
rect 15844 18566 15896 18572
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15764 16794 15792 17138
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15856 16674 15884 18566
rect 15764 16646 15884 16674
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 14936 13530 14964 15098
rect 15028 14550 15056 15982
rect 15120 15638 15148 15982
rect 15108 15632 15160 15638
rect 15108 15574 15160 15580
rect 15120 15314 15148 15574
rect 15396 15502 15424 15982
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15120 15286 15240 15314
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 15016 14544 15068 14550
rect 15016 14486 15068 14492
rect 15120 13938 15148 14758
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14924 13524 14976 13530
rect 14924 13466 14976 13472
rect 14832 13388 14884 13394
rect 14832 13330 14884 13336
rect 14844 12238 14872 13330
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 14936 11354 14964 11698
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14844 10810 14872 10950
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14476 10062 14504 10202
rect 14568 10130 14596 10542
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14384 8634 14412 9590
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14476 8634 14504 8910
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14476 7546 14504 8570
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 13820 7472 13872 7478
rect 13820 7414 13872 7420
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 14188 6724 14240 6730
rect 14188 6666 14240 6672
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 14200 6458 14228 6666
rect 14568 6458 14596 7346
rect 14660 6662 14688 8910
rect 14752 7886 14780 10678
rect 14844 10130 14872 10746
rect 14832 10124 14884 10130
rect 14832 10066 14884 10072
rect 14844 9722 14872 10066
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 14936 9178 14964 9318
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 15028 8974 15056 13806
rect 15120 13394 15148 13874
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15212 12434 15240 15286
rect 15672 15162 15700 16050
rect 15764 15502 15792 16646
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15948 16182 15976 16526
rect 15936 16176 15988 16182
rect 15936 16118 15988 16124
rect 16040 15994 16068 18838
rect 16592 18290 16620 19790
rect 16684 19786 16712 20198
rect 16764 20052 16816 20058
rect 16764 19994 16816 20000
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16684 19378 16712 19450
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 15948 15966 16068 15994
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 15856 15502 15884 15846
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15672 14414 15700 15098
rect 15764 14822 15792 15438
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15660 13252 15712 13258
rect 15660 13194 15712 13200
rect 15672 12986 15700 13194
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15948 12646 15976 15966
rect 16132 15586 16160 16186
rect 16040 15558 16160 15586
rect 16040 13705 16068 15558
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16132 14958 16160 15438
rect 16224 15162 16252 16390
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 16132 14618 16160 14894
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 16026 13696 16082 13705
rect 16026 13631 16082 13640
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 16040 12986 16068 13126
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 16316 12442 16344 18022
rect 16776 17678 16804 19994
rect 16868 17746 16896 22066
rect 17040 21888 17092 21894
rect 17040 21830 17092 21836
rect 17052 21690 17080 21830
rect 17236 21690 17264 22102
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18788 21888 18840 21894
rect 18788 21830 18840 21836
rect 17040 21684 17092 21690
rect 17040 21626 17092 21632
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 18604 21684 18656 21690
rect 18604 21626 18656 21632
rect 17500 21616 17552 21622
rect 17500 21558 17552 21564
rect 17316 21480 17368 21486
rect 17316 21422 17368 21428
rect 17328 20874 17356 21422
rect 17512 20924 17540 21558
rect 18144 21548 18196 21554
rect 18144 21490 18196 21496
rect 18156 21146 18184 21490
rect 18512 21344 18564 21350
rect 18512 21286 18564 21292
rect 18144 21140 18196 21146
rect 18144 21082 18196 21088
rect 17684 20936 17736 20942
rect 17512 20896 17684 20924
rect 17316 20868 17368 20874
rect 17316 20810 17368 20816
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 17052 20058 17080 20402
rect 17224 20392 17276 20398
rect 17144 20352 17224 20380
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 17052 19446 17080 19994
rect 17040 19440 17092 19446
rect 17040 19382 17092 19388
rect 17144 19258 17172 20352
rect 17224 20334 17276 20340
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 17052 19230 17172 19258
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16960 17882 16988 18226
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16580 17060 16632 17066
rect 16580 17002 16632 17008
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 16500 16590 16528 16934
rect 16592 16590 16620 17002
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16776 16114 16804 16390
rect 16764 16108 16816 16114
rect 16764 16050 16816 16056
rect 16488 15632 16540 15638
rect 16488 15574 16540 15580
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16408 15094 16436 15302
rect 16396 15088 16448 15094
rect 16396 15030 16448 15036
rect 16500 14940 16528 15574
rect 16408 14912 16528 14940
rect 16408 14618 16436 14912
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16500 13734 16528 14758
rect 16776 14414 16804 14758
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16488 13728 16540 13734
rect 16394 13696 16450 13705
rect 16488 13670 16540 13676
rect 16394 13631 16450 13640
rect 16408 12730 16436 13631
rect 16592 13326 16620 14010
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16580 12776 16632 12782
rect 16408 12724 16580 12730
rect 16408 12718 16632 12724
rect 16408 12702 16620 12718
rect 15120 12406 15240 12434
rect 16304 12436 16356 12442
rect 15120 11150 15148 12406
rect 16304 12378 16356 12384
rect 15476 11824 15528 11830
rect 15476 11766 15528 11772
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14936 7834 14964 8230
rect 15120 7954 15148 11086
rect 15212 9586 15240 11494
rect 15488 11082 15516 11766
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 15488 10742 15516 11018
rect 15764 10810 15792 11018
rect 16132 10810 16160 11290
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 15476 10736 15528 10742
rect 15476 10678 15528 10684
rect 15488 10130 15516 10678
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15488 9586 15516 10066
rect 16040 10062 16068 10406
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15488 8566 15516 9522
rect 15568 9104 15620 9110
rect 15568 9046 15620 9052
rect 15580 8566 15608 9046
rect 16408 9042 16436 12702
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16592 11762 16620 12106
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16684 11694 16712 14214
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16776 12986 16804 13126
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16948 12912 17000 12918
rect 16948 12854 17000 12860
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16672 11688 16724 11694
rect 16670 11656 16672 11665
rect 16724 11656 16726 11665
rect 16670 11591 16726 11600
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16684 11150 16712 11494
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16776 9518 16804 10610
rect 16868 10606 16896 12582
rect 16960 11898 16988 12854
rect 17052 12238 17080 19230
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17144 18766 17172 19110
rect 17236 18834 17264 19654
rect 17604 19514 17632 20896
rect 17684 20878 17736 20884
rect 18236 19780 18288 19786
rect 18236 19722 18288 19728
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17500 19372 17552 19378
rect 17500 19314 17552 19320
rect 17512 19174 17540 19314
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 17132 18760 17184 18766
rect 17408 18760 17460 18766
rect 17132 18702 17184 18708
rect 17328 18720 17408 18748
rect 17328 18086 17356 18720
rect 17408 18702 17460 18708
rect 17512 18612 17540 19110
rect 17420 18584 17540 18612
rect 17316 18080 17368 18086
rect 17316 18022 17368 18028
rect 17132 17876 17184 17882
rect 17132 17818 17184 17824
rect 17144 17746 17172 17818
rect 17328 17746 17356 18022
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 17224 16584 17276 16590
rect 17222 16552 17224 16561
rect 17276 16552 17278 16561
rect 17222 16487 17278 16496
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17328 13530 17356 13874
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17420 13410 17448 18584
rect 17604 18578 17632 19450
rect 18144 19372 18196 19378
rect 18144 19314 18196 19320
rect 18156 19174 18184 19314
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 17682 18728 17738 18737
rect 17682 18663 17684 18672
rect 17736 18663 17738 18672
rect 17960 18692 18012 18698
rect 17684 18634 17736 18640
rect 17960 18634 18012 18640
rect 17604 18550 17724 18578
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17500 17604 17552 17610
rect 17500 17546 17552 17552
rect 17512 17202 17540 17546
rect 17604 17542 17632 17682
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17512 16114 17540 17138
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17512 15570 17540 16050
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 17512 14482 17540 15506
rect 17604 14822 17632 17478
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17512 13938 17540 14418
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17604 13462 17632 14758
rect 17328 13382 17448 13410
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 16948 11892 17000 11898
rect 16948 11834 17000 11840
rect 16948 11620 17000 11626
rect 16948 11562 17000 11568
rect 16960 11286 16988 11562
rect 16948 11280 17000 11286
rect 16948 11222 17000 11228
rect 17052 10792 17080 12174
rect 17144 11898 17172 12786
rect 17328 12170 17356 13382
rect 17696 13308 17724 18550
rect 17972 16250 18000 18634
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 18064 16794 18092 17138
rect 18052 16788 18104 16794
rect 18052 16730 18104 16736
rect 17960 16244 18012 16250
rect 18012 16204 18092 16232
rect 17960 16186 18012 16192
rect 18064 15502 18092 16204
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17972 15162 18000 15370
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17776 14884 17828 14890
rect 17776 14826 17828 14832
rect 17420 13280 17724 13308
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17144 11354 17172 11834
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 17328 11218 17356 11698
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 16960 10764 17080 10792
rect 16960 10674 16988 10764
rect 17132 10736 17184 10742
rect 17130 10704 17132 10713
rect 17184 10704 17186 10713
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 17040 10668 17092 10674
rect 17130 10639 17186 10648
rect 17040 10610 17092 10616
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 17052 10266 17080 10610
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 17420 10198 17448 13280
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 17512 11762 17540 13126
rect 17590 12880 17646 12889
rect 17590 12815 17592 12824
rect 17644 12815 17646 12824
rect 17592 12786 17644 12792
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17696 11830 17724 12174
rect 17684 11824 17736 11830
rect 17684 11766 17736 11772
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17590 11656 17646 11665
rect 17590 11591 17592 11600
rect 17644 11591 17646 11600
rect 17592 11562 17644 11568
rect 17604 11354 17632 11562
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17788 11014 17816 14826
rect 17960 13728 18012 13734
rect 17960 13670 18012 13676
rect 17972 13326 18000 13670
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17972 12918 18000 13262
rect 17960 12912 18012 12918
rect 17960 12854 18012 12860
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17880 11354 17908 11698
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 17408 10192 17460 10198
rect 17408 10134 17460 10140
rect 17420 10062 17448 10134
rect 17408 10056 17460 10062
rect 16946 10024 17002 10033
rect 17408 9998 17460 10004
rect 16946 9959 17002 9968
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16868 8838 16896 8978
rect 16960 8838 16988 9959
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 15568 8560 15620 8566
rect 15568 8502 15620 8508
rect 16960 8498 16988 8774
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15016 7880 15068 7886
rect 14936 7828 15016 7834
rect 14936 7822 15068 7828
rect 14936 7806 15056 7822
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14660 6458 14688 6598
rect 15028 6458 15056 7806
rect 15120 7546 15148 7890
rect 16960 7886 16988 8434
rect 17328 7886 17356 9862
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 17696 9178 17724 9522
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17788 8634 17816 10202
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17420 7886 17448 8570
rect 17512 7954 17540 8570
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17408 7880 17460 7886
rect 17696 7834 17724 7890
rect 17880 7886 17908 8910
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 18064 8090 18092 8434
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 17408 7822 17460 7828
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15120 7342 15148 7482
rect 15948 7342 15976 7754
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 15948 6866 15976 7278
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 16500 6798 16528 7686
rect 16960 6798 16988 7822
rect 17604 7818 17724 7834
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17592 7812 17724 7818
rect 17644 7806 17724 7812
rect 17592 7754 17644 7760
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 17328 7002 17356 7686
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17696 7002 17724 7346
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 17684 6996 17736 7002
rect 17684 6938 17736 6944
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 15028 6254 15056 6394
rect 15016 6248 15068 6254
rect 15016 6190 15068 6196
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 1308 5228 1360 5234
rect 1308 5170 1360 5176
rect 1320 5001 1348 5170
rect 1860 5024 1912 5030
rect 1306 4992 1362 5001
rect 1860 4966 1912 4972
rect 1306 4927 1362 4936
rect 1872 4826 1900 4966
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1320 3097 1348 3470
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 1306 3088 1362 3097
rect 1306 3023 1362 3032
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 18156 1193 18184 19110
rect 18248 18970 18276 19722
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 18524 18612 18552 21286
rect 18616 21010 18644 21626
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18708 20806 18736 21830
rect 18800 21078 18828 21830
rect 18984 21554 19012 22102
rect 18972 21548 19024 21554
rect 18972 21490 19024 21496
rect 18788 21072 18840 21078
rect 18788 21014 18840 21020
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18616 18766 18644 19654
rect 18708 19446 18736 20742
rect 18696 19440 18748 19446
rect 18696 19382 18748 19388
rect 18708 18834 18736 19382
rect 18696 18828 18748 18834
rect 18696 18770 18748 18776
rect 18880 18828 18932 18834
rect 18880 18770 18932 18776
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18524 18584 18644 18612
rect 18512 13456 18564 13462
rect 18512 13398 18564 13404
rect 18524 12850 18552 13398
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18432 11898 18460 12786
rect 18616 12306 18644 18584
rect 18892 18086 18920 18770
rect 18880 18080 18932 18086
rect 18880 18022 18932 18028
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18984 17202 19012 17478
rect 18972 17196 19024 17202
rect 18972 17138 19024 17144
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18892 16590 18920 16934
rect 19168 16658 19196 23802
rect 19260 23526 19288 24142
rect 19524 24132 19576 24138
rect 19524 24074 19576 24080
rect 19536 23866 19564 24074
rect 19904 24070 19932 24346
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19524 23860 19576 23866
rect 19524 23802 19576 23808
rect 19340 23792 19392 23798
rect 19340 23734 19392 23740
rect 19248 23520 19300 23526
rect 19248 23462 19300 23468
rect 19352 22778 19380 23734
rect 19536 22778 19564 23802
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19524 22772 19576 22778
rect 19524 22714 19576 22720
rect 19246 22536 19302 22545
rect 19246 22471 19302 22480
rect 19260 22438 19288 22471
rect 19248 22432 19300 22438
rect 19248 22374 19300 22380
rect 19260 22030 19288 22374
rect 20088 22030 20116 24142
rect 20180 24138 20208 24550
rect 20168 24132 20220 24138
rect 20168 24074 20220 24080
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 19260 21457 19288 21966
rect 19616 21548 19668 21554
rect 19616 21490 19668 21496
rect 19246 21448 19302 21457
rect 19246 21383 19302 21392
rect 19628 21146 19656 21490
rect 19982 21312 20038 21321
rect 19982 21247 20038 21256
rect 19616 21140 19668 21146
rect 19616 21082 19668 21088
rect 19340 21004 19392 21010
rect 19340 20946 19392 20952
rect 19352 20806 19380 20946
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19352 18902 19380 20742
rect 19996 20602 20024 21247
rect 20088 21078 20116 21966
rect 20272 21962 20300 26386
rect 20364 24750 20392 28630
rect 20456 28014 20484 32166
rect 20916 31890 20944 33934
rect 22008 33584 22060 33590
rect 22008 33526 22060 33532
rect 20996 33516 21048 33522
rect 20996 33458 21048 33464
rect 21008 32570 21036 33458
rect 21088 33312 21140 33318
rect 21088 33254 21140 33260
rect 22020 33266 22048 33526
rect 20996 32564 21048 32570
rect 20996 32506 21048 32512
rect 20904 31884 20956 31890
rect 20904 31826 20956 31832
rect 21100 31482 21128 33254
rect 22020 33238 22140 33266
rect 22112 32978 22140 33238
rect 22100 32972 22152 32978
rect 22100 32914 22152 32920
rect 21180 32836 21232 32842
rect 21180 32778 21232 32784
rect 21456 32836 21508 32842
rect 21456 32778 21508 32784
rect 21192 32570 21220 32778
rect 21272 32768 21324 32774
rect 21272 32710 21324 32716
rect 21180 32564 21232 32570
rect 21180 32506 21232 32512
rect 21284 32434 21312 32710
rect 21272 32428 21324 32434
rect 21272 32370 21324 32376
rect 21364 32428 21416 32434
rect 21364 32370 21416 32376
rect 21180 31884 21232 31890
rect 21180 31826 21232 31832
rect 21088 31476 21140 31482
rect 21088 31418 21140 31424
rect 20536 30592 20588 30598
rect 20812 30592 20864 30598
rect 20588 30540 20760 30546
rect 20536 30534 20760 30540
rect 20812 30534 20864 30540
rect 20548 30518 20760 30534
rect 20628 30184 20680 30190
rect 20628 30126 20680 30132
rect 20640 29850 20668 30126
rect 20732 30054 20760 30518
rect 20824 30394 20852 30534
rect 20812 30388 20864 30394
rect 20812 30330 20864 30336
rect 21192 30326 21220 31826
rect 21284 31822 21312 32370
rect 21272 31816 21324 31822
rect 21272 31758 21324 31764
rect 21272 31408 21324 31414
rect 21272 31350 21324 31356
rect 21284 30598 21312 31350
rect 21272 30592 21324 30598
rect 21272 30534 21324 30540
rect 21284 30394 21312 30534
rect 21272 30388 21324 30394
rect 21272 30330 21324 30336
rect 20904 30320 20956 30326
rect 20904 30262 20956 30268
rect 21180 30320 21232 30326
rect 21180 30262 21232 30268
rect 20720 30048 20772 30054
rect 20720 29990 20772 29996
rect 20536 29844 20588 29850
rect 20536 29786 20588 29792
rect 20628 29844 20680 29850
rect 20628 29786 20680 29792
rect 20548 29730 20576 29786
rect 20548 29702 20760 29730
rect 20732 28966 20760 29702
rect 20720 28960 20772 28966
rect 20720 28902 20772 28908
rect 20444 28008 20496 28014
rect 20444 27950 20496 27956
rect 20628 27872 20680 27878
rect 20628 27814 20680 27820
rect 20536 27668 20588 27674
rect 20536 27610 20588 27616
rect 20548 26994 20576 27610
rect 20536 26988 20588 26994
rect 20536 26930 20588 26936
rect 20640 26058 20668 27814
rect 20916 27674 20944 30262
rect 21376 29850 21404 32370
rect 21468 32026 21496 32778
rect 21732 32360 21784 32366
rect 21732 32302 21784 32308
rect 21456 32020 21508 32026
rect 21456 31962 21508 31968
rect 21744 31754 21772 32302
rect 22100 32020 22152 32026
rect 22100 31962 22152 31968
rect 22112 31890 22140 31962
rect 22100 31884 22152 31890
rect 22100 31826 22152 31832
rect 21560 31726 21772 31754
rect 22480 31754 22508 34342
rect 22572 33454 22600 34614
rect 23584 34490 23612 34682
rect 23756 34604 23808 34610
rect 23756 34546 23808 34552
rect 23492 34462 23612 34490
rect 23204 34400 23256 34406
rect 23204 34342 23256 34348
rect 23216 33998 23244 34342
rect 23296 34060 23348 34066
rect 23296 34002 23348 34008
rect 23204 33992 23256 33998
rect 23204 33934 23256 33940
rect 23308 33862 23336 34002
rect 23492 33998 23520 34462
rect 23768 34134 23796 34546
rect 23756 34128 23808 34134
rect 23756 34070 23808 34076
rect 23480 33992 23532 33998
rect 23480 33934 23532 33940
rect 23664 33924 23716 33930
rect 23664 33866 23716 33872
rect 22928 33856 22980 33862
rect 22926 33824 22928 33833
rect 23296 33856 23348 33862
rect 22980 33824 22982 33833
rect 23676 33833 23704 33866
rect 23296 33798 23348 33804
rect 23662 33824 23718 33833
rect 22926 33759 22982 33768
rect 23112 33516 23164 33522
rect 23112 33458 23164 33464
rect 22560 33448 22612 33454
rect 22560 33390 22612 33396
rect 22572 32842 22600 33390
rect 23124 33318 23152 33458
rect 23112 33312 23164 33318
rect 23112 33254 23164 33260
rect 22560 32836 22612 32842
rect 22560 32778 22612 32784
rect 22572 32434 22600 32778
rect 22560 32428 22612 32434
rect 22560 32370 22612 32376
rect 22836 32428 22888 32434
rect 22836 32370 22888 32376
rect 22848 32026 22876 32370
rect 22836 32020 22888 32026
rect 22836 31962 22888 31968
rect 22928 31952 22980 31958
rect 22928 31894 22980 31900
rect 22480 31726 22600 31754
rect 21364 29844 21416 29850
rect 21364 29786 21416 29792
rect 21088 29776 21140 29782
rect 21088 29718 21140 29724
rect 21100 29034 21128 29718
rect 21088 29028 21140 29034
rect 21088 28970 21140 28976
rect 21100 28558 21128 28970
rect 21088 28552 21140 28558
rect 21088 28494 21140 28500
rect 20904 27668 20956 27674
rect 20444 26036 20496 26042
rect 20444 25978 20496 25984
rect 20548 26030 20668 26058
rect 20732 27628 20904 27656
rect 20456 25294 20484 25978
rect 20444 25288 20496 25294
rect 20444 25230 20496 25236
rect 20352 24744 20404 24750
rect 20352 24686 20404 24692
rect 20444 22568 20496 22574
rect 20444 22510 20496 22516
rect 20456 22098 20484 22510
rect 20444 22092 20496 22098
rect 20444 22034 20496 22040
rect 20260 21956 20312 21962
rect 20260 21898 20312 21904
rect 20076 21072 20128 21078
rect 20076 21014 20128 21020
rect 20076 20800 20128 20806
rect 20076 20742 20128 20748
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 19432 20324 19484 20330
rect 19432 20266 19484 20272
rect 19444 19854 19472 20266
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19996 19786 20024 20538
rect 19524 19780 19576 19786
rect 19524 19722 19576 19728
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 19536 19378 19564 19722
rect 20088 19446 20116 20742
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 19536 18970 19564 19314
rect 19616 19168 19668 19174
rect 19616 19110 19668 19116
rect 19524 18964 19576 18970
rect 19524 18906 19576 18912
rect 19340 18896 19392 18902
rect 19340 18838 19392 18844
rect 19628 18154 19656 19110
rect 19616 18148 19668 18154
rect 19616 18090 19668 18096
rect 19892 17604 19944 17610
rect 19892 17546 19944 17552
rect 19904 17338 19932 17546
rect 19892 17332 19944 17338
rect 19892 17274 19944 17280
rect 19340 17264 19392 17270
rect 19340 17206 19392 17212
rect 19352 16726 19380 17206
rect 19800 17128 19852 17134
rect 19800 17070 19852 17076
rect 19340 16720 19392 16726
rect 19340 16662 19392 16668
rect 19156 16652 19208 16658
rect 19156 16594 19208 16600
rect 18880 16584 18932 16590
rect 18880 16526 18932 16532
rect 18788 16108 18840 16114
rect 18892 16096 18920 16526
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 18840 16068 18920 16096
rect 18972 16108 19024 16114
rect 18788 16050 18840 16056
rect 18972 16050 19024 16056
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 18984 15706 19012 16050
rect 19260 15858 19288 16050
rect 19352 16046 19380 16390
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19432 16040 19484 16046
rect 19432 15982 19484 15988
rect 19340 15904 19392 15910
rect 19260 15852 19340 15858
rect 19260 15846 19392 15852
rect 19260 15830 19380 15846
rect 18972 15700 19024 15706
rect 18972 15642 19024 15648
rect 18984 15162 19012 15642
rect 19352 15638 19380 15830
rect 19340 15632 19392 15638
rect 19340 15574 19392 15580
rect 19444 15502 19472 15982
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 18696 13728 18748 13734
rect 18748 13688 18828 13716
rect 18696 13670 18748 13676
rect 18800 12850 18828 13688
rect 19076 13410 19104 15438
rect 19444 14414 19472 15438
rect 19536 15026 19564 15846
rect 19524 15020 19576 15026
rect 19524 14962 19576 14968
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19168 13530 19196 13874
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 19076 13382 19196 13410
rect 19062 13016 19118 13025
rect 19062 12951 19118 12960
rect 19076 12850 19104 12951
rect 19168 12850 19196 13382
rect 19444 13326 19472 14350
rect 19708 13728 19760 13734
rect 19708 13670 19760 13676
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 18800 12714 18828 12786
rect 18788 12708 18840 12714
rect 18788 12650 18840 12656
rect 19168 12617 19196 12786
rect 19248 12776 19300 12782
rect 19248 12718 19300 12724
rect 19154 12608 19210 12617
rect 19154 12543 19210 12552
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18432 11150 18460 11834
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18326 10704 18382 10713
rect 18326 10639 18328 10648
rect 18380 10639 18382 10648
rect 18328 10610 18380 10616
rect 18420 10192 18472 10198
rect 18420 10134 18472 10140
rect 18432 10062 18460 10134
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18788 9988 18840 9994
rect 18788 9930 18840 9936
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 18340 9042 18368 9862
rect 18800 9450 18828 9930
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18800 8974 18828 9386
rect 18788 8968 18840 8974
rect 18788 8910 18840 8916
rect 18880 8968 18932 8974
rect 18880 8910 18932 8916
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 18432 7546 18460 8434
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18432 6730 18460 7482
rect 18616 6905 18644 8298
rect 18892 7410 18920 8910
rect 19168 8838 19196 12543
rect 19156 8832 19208 8838
rect 19156 8774 19208 8780
rect 19168 8634 19196 8774
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19260 8566 19288 12718
rect 19338 12336 19394 12345
rect 19444 12306 19472 13262
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 19338 12271 19340 12280
rect 19392 12271 19394 12280
rect 19432 12300 19484 12306
rect 19340 12242 19392 12248
rect 19432 12242 19484 12248
rect 19444 10742 19472 12242
rect 19536 11257 19564 12582
rect 19628 12458 19656 13330
rect 19720 13190 19748 13670
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19720 12850 19748 13126
rect 19708 12844 19760 12850
rect 19708 12786 19760 12792
rect 19708 12640 19760 12646
rect 19706 12608 19708 12617
rect 19760 12608 19762 12617
rect 19706 12543 19762 12552
rect 19628 12430 19748 12458
rect 19616 12368 19668 12374
rect 19616 12310 19668 12316
rect 19628 12102 19656 12310
rect 19616 12096 19668 12102
rect 19616 12038 19668 12044
rect 19628 11354 19656 12038
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19522 11248 19578 11257
rect 19628 11218 19656 11290
rect 19522 11183 19578 11192
rect 19616 11212 19668 11218
rect 19616 11154 19668 11160
rect 19614 11112 19670 11121
rect 19614 11047 19616 11056
rect 19668 11047 19670 11056
rect 19616 11018 19668 11024
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 19260 8362 19288 8502
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 19628 8022 19656 8230
rect 19720 8022 19748 12430
rect 19812 10062 19840 17070
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 19892 16652 19944 16658
rect 19892 16594 19944 16600
rect 19800 10056 19852 10062
rect 19800 9998 19852 10004
rect 19904 9586 19932 16594
rect 20076 16108 20128 16114
rect 20076 16050 20128 16056
rect 20088 15706 20116 16050
rect 20076 15700 20128 15706
rect 20076 15642 20128 15648
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19996 14414 20024 14758
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 20180 12102 20208 16934
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19904 8566 19932 9522
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19996 9178 20024 9318
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19892 8560 19944 8566
rect 19892 8502 19944 8508
rect 19984 8424 20036 8430
rect 20088 8412 20116 11630
rect 20036 8384 20116 8412
rect 19984 8366 20036 8372
rect 19996 8090 20024 8366
rect 20272 8090 20300 21898
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 20942 20484 21286
rect 20444 20936 20496 20942
rect 20548 20913 20576 26030
rect 20628 25968 20680 25974
rect 20628 25910 20680 25916
rect 20640 25702 20668 25910
rect 20628 25696 20680 25702
rect 20628 25638 20680 25644
rect 20444 20878 20496 20884
rect 20534 20904 20590 20913
rect 20640 20874 20668 25638
rect 20732 22030 20760 27628
rect 20904 27610 20956 27616
rect 21456 27396 21508 27402
rect 21456 27338 21508 27344
rect 20996 26920 21048 26926
rect 20994 26888 20996 26897
rect 21048 26888 21050 26897
rect 20994 26823 21050 26832
rect 21468 26586 21496 27338
rect 21456 26580 21508 26586
rect 21456 26522 21508 26528
rect 21560 26246 21588 31726
rect 21824 30728 21876 30734
rect 21824 30670 21876 30676
rect 21640 30184 21692 30190
rect 21640 30126 21692 30132
rect 21652 29102 21680 30126
rect 21836 29170 21864 30670
rect 21916 30116 21968 30122
rect 21916 30058 21968 30064
rect 21928 30002 21956 30058
rect 21928 29974 22048 30002
rect 22020 29714 22048 29974
rect 22008 29708 22060 29714
rect 22008 29650 22060 29656
rect 21824 29164 21876 29170
rect 21824 29106 21876 29112
rect 21640 29096 21692 29102
rect 21640 29038 21692 29044
rect 21836 28558 21864 29106
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 21640 27872 21692 27878
rect 21640 27814 21692 27820
rect 21652 26382 21680 27814
rect 21824 27056 21876 27062
rect 21876 27016 21956 27044
rect 21824 26998 21876 27004
rect 21928 27010 21956 27016
rect 22020 27010 22048 29650
rect 22100 29504 22152 29510
rect 22100 29446 22152 29452
rect 22376 29504 22428 29510
rect 22376 29446 22428 29452
rect 22112 29238 22140 29446
rect 22388 29238 22416 29446
rect 22100 29232 22152 29238
rect 22100 29174 22152 29180
rect 22376 29232 22428 29238
rect 22376 29174 22428 29180
rect 22284 28552 22336 28558
rect 22284 28494 22336 28500
rect 22296 28014 22324 28494
rect 22284 28008 22336 28014
rect 22284 27950 22336 27956
rect 22100 27872 22152 27878
rect 22100 27814 22152 27820
rect 22112 27470 22140 27814
rect 22100 27464 22152 27470
rect 22100 27406 22152 27412
rect 21928 26982 22048 27010
rect 21824 26852 21876 26858
rect 21824 26794 21876 26800
rect 21836 26586 21864 26794
rect 21824 26580 21876 26586
rect 21824 26522 21876 26528
rect 22020 26450 22048 26982
rect 22112 26761 22140 27406
rect 22296 27402 22324 27950
rect 22376 27668 22428 27674
rect 22376 27610 22428 27616
rect 22388 27520 22416 27610
rect 22468 27532 22520 27538
rect 22388 27492 22468 27520
rect 22284 27396 22336 27402
rect 22284 27338 22336 27344
rect 22296 26926 22324 27338
rect 22284 26920 22336 26926
rect 22284 26862 22336 26868
rect 22098 26752 22154 26761
rect 22098 26687 22154 26696
rect 22008 26444 22060 26450
rect 22008 26386 22060 26392
rect 21640 26376 21692 26382
rect 21640 26318 21692 26324
rect 21548 26240 21600 26246
rect 21548 26182 21600 26188
rect 21652 24818 21680 26318
rect 21732 26240 21784 26246
rect 21732 26182 21784 26188
rect 21744 25838 21772 26182
rect 21916 25900 21968 25906
rect 21916 25842 21968 25848
rect 21732 25832 21784 25838
rect 21928 25809 21956 25842
rect 21732 25774 21784 25780
rect 21914 25800 21970 25809
rect 21914 25735 21970 25744
rect 22020 25684 22048 26386
rect 22100 26240 22152 26246
rect 22100 26182 22152 26188
rect 22112 25702 22140 26182
rect 21928 25656 22048 25684
rect 22100 25696 22152 25702
rect 21824 25220 21876 25226
rect 21824 25162 21876 25168
rect 21836 24954 21864 25162
rect 21824 24948 21876 24954
rect 21824 24890 21876 24896
rect 21640 24812 21692 24818
rect 21640 24754 21692 24760
rect 21652 23662 21680 24754
rect 21732 24336 21784 24342
rect 21730 24304 21732 24313
rect 21784 24304 21786 24313
rect 21730 24239 21786 24248
rect 21744 23798 21772 24239
rect 21732 23792 21784 23798
rect 21732 23734 21784 23740
rect 21640 23656 21692 23662
rect 21640 23598 21692 23604
rect 21732 23520 21784 23526
rect 21732 23462 21784 23468
rect 21744 23118 21772 23462
rect 21732 23112 21784 23118
rect 21732 23054 21784 23060
rect 21928 22778 21956 25656
rect 22100 25638 22152 25644
rect 22112 25430 22140 25638
rect 22100 25424 22152 25430
rect 22100 25366 22152 25372
rect 22112 24750 22140 25366
rect 22192 25356 22244 25362
rect 22192 25298 22244 25304
rect 22100 24744 22152 24750
rect 22100 24686 22152 24692
rect 22008 24268 22060 24274
rect 22008 24210 22060 24216
rect 22020 23866 22048 24210
rect 22100 24200 22152 24206
rect 22100 24142 22152 24148
rect 22008 23860 22060 23866
rect 22008 23802 22060 23808
rect 22112 23730 22140 24142
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 21916 22772 21968 22778
rect 21916 22714 21968 22720
rect 22204 22574 22232 25298
rect 22296 25294 22324 26862
rect 22388 26518 22416 27492
rect 22468 27474 22520 27480
rect 22376 26512 22428 26518
rect 22376 26454 22428 26460
rect 22466 25800 22522 25809
rect 22572 25786 22600 31726
rect 22744 31680 22796 31686
rect 22744 31622 22796 31628
rect 22756 28422 22784 31622
rect 22836 30660 22888 30666
rect 22836 30602 22888 30608
rect 22848 30394 22876 30602
rect 22836 30388 22888 30394
rect 22836 30330 22888 30336
rect 22744 28416 22796 28422
rect 22744 28358 22796 28364
rect 22652 28076 22704 28082
rect 22652 28018 22704 28024
rect 22664 27470 22692 28018
rect 22652 27464 22704 27470
rect 22652 27406 22704 27412
rect 22836 26988 22888 26994
rect 22836 26930 22888 26936
rect 22650 26752 22706 26761
rect 22650 26687 22706 26696
rect 22522 25758 22600 25786
rect 22466 25735 22522 25744
rect 22480 25702 22508 25735
rect 22468 25696 22520 25702
rect 22468 25638 22520 25644
rect 22480 25362 22508 25638
rect 22664 25514 22692 26687
rect 22848 26586 22876 26930
rect 22940 26586 22968 31894
rect 23124 31754 23152 33254
rect 23020 31748 23072 31754
rect 23020 31690 23072 31696
rect 23112 31748 23164 31754
rect 23112 31690 23164 31696
rect 23032 31385 23060 31690
rect 23018 31376 23074 31385
rect 23018 31311 23074 31320
rect 23020 30252 23072 30258
rect 23020 30194 23072 30200
rect 23032 29510 23060 30194
rect 23020 29504 23072 29510
rect 23020 29446 23072 29452
rect 23020 28960 23072 28966
rect 23020 28902 23072 28908
rect 22836 26580 22888 26586
rect 22836 26522 22888 26528
rect 22928 26580 22980 26586
rect 22928 26522 22980 26528
rect 22744 26444 22796 26450
rect 22744 26386 22796 26392
rect 22756 26042 22784 26386
rect 22744 26036 22796 26042
rect 22744 25978 22796 25984
rect 23032 25974 23060 28902
rect 23124 28218 23152 31690
rect 23308 31686 23336 33798
rect 23662 33759 23718 33768
rect 23768 33046 23796 34070
rect 25332 33998 25360 34682
rect 25608 33998 25636 35226
rect 23848 33992 23900 33998
rect 23848 33934 23900 33940
rect 25320 33992 25372 33998
rect 25320 33934 25372 33940
rect 25596 33992 25648 33998
rect 25596 33934 25648 33940
rect 23860 33862 23888 33934
rect 23848 33856 23900 33862
rect 24124 33856 24176 33862
rect 23848 33798 23900 33804
rect 24122 33824 24124 33833
rect 24176 33824 24178 33833
rect 23756 33040 23808 33046
rect 23756 32982 23808 32988
rect 23572 32904 23624 32910
rect 23572 32846 23624 32852
rect 23296 31680 23348 31686
rect 23296 31622 23348 31628
rect 23480 31680 23532 31686
rect 23480 31622 23532 31628
rect 23388 31272 23440 31278
rect 23388 31214 23440 31220
rect 23296 31136 23348 31142
rect 23296 31078 23348 31084
rect 23204 30592 23256 30598
rect 23204 30534 23256 30540
rect 23216 30394 23244 30534
rect 23204 30388 23256 30394
rect 23204 30330 23256 30336
rect 23308 30190 23336 31078
rect 23400 30938 23428 31214
rect 23492 30938 23520 31622
rect 23584 31278 23612 32846
rect 23768 32434 23796 32982
rect 23756 32428 23808 32434
rect 23756 32370 23808 32376
rect 23768 31822 23796 32370
rect 23756 31816 23808 31822
rect 23756 31758 23808 31764
rect 23572 31272 23624 31278
rect 23572 31214 23624 31220
rect 23388 30932 23440 30938
rect 23388 30874 23440 30880
rect 23480 30932 23532 30938
rect 23480 30874 23532 30880
rect 23296 30184 23348 30190
rect 23296 30126 23348 30132
rect 23204 29640 23256 29646
rect 23204 29582 23256 29588
rect 23216 29306 23244 29582
rect 23204 29300 23256 29306
rect 23204 29242 23256 29248
rect 23308 29238 23336 30126
rect 23296 29232 23348 29238
rect 23296 29174 23348 29180
rect 23296 28960 23348 28966
rect 23296 28902 23348 28908
rect 23308 28558 23336 28902
rect 23400 28558 23428 30874
rect 23664 30728 23716 30734
rect 23664 30670 23716 30676
rect 23676 29850 23704 30670
rect 23664 29844 23716 29850
rect 23664 29786 23716 29792
rect 23572 29640 23624 29646
rect 23572 29582 23624 29588
rect 23480 29096 23532 29102
rect 23480 29038 23532 29044
rect 23492 28762 23520 29038
rect 23480 28756 23532 28762
rect 23480 28698 23532 28704
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 23388 28552 23440 28558
rect 23388 28494 23440 28500
rect 23112 28212 23164 28218
rect 23112 28154 23164 28160
rect 23296 27940 23348 27946
rect 23296 27882 23348 27888
rect 23204 27464 23256 27470
rect 23204 27406 23256 27412
rect 23216 26042 23244 27406
rect 23204 26036 23256 26042
rect 23204 25978 23256 25984
rect 23020 25968 23072 25974
rect 23020 25910 23072 25916
rect 22664 25486 22784 25514
rect 22468 25356 22520 25362
rect 22468 25298 22520 25304
rect 22284 25288 22336 25294
rect 22284 25230 22336 25236
rect 22560 25288 22612 25294
rect 22560 25230 22612 25236
rect 22284 25152 22336 25158
rect 22284 25094 22336 25100
rect 22296 24954 22324 25094
rect 22284 24948 22336 24954
rect 22284 24890 22336 24896
rect 22296 24274 22324 24890
rect 22468 24744 22520 24750
rect 22468 24686 22520 24692
rect 22376 24608 22428 24614
rect 22480 24562 22508 24686
rect 22428 24556 22508 24562
rect 22376 24550 22508 24556
rect 22388 24534 22508 24550
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 22480 24313 22508 24346
rect 22466 24304 22522 24313
rect 22284 24268 22336 24274
rect 22466 24239 22522 24248
rect 22284 24210 22336 24216
rect 22468 23860 22520 23866
rect 22468 23802 22520 23808
rect 22284 23724 22336 23730
rect 22284 23666 22336 23672
rect 22296 22982 22324 23666
rect 22480 23526 22508 23802
rect 22572 23730 22600 25230
rect 22652 24608 22704 24614
rect 22652 24550 22704 24556
rect 22664 24138 22692 24550
rect 22652 24132 22704 24138
rect 22652 24074 22704 24080
rect 22560 23724 22612 23730
rect 22560 23666 22612 23672
rect 22468 23520 22520 23526
rect 22468 23462 22520 23468
rect 22756 23254 22784 25486
rect 23112 25220 23164 25226
rect 23112 25162 23164 25168
rect 23124 24954 23152 25162
rect 23112 24948 23164 24954
rect 23112 24890 23164 24896
rect 22928 24812 22980 24818
rect 22928 24754 22980 24760
rect 23020 24812 23072 24818
rect 23020 24754 23072 24760
rect 22940 24682 22968 24754
rect 22928 24676 22980 24682
rect 22928 24618 22980 24624
rect 23032 24342 23060 24754
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 23216 24342 23244 24550
rect 23020 24336 23072 24342
rect 23020 24278 23072 24284
rect 23204 24336 23256 24342
rect 23204 24278 23256 24284
rect 23308 24206 23336 27882
rect 23492 27130 23520 28698
rect 23584 27577 23612 29582
rect 23664 29572 23716 29578
rect 23664 29514 23716 29520
rect 23676 29170 23704 29514
rect 23664 29164 23716 29170
rect 23664 29106 23716 29112
rect 23676 28762 23704 29106
rect 23664 28756 23716 28762
rect 23664 28698 23716 28704
rect 23860 27946 23888 33798
rect 24122 33759 24178 33768
rect 24400 32904 24452 32910
rect 24400 32846 24452 32852
rect 23940 32224 23992 32230
rect 23940 32166 23992 32172
rect 23952 30938 23980 32166
rect 24412 31278 24440 32846
rect 24492 32836 24544 32842
rect 24492 32778 24544 32784
rect 24504 32298 24532 32778
rect 24492 32292 24544 32298
rect 24492 32234 24544 32240
rect 25596 31476 25648 31482
rect 25596 31418 25648 31424
rect 24676 31408 24728 31414
rect 24676 31350 24728 31356
rect 24400 31272 24452 31278
rect 24400 31214 24452 31220
rect 23940 30932 23992 30938
rect 23940 30874 23992 30880
rect 24032 30048 24084 30054
rect 24032 29990 24084 29996
rect 23848 27940 23900 27946
rect 23848 27882 23900 27888
rect 23570 27568 23626 27577
rect 23570 27503 23626 27512
rect 23756 27532 23808 27538
rect 23480 27124 23532 27130
rect 23480 27066 23532 27072
rect 23480 26308 23532 26314
rect 23480 26250 23532 26256
rect 23492 24732 23520 26250
rect 23584 25906 23612 27503
rect 23756 27474 23808 27480
rect 23664 27464 23716 27470
rect 23662 27432 23664 27441
rect 23716 27432 23718 27441
rect 23662 27367 23718 27376
rect 23664 26784 23716 26790
rect 23768 26772 23796 27474
rect 23848 27328 23900 27334
rect 23848 27270 23900 27276
rect 23716 26744 23796 26772
rect 23664 26726 23716 26732
rect 23676 26382 23704 26726
rect 23664 26376 23716 26382
rect 23664 26318 23716 26324
rect 23860 26314 23888 27270
rect 23848 26308 23900 26314
rect 23848 26250 23900 26256
rect 23756 26240 23808 26246
rect 24044 26194 24072 29990
rect 24412 29714 24440 31214
rect 24688 30666 24716 31350
rect 25136 31340 25188 31346
rect 25136 31282 25188 31288
rect 25148 30938 25176 31282
rect 25228 31136 25280 31142
rect 25228 31078 25280 31084
rect 25240 30938 25268 31078
rect 25136 30932 25188 30938
rect 25136 30874 25188 30880
rect 25228 30932 25280 30938
rect 25228 30874 25280 30880
rect 25320 30796 25372 30802
rect 25320 30738 25372 30744
rect 24860 30728 24912 30734
rect 24860 30670 24912 30676
rect 24676 30660 24728 30666
rect 24676 30602 24728 30608
rect 24688 30394 24716 30602
rect 24872 30598 24900 30670
rect 24860 30592 24912 30598
rect 24860 30534 24912 30540
rect 24676 30388 24728 30394
rect 24676 30330 24728 30336
rect 24492 30320 24544 30326
rect 24492 30262 24544 30268
rect 24504 30122 24532 30262
rect 24492 30116 24544 30122
rect 24492 30058 24544 30064
rect 24400 29708 24452 29714
rect 24400 29650 24452 29656
rect 24504 29594 24532 30058
rect 25332 30054 25360 30738
rect 25608 30054 25636 31418
rect 25700 30666 25728 35634
rect 27988 35624 28040 35630
rect 27988 35566 28040 35572
rect 26056 35488 26108 35494
rect 26056 35430 26108 35436
rect 26240 35488 26292 35494
rect 27436 35488 27488 35494
rect 26240 35430 26292 35436
rect 27434 35456 27436 35465
rect 27620 35488 27672 35494
rect 27488 35456 27490 35465
rect 26068 35086 26096 35430
rect 26252 35193 26280 35430
rect 27620 35430 27672 35436
rect 27434 35391 27490 35400
rect 26238 35184 26294 35193
rect 26238 35119 26294 35128
rect 27632 35086 27660 35430
rect 28000 35290 28028 35566
rect 28736 35290 28764 35634
rect 34336 35624 34388 35630
rect 34334 35592 34336 35601
rect 34388 35592 34390 35601
rect 34334 35527 34390 35536
rect 27988 35284 28040 35290
rect 27988 35226 28040 35232
rect 28448 35284 28500 35290
rect 28448 35226 28500 35232
rect 28724 35284 28776 35290
rect 28724 35226 28776 35232
rect 26056 35080 26108 35086
rect 26056 35022 26108 35028
rect 27252 35080 27304 35086
rect 27252 35022 27304 35028
rect 27620 35080 27672 35086
rect 27620 35022 27672 35028
rect 25780 34944 25832 34950
rect 25780 34886 25832 34892
rect 25792 34746 25820 34886
rect 25780 34740 25832 34746
rect 25780 34682 25832 34688
rect 25780 34196 25832 34202
rect 25780 34138 25832 34144
rect 26332 34196 26384 34202
rect 26332 34138 26384 34144
rect 25792 33998 25820 34138
rect 25780 33992 25832 33998
rect 25780 33934 25832 33940
rect 25792 33658 25820 33934
rect 25872 33856 25924 33862
rect 25872 33798 25924 33804
rect 25780 33652 25832 33658
rect 25780 33594 25832 33600
rect 25884 32910 25912 33798
rect 25872 32904 25924 32910
rect 25872 32846 25924 32852
rect 25780 32768 25832 32774
rect 25780 32710 25832 32716
rect 26056 32768 26108 32774
rect 26056 32710 26108 32716
rect 25792 32570 25820 32710
rect 25780 32564 25832 32570
rect 25780 32506 25832 32512
rect 26068 32026 26096 32710
rect 26148 32360 26200 32366
rect 26148 32302 26200 32308
rect 26056 32020 26108 32026
rect 26056 31962 26108 31968
rect 25872 31816 25924 31822
rect 25872 31758 25924 31764
rect 25964 31816 26016 31822
rect 25964 31758 26016 31764
rect 25884 31482 25912 31758
rect 25872 31476 25924 31482
rect 25872 31418 25924 31424
rect 25976 31226 26004 31758
rect 25884 31198 26004 31226
rect 25884 30870 25912 31198
rect 25964 31136 26016 31142
rect 25964 31078 26016 31084
rect 25872 30864 25924 30870
rect 25872 30806 25924 30812
rect 25976 30734 26004 31078
rect 25964 30728 26016 30734
rect 25964 30670 26016 30676
rect 25688 30660 25740 30666
rect 25688 30602 25740 30608
rect 25780 30660 25832 30666
rect 25780 30602 25832 30608
rect 25320 30048 25372 30054
rect 25320 29990 25372 29996
rect 25596 30048 25648 30054
rect 25596 29990 25648 29996
rect 25044 29844 25096 29850
rect 25044 29786 25096 29792
rect 24412 29566 24532 29594
rect 24676 29572 24728 29578
rect 24124 28008 24176 28014
rect 24124 27950 24176 27956
rect 24136 26994 24164 27950
rect 24216 27600 24268 27606
rect 24216 27542 24268 27548
rect 24124 26988 24176 26994
rect 24124 26930 24176 26936
rect 23756 26182 23808 26188
rect 23572 25900 23624 25906
rect 23572 25842 23624 25848
rect 23768 25226 23796 26182
rect 23860 26166 24072 26194
rect 23756 25220 23808 25226
rect 23756 25162 23808 25168
rect 23664 24948 23716 24954
rect 23664 24890 23716 24896
rect 23572 24744 23624 24750
rect 23400 24704 23572 24732
rect 22928 24200 22980 24206
rect 22928 24142 22980 24148
rect 23112 24200 23164 24206
rect 23296 24200 23348 24206
rect 23164 24148 23296 24154
rect 23112 24142 23348 24148
rect 22836 23724 22888 23730
rect 22836 23666 22888 23672
rect 22848 23322 22876 23666
rect 22836 23316 22888 23322
rect 22836 23258 22888 23264
rect 22744 23248 22796 23254
rect 22744 23190 22796 23196
rect 22284 22976 22336 22982
rect 22284 22918 22336 22924
rect 22192 22568 22244 22574
rect 22192 22510 22244 22516
rect 22836 22568 22888 22574
rect 22836 22510 22888 22516
rect 20812 22432 20864 22438
rect 20812 22374 20864 22380
rect 22744 22432 22796 22438
rect 22744 22374 22796 22380
rect 20824 22094 20852 22374
rect 20824 22066 20944 22094
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20732 21486 20760 21966
rect 20916 21554 20944 22066
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 21180 21888 21232 21894
rect 21180 21830 21232 21836
rect 21192 21690 21220 21830
rect 21180 21684 21232 21690
rect 21180 21626 21232 21632
rect 22100 21684 22152 21690
rect 22100 21626 22152 21632
rect 22008 21616 22060 21622
rect 22008 21558 22060 21564
rect 20904 21548 20956 21554
rect 20824 21508 20904 21536
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20824 21146 20852 21508
rect 20904 21490 20956 21496
rect 22020 21350 22048 21558
rect 22112 21350 22140 21626
rect 22480 21554 22508 21966
rect 22756 21962 22784 22374
rect 22848 22098 22876 22510
rect 22836 22092 22888 22098
rect 22836 22034 22888 22040
rect 22744 21956 22796 21962
rect 22744 21898 22796 21904
rect 22756 21706 22784 21898
rect 22664 21678 22784 21706
rect 22284 21548 22336 21554
rect 22284 21490 22336 21496
rect 22468 21548 22520 21554
rect 22468 21490 22520 21496
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 22100 21344 22152 21350
rect 22100 21286 22152 21292
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 20534 20839 20536 20848
rect 20588 20839 20590 20848
rect 20628 20868 20680 20874
rect 20536 20810 20588 20816
rect 20628 20810 20680 20816
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20536 19780 20588 19786
rect 20536 19722 20588 19728
rect 20548 19514 20576 19722
rect 20536 19508 20588 19514
rect 20536 19450 20588 19456
rect 20640 19446 20668 19790
rect 20628 19440 20680 19446
rect 20628 19382 20680 19388
rect 20444 19304 20496 19310
rect 20444 19246 20496 19252
rect 20456 18970 20484 19246
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 20548 18766 20576 19110
rect 20640 18766 20668 19382
rect 20916 18850 20944 21286
rect 22008 21072 22060 21078
rect 22008 21014 22060 21020
rect 20994 20224 21050 20233
rect 20994 20159 21050 20168
rect 20824 18822 20944 18850
rect 20536 18760 20588 18766
rect 20536 18702 20588 18708
rect 20628 18760 20680 18766
rect 20628 18702 20680 18708
rect 20536 17264 20588 17270
rect 20536 17206 20588 17212
rect 20548 15570 20576 17206
rect 20640 16658 20668 18702
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20732 17202 20760 17478
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20536 15564 20588 15570
rect 20536 15506 20588 15512
rect 20548 15162 20576 15506
rect 20732 15434 20760 15846
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20732 15162 20760 15370
rect 20824 15366 20852 18822
rect 21008 16998 21036 20159
rect 21456 19848 21508 19854
rect 21456 19790 21508 19796
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 21284 19514 21312 19654
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 21376 19378 21404 19450
rect 21364 19372 21416 19378
rect 21364 19314 21416 19320
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 21468 16794 21496 19790
rect 21640 19304 21692 19310
rect 21640 19246 21692 19252
rect 21548 18760 21600 18766
rect 21548 18702 21600 18708
rect 21560 18630 21588 18702
rect 21652 18630 21680 19246
rect 21548 18624 21600 18630
rect 21546 18592 21548 18601
rect 21640 18624 21692 18630
rect 21600 18592 21602 18601
rect 21640 18566 21692 18572
rect 21546 18527 21602 18536
rect 21548 18420 21600 18426
rect 21548 18362 21600 18368
rect 21560 18222 21588 18362
rect 21744 18358 21772 19790
rect 21916 19508 21968 19514
rect 21916 19450 21968 19456
rect 21822 19000 21878 19009
rect 21928 18970 21956 19450
rect 21822 18935 21824 18944
rect 21876 18935 21878 18944
rect 21916 18964 21968 18970
rect 21824 18906 21876 18912
rect 21916 18906 21968 18912
rect 22020 18578 22048 21014
rect 22098 20632 22154 20641
rect 22098 20567 22154 20576
rect 22112 20534 22140 20567
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 22100 19984 22152 19990
rect 22100 19926 22152 19932
rect 22112 19854 22140 19926
rect 22100 19848 22152 19854
rect 22100 19790 22152 19796
rect 22296 19258 22324 21490
rect 22466 20496 22522 20505
rect 22664 20466 22692 21678
rect 22744 21548 22796 21554
rect 22744 21490 22796 21496
rect 22756 20806 22784 21490
rect 22744 20800 22796 20806
rect 22744 20742 22796 20748
rect 22756 20602 22784 20742
rect 22744 20596 22796 20602
rect 22744 20538 22796 20544
rect 22466 20431 22522 20440
rect 22652 20460 22704 20466
rect 22480 20398 22508 20431
rect 22652 20402 22704 20408
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22664 19922 22692 20402
rect 22652 19916 22704 19922
rect 22652 19858 22704 19864
rect 22376 19712 22428 19718
rect 22376 19654 22428 19660
rect 22744 19712 22796 19718
rect 22744 19654 22796 19660
rect 22388 19446 22416 19654
rect 22756 19514 22784 19654
rect 22744 19508 22796 19514
rect 22744 19450 22796 19456
rect 22376 19440 22428 19446
rect 22376 19382 22428 19388
rect 22296 19230 22416 19258
rect 22192 19168 22244 19174
rect 22244 19116 22324 19122
rect 22192 19110 22324 19116
rect 22204 19094 22324 19110
rect 22296 18766 22324 19094
rect 22192 18760 22244 18766
rect 22192 18702 22244 18708
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 21928 18550 22048 18578
rect 21732 18352 21784 18358
rect 21732 18294 21784 18300
rect 21548 18216 21600 18222
rect 21548 18158 21600 18164
rect 21560 17338 21588 18158
rect 21548 17332 21600 17338
rect 21548 17274 21600 17280
rect 21560 17066 21588 17274
rect 21548 17060 21600 17066
rect 21548 17002 21600 17008
rect 21456 16788 21508 16794
rect 21456 16730 21508 16736
rect 21928 16402 21956 18550
rect 22204 18426 22232 18702
rect 22192 18420 22244 18426
rect 22192 18362 22244 18368
rect 22098 18320 22154 18329
rect 22098 18255 22154 18264
rect 22112 18086 22140 18255
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 22112 17270 22140 17478
rect 22100 17264 22152 17270
rect 22100 17206 22152 17212
rect 22112 16794 22140 17206
rect 22100 16788 22152 16794
rect 22100 16730 22152 16736
rect 22204 16590 22232 18022
rect 22296 17678 22324 18702
rect 22388 17882 22416 19230
rect 22652 18896 22704 18902
rect 22652 18838 22704 18844
rect 22664 18426 22692 18838
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22652 18420 22704 18426
rect 22652 18362 22704 18368
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22284 17672 22336 17678
rect 22284 17614 22336 17620
rect 22296 17082 22324 17614
rect 22480 17610 22508 18362
rect 22468 17604 22520 17610
rect 22468 17546 22520 17552
rect 22664 17338 22692 18362
rect 22744 18216 22796 18222
rect 22744 18158 22796 18164
rect 22756 17542 22784 18158
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 22848 17354 22876 22034
rect 22940 21690 22968 24142
rect 23124 24126 23336 24142
rect 23204 24064 23256 24070
rect 23204 24006 23256 24012
rect 23216 23730 23244 24006
rect 23204 23724 23256 23730
rect 23204 23666 23256 23672
rect 23400 23254 23428 24704
rect 23572 24686 23624 24692
rect 23480 24200 23532 24206
rect 23480 24142 23532 24148
rect 23388 23248 23440 23254
rect 23388 23190 23440 23196
rect 23492 22982 23520 24142
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23584 23186 23612 24006
rect 23572 23180 23624 23186
rect 23572 23122 23624 23128
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23584 22506 23612 23122
rect 23572 22500 23624 22506
rect 23572 22442 23624 22448
rect 23676 22166 23704 24890
rect 23768 24750 23796 25162
rect 23756 24744 23808 24750
rect 23756 24686 23808 24692
rect 23768 24410 23796 24686
rect 23756 24404 23808 24410
rect 23756 24346 23808 24352
rect 23860 24290 23888 26166
rect 24136 25906 24164 26930
rect 24228 26790 24256 27542
rect 24216 26784 24268 26790
rect 24216 26726 24268 26732
rect 24124 25900 24176 25906
rect 24124 25842 24176 25848
rect 23940 25152 23992 25158
rect 23940 25094 23992 25100
rect 23952 24800 23980 25094
rect 24032 24812 24084 24818
rect 23952 24772 24032 24800
rect 24032 24754 24084 24760
rect 24308 24812 24360 24818
rect 24308 24754 24360 24760
rect 24032 24608 24084 24614
rect 24032 24550 24084 24556
rect 23768 24262 23888 24290
rect 23768 24206 23796 24262
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 23848 24200 23900 24206
rect 23848 24142 23900 24148
rect 23860 23866 23888 24142
rect 24044 24070 24072 24550
rect 24032 24064 24084 24070
rect 24032 24006 24084 24012
rect 23848 23860 23900 23866
rect 23848 23802 23900 23808
rect 23940 22976 23992 22982
rect 23940 22918 23992 22924
rect 23756 22636 23808 22642
rect 23756 22578 23808 22584
rect 23664 22160 23716 22166
rect 23664 22102 23716 22108
rect 23386 21992 23442 22001
rect 23386 21927 23442 21936
rect 23400 21894 23428 21927
rect 23676 21894 23704 22102
rect 23020 21888 23072 21894
rect 23020 21830 23072 21836
rect 23388 21888 23440 21894
rect 23388 21830 23440 21836
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 22928 21684 22980 21690
rect 22928 21626 22980 21632
rect 23032 21554 23060 21830
rect 23020 21548 23072 21554
rect 23020 21490 23072 21496
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 23492 21010 23520 21286
rect 23480 21004 23532 21010
rect 23480 20946 23532 20952
rect 22928 20868 22980 20874
rect 22928 20810 22980 20816
rect 22940 20602 22968 20810
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 23676 20262 23704 20742
rect 23768 20534 23796 22578
rect 23848 21072 23900 21078
rect 23848 21014 23900 21020
rect 23860 20942 23888 21014
rect 23848 20936 23900 20942
rect 23848 20878 23900 20884
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23572 20256 23624 20262
rect 23572 20198 23624 20204
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23584 19990 23612 20198
rect 23572 19984 23624 19990
rect 23572 19926 23624 19932
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23296 19916 23348 19922
rect 23296 19858 23348 19864
rect 23216 19718 23244 19858
rect 23204 19712 23256 19718
rect 23202 19680 23204 19689
rect 23256 19680 23258 19689
rect 23202 19615 23258 19624
rect 23112 19304 23164 19310
rect 23112 19246 23164 19252
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 22928 18352 22980 18358
rect 22928 18294 22980 18300
rect 22652 17332 22704 17338
rect 22652 17274 22704 17280
rect 22756 17326 22876 17354
rect 22376 17128 22428 17134
rect 22296 17076 22376 17082
rect 22296 17070 22428 17076
rect 22296 17054 22416 17070
rect 22296 16590 22324 17054
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22192 16584 22244 16590
rect 22192 16526 22244 16532
rect 22284 16584 22336 16590
rect 22284 16526 22336 16532
rect 22100 16448 22152 16454
rect 21928 16374 22048 16402
rect 22100 16390 22152 16396
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 21008 15366 21036 15506
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 20536 15156 20588 15162
rect 20536 15098 20588 15104
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20548 14822 20576 14894
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20548 13258 20576 14758
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 20536 13252 20588 13258
rect 20536 13194 20588 13200
rect 20640 12714 20668 14214
rect 20824 12714 20852 15302
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 21088 15020 21140 15026
rect 21088 14962 21140 14968
rect 20916 14618 20944 14962
rect 20904 14612 20956 14618
rect 20904 14554 20956 14560
rect 20904 14340 20956 14346
rect 20904 14282 20956 14288
rect 20916 12850 20944 14282
rect 21100 14278 21128 14962
rect 21088 14272 21140 14278
rect 21088 14214 21140 14220
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 21008 12918 21036 13262
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 20628 12708 20680 12714
rect 20628 12650 20680 12656
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20916 12374 20944 12786
rect 21100 12442 21128 12786
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 20904 12368 20956 12374
rect 20904 12310 20956 12316
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20352 12164 20404 12170
rect 20352 12106 20404 12112
rect 20364 11898 20392 12106
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20352 11620 20404 11626
rect 20352 11562 20404 11568
rect 20364 10674 20392 11562
rect 20732 11558 20760 11834
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20628 11008 20680 11014
rect 20628 10950 20680 10956
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20364 10130 20392 10610
rect 20640 10606 20668 10950
rect 20628 10600 20680 10606
rect 20548 10560 20628 10588
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20352 9648 20404 9654
rect 20350 9616 20352 9625
rect 20404 9616 20406 9625
rect 20350 9551 20406 9560
rect 20548 9518 20576 10560
rect 20628 10542 20680 10548
rect 20824 10470 20852 12242
rect 21008 11354 21036 12378
rect 21100 11898 21128 12378
rect 21272 12368 21324 12374
rect 21272 12310 21324 12316
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 21088 10464 21140 10470
rect 21088 10406 21140 10412
rect 20628 9988 20680 9994
rect 20628 9930 20680 9936
rect 20640 9722 20668 9930
rect 20996 9920 21048 9926
rect 20996 9862 21048 9868
rect 21008 9722 21036 9862
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20996 9716 21048 9722
rect 20996 9658 21048 9664
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20536 9512 20588 9518
rect 20364 9472 20536 9500
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 20260 8084 20312 8090
rect 20260 8026 20312 8032
rect 19616 8016 19668 8022
rect 19616 7958 19668 7964
rect 19708 8016 19760 8022
rect 19708 7958 19760 7964
rect 19628 7750 19656 7958
rect 19616 7744 19668 7750
rect 19616 7686 19668 7692
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18602 6896 18658 6905
rect 18892 6866 18920 7346
rect 18602 6831 18658 6840
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 19720 6798 19748 7958
rect 19996 7954 20024 8026
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 20272 7886 20300 8026
rect 20364 7886 20392 9472
rect 20536 9454 20588 9460
rect 20626 9072 20682 9081
rect 20626 9007 20682 9016
rect 20640 8838 20668 9007
rect 20732 8974 20760 9590
rect 20996 9512 21048 9518
rect 20996 9454 21048 9460
rect 21008 9042 21036 9454
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 20996 9036 21048 9042
rect 20996 8978 21048 8984
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20824 8566 20852 8978
rect 20812 8560 20864 8566
rect 20812 8502 20864 8508
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20444 7948 20496 7954
rect 20444 7890 20496 7896
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 20364 7410 20392 7822
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 20456 7342 20484 7890
rect 20640 7546 20668 8434
rect 20732 8276 20760 8434
rect 21100 8430 21128 10406
rect 21284 9674 21312 12310
rect 21376 11694 21404 15438
rect 21468 15162 21496 16050
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 21836 15162 21864 15370
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21456 15156 21508 15162
rect 21456 15098 21508 15104
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21732 15020 21784 15026
rect 21732 14962 21784 14968
rect 21744 14657 21772 14962
rect 21730 14648 21786 14657
rect 21730 14583 21732 14592
rect 21784 14583 21786 14592
rect 21732 14554 21784 14560
rect 21732 13796 21784 13802
rect 21732 13738 21784 13744
rect 21744 12850 21772 13738
rect 21824 13252 21876 13258
rect 21824 13194 21876 13200
rect 21732 12844 21784 12850
rect 21732 12786 21784 12792
rect 21836 12442 21864 13194
rect 21824 12436 21876 12442
rect 21824 12378 21876 12384
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21928 11370 21956 15302
rect 22020 14618 22048 16374
rect 22112 16250 22140 16390
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22296 16182 22324 16526
rect 22388 16250 22416 16934
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 22468 16244 22520 16250
rect 22468 16186 22520 16192
rect 22284 16176 22336 16182
rect 22190 16144 22246 16153
rect 22284 16118 22336 16124
rect 22480 16114 22508 16186
rect 22190 16079 22192 16088
rect 22244 16079 22246 16088
rect 22468 16108 22520 16114
rect 22192 16050 22244 16056
rect 22468 16050 22520 16056
rect 22480 15638 22508 16050
rect 22560 16040 22612 16046
rect 22560 15982 22612 15988
rect 22572 15706 22600 15982
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22468 15632 22520 15638
rect 22466 15600 22468 15609
rect 22520 15600 22522 15609
rect 22466 15535 22522 15544
rect 22572 15162 22600 15642
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22664 15026 22692 17274
rect 22652 15020 22704 15026
rect 22652 14962 22704 14968
rect 22468 14952 22520 14958
rect 22468 14894 22520 14900
rect 22480 14822 22508 14894
rect 22468 14816 22520 14822
rect 22468 14758 22520 14764
rect 22008 14612 22060 14618
rect 22008 14554 22060 14560
rect 22020 12238 22048 14554
rect 22480 14550 22508 14758
rect 22468 14544 22520 14550
rect 22468 14486 22520 14492
rect 22376 14408 22428 14414
rect 22376 14350 22428 14356
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22112 12442 22140 13670
rect 22192 13456 22244 13462
rect 22192 13398 22244 13404
rect 22204 12918 22232 13398
rect 22192 12912 22244 12918
rect 22192 12854 22244 12860
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22112 12306 22140 12378
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 22204 12238 22232 12854
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 21732 11348 21784 11354
rect 21928 11342 22048 11370
rect 22112 11354 22140 11698
rect 21732 11290 21784 11296
rect 21744 10674 21772 11290
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 21732 10668 21784 10674
rect 21732 10610 21784 10616
rect 21376 9926 21404 10610
rect 21916 10600 21968 10606
rect 21836 10560 21916 10588
rect 21836 10470 21864 10560
rect 21916 10542 21968 10548
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21192 9646 21312 9674
rect 21192 8430 21220 9646
rect 21836 9518 21864 10406
rect 21916 9988 21968 9994
rect 21916 9930 21968 9936
rect 21824 9512 21876 9518
rect 21824 9454 21876 9460
rect 21362 9208 21418 9217
rect 21362 9143 21418 9152
rect 21824 9172 21876 9178
rect 21376 9058 21404 9143
rect 21824 9114 21876 9120
rect 21284 9042 21404 9058
rect 21836 9042 21864 9114
rect 21272 9036 21404 9042
rect 21324 9030 21404 9036
rect 21272 8978 21324 8984
rect 21272 8900 21324 8906
rect 21272 8842 21324 8848
rect 21088 8424 21140 8430
rect 21088 8366 21140 8372
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 21192 8276 21220 8366
rect 20732 8248 21220 8276
rect 20732 7818 20760 8248
rect 21284 7954 21312 8842
rect 21376 8294 21404 9030
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 21732 8968 21784 8974
rect 21732 8910 21784 8916
rect 21548 8832 21600 8838
rect 21548 8774 21600 8780
rect 21560 8498 21588 8774
rect 21652 8673 21680 8910
rect 21638 8664 21694 8673
rect 21744 8634 21772 8910
rect 21638 8599 21694 8608
rect 21732 8628 21784 8634
rect 21548 8492 21600 8498
rect 21548 8434 21600 8440
rect 21548 8356 21600 8362
rect 21652 8344 21680 8599
rect 21732 8570 21784 8576
rect 21928 8498 21956 9930
rect 22020 9178 22048 11342
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22100 11212 22152 11218
rect 22100 11154 22152 11160
rect 22112 11082 22140 11154
rect 22100 11076 22152 11082
rect 22100 11018 22152 11024
rect 22112 9382 22140 11018
rect 22296 10266 22324 13874
rect 22388 13870 22416 14350
rect 22376 13864 22428 13870
rect 22376 13806 22428 13812
rect 22388 13394 22416 13806
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22388 12434 22416 13330
rect 22560 12776 22612 12782
rect 22560 12718 22612 12724
rect 22572 12434 22600 12718
rect 22756 12714 22784 17326
rect 22940 16114 22968 18294
rect 23032 18222 23060 18566
rect 23020 18216 23072 18222
rect 23020 18158 23072 18164
rect 23124 17202 23152 19246
rect 23308 18816 23336 19858
rect 23848 19780 23900 19786
rect 23848 19722 23900 19728
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23676 19446 23704 19654
rect 23664 19440 23716 19446
rect 23664 19382 23716 19388
rect 23756 19372 23808 19378
rect 23756 19314 23808 19320
rect 23768 18970 23796 19314
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23756 18964 23808 18970
rect 23756 18906 23808 18912
rect 23216 18788 23336 18816
rect 23216 18426 23244 18788
rect 23296 18692 23348 18698
rect 23296 18634 23348 18640
rect 23308 18426 23336 18634
rect 23676 18426 23704 18906
rect 23768 18426 23796 18906
rect 23860 18902 23888 19722
rect 23848 18896 23900 18902
rect 23848 18838 23900 18844
rect 23204 18420 23256 18426
rect 23204 18362 23256 18368
rect 23296 18420 23348 18426
rect 23296 18362 23348 18368
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23756 18420 23808 18426
rect 23756 18362 23808 18368
rect 23952 18329 23980 22918
rect 24044 22098 24072 24006
rect 24320 23866 24348 24754
rect 24308 23860 24360 23866
rect 24308 23802 24360 23808
rect 24320 23118 24348 23802
rect 24308 23112 24360 23118
rect 24308 23054 24360 23060
rect 24032 22092 24084 22098
rect 24032 22034 24084 22040
rect 24308 22024 24360 22030
rect 24308 21966 24360 21972
rect 24032 21888 24084 21894
rect 24032 21830 24084 21836
rect 24044 21554 24072 21830
rect 24216 21684 24268 21690
rect 24216 21626 24268 21632
rect 24032 21548 24084 21554
rect 24032 21490 24084 21496
rect 24122 21176 24178 21185
rect 24122 21111 24178 21120
rect 24136 21078 24164 21111
rect 24124 21072 24176 21078
rect 24124 21014 24176 21020
rect 24228 20466 24256 21626
rect 24320 21593 24348 21966
rect 24306 21584 24362 21593
rect 24306 21519 24362 21528
rect 24308 21412 24360 21418
rect 24308 21354 24360 21360
rect 24320 20942 24348 21354
rect 24308 20936 24360 20942
rect 24308 20878 24360 20884
rect 24308 20800 24360 20806
rect 24412 20754 24440 29566
rect 24676 29514 24728 29520
rect 24688 29306 24716 29514
rect 25056 29306 25084 29786
rect 24676 29300 24728 29306
rect 24676 29242 24728 29248
rect 25044 29300 25096 29306
rect 25044 29242 25096 29248
rect 24768 28212 24820 28218
rect 24768 28154 24820 28160
rect 24584 26988 24636 26994
rect 24584 26930 24636 26936
rect 24596 26586 24624 26930
rect 24584 26580 24636 26586
rect 24584 26522 24636 26528
rect 24584 25152 24636 25158
rect 24584 25094 24636 25100
rect 24492 24404 24544 24410
rect 24492 24346 24544 24352
rect 24360 20748 24440 20754
rect 24308 20742 24440 20748
rect 24320 20726 24440 20742
rect 24032 20460 24084 20466
rect 24032 20402 24084 20408
rect 24216 20460 24268 20466
rect 24216 20402 24268 20408
rect 24044 20058 24072 20402
rect 24124 20392 24176 20398
rect 24124 20334 24176 20340
rect 24032 20052 24084 20058
rect 24032 19994 24084 20000
rect 24032 19712 24084 19718
rect 24032 19654 24084 19660
rect 24044 19242 24072 19654
rect 24136 19514 24164 20334
rect 24320 20262 24348 20726
rect 24400 20596 24452 20602
rect 24400 20538 24452 20544
rect 24412 20369 24440 20538
rect 24398 20360 24454 20369
rect 24398 20295 24454 20304
rect 24308 20256 24360 20262
rect 24308 20198 24360 20204
rect 24124 19508 24176 19514
rect 24124 19450 24176 19456
rect 24504 19258 24532 24346
rect 24032 19236 24084 19242
rect 24032 19178 24084 19184
rect 24228 19230 24532 19258
rect 23938 18320 23994 18329
rect 23938 18255 23994 18264
rect 23952 17542 23980 18255
rect 23940 17536 23992 17542
rect 23940 17478 23992 17484
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 23112 17196 23164 17202
rect 23112 17138 23164 17144
rect 23388 17196 23440 17202
rect 23388 17138 23440 17144
rect 22928 16108 22980 16114
rect 22928 16050 22980 16056
rect 23124 15910 23152 17138
rect 23400 16522 23428 17138
rect 23940 17128 23992 17134
rect 23940 17070 23992 17076
rect 24032 17128 24084 17134
rect 24032 17070 24084 17076
rect 23480 16992 23532 16998
rect 23480 16934 23532 16940
rect 23848 16992 23900 16998
rect 23848 16934 23900 16940
rect 23492 16590 23520 16934
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 23388 16516 23440 16522
rect 23388 16458 23440 16464
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 22928 15564 22980 15570
rect 22848 15524 22928 15552
rect 22848 13190 22876 15524
rect 22928 15506 22980 15512
rect 22836 13184 22888 13190
rect 22836 13126 22888 13132
rect 22744 12708 22796 12714
rect 22744 12650 22796 12656
rect 22756 12442 22784 12650
rect 22744 12436 22796 12442
rect 22388 12406 22508 12434
rect 22572 12406 22692 12434
rect 22480 12238 22508 12406
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22480 11830 22508 12174
rect 22664 12102 22692 12406
rect 22744 12378 22796 12384
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22468 11824 22520 11830
rect 22468 11766 22520 11772
rect 22560 11552 22612 11558
rect 22664 11506 22692 12038
rect 22612 11500 22692 11506
rect 22560 11494 22692 11500
rect 22572 11478 22692 11494
rect 22468 11144 22520 11150
rect 22468 11086 22520 11092
rect 22376 11008 22428 11014
rect 22376 10950 22428 10956
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22388 10062 22416 10950
rect 22480 10130 22508 11086
rect 22664 11082 22692 11478
rect 22652 11076 22704 11082
rect 22652 11018 22704 11024
rect 22468 10124 22520 10130
rect 22468 10066 22520 10072
rect 22376 10056 22428 10062
rect 22376 9998 22428 10004
rect 22560 10056 22612 10062
rect 22560 9998 22612 10004
rect 22572 9722 22600 9998
rect 22560 9716 22612 9722
rect 22560 9658 22612 9664
rect 22468 9648 22520 9654
rect 22468 9590 22520 9596
rect 22376 9580 22428 9586
rect 22376 9522 22428 9528
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 22008 9172 22060 9178
rect 22008 9114 22060 9120
rect 22006 9072 22062 9081
rect 22388 9042 22416 9522
rect 22480 9489 22508 9590
rect 22466 9480 22522 9489
rect 22466 9415 22522 9424
rect 22006 9007 22008 9016
rect 22060 9007 22062 9016
rect 22376 9036 22428 9042
rect 22008 8978 22060 8984
rect 22376 8978 22428 8984
rect 22100 8832 22152 8838
rect 22284 8832 22336 8838
rect 22100 8774 22152 8780
rect 22282 8800 22284 8809
rect 22468 8832 22520 8838
rect 22336 8800 22338 8809
rect 22112 8634 22140 8774
rect 22468 8774 22520 8780
rect 22282 8735 22338 8744
rect 22480 8673 22508 8774
rect 22466 8664 22522 8673
rect 22100 8628 22152 8634
rect 22466 8599 22522 8608
rect 22100 8570 22152 8576
rect 21916 8492 21968 8498
rect 21916 8434 21968 8440
rect 22192 8424 22244 8430
rect 22192 8366 22244 8372
rect 21600 8316 21680 8344
rect 21916 8356 21968 8362
rect 21548 8298 21600 8304
rect 21916 8298 21968 8304
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 21928 8022 21956 8298
rect 22204 8090 22232 8366
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 21916 8016 21968 8022
rect 21916 7958 21968 7964
rect 21272 7948 21324 7954
rect 21272 7890 21324 7896
rect 20720 7812 20772 7818
rect 20720 7754 20772 7760
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20444 7336 20496 7342
rect 20444 7278 20496 7284
rect 20456 7018 20484 7278
rect 20640 7274 20668 7482
rect 20628 7268 20680 7274
rect 20628 7210 20680 7216
rect 20364 7002 20484 7018
rect 20352 6996 20484 7002
rect 20404 6990 20484 6996
rect 20352 6938 20404 6944
rect 19708 6792 19760 6798
rect 19708 6734 19760 6740
rect 20824 6730 20852 7686
rect 21284 7002 21312 7890
rect 21824 7744 21876 7750
rect 21824 7686 21876 7692
rect 21836 7546 21864 7686
rect 21928 7546 21956 7958
rect 22204 7750 22232 8026
rect 22480 7818 22508 8599
rect 22572 8498 22600 9658
rect 22652 9648 22704 9654
rect 22650 9616 22652 9625
rect 22704 9616 22706 9625
rect 22650 9551 22706 9560
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22664 9178 22692 9318
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 22742 9072 22798 9081
rect 22742 9007 22798 9016
rect 22652 8900 22704 8906
rect 22652 8842 22704 8848
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 22468 7812 22520 7818
rect 22468 7754 22520 7760
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 21916 7540 21968 7546
rect 21916 7482 21968 7488
rect 21548 7404 21600 7410
rect 21548 7346 21600 7352
rect 21560 7206 21588 7346
rect 22664 7342 22692 8842
rect 22756 8634 22784 9007
rect 22848 8634 22876 13126
rect 22928 12232 22980 12238
rect 22928 12174 22980 12180
rect 22940 11218 22968 12174
rect 22928 11212 22980 11218
rect 22928 11154 22980 11160
rect 23124 10849 23152 15846
rect 23572 15700 23624 15706
rect 23572 15642 23624 15648
rect 23584 15162 23612 15642
rect 23572 15156 23624 15162
rect 23572 15098 23624 15104
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 23204 14816 23256 14822
rect 23204 14758 23256 14764
rect 23110 10840 23166 10849
rect 23110 10775 23166 10784
rect 22926 10568 22982 10577
rect 22926 10503 22982 10512
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 22836 8628 22888 8634
rect 22836 8570 22888 8576
rect 22756 7546 22784 8570
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22652 7336 22704 7342
rect 22652 7278 22704 7284
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 18420 6724 18472 6730
rect 18420 6666 18472 6672
rect 20812 6724 20864 6730
rect 20812 6666 20864 6672
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 21100 6322 21128 6598
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 21560 3398 21588 7142
rect 22756 7002 22784 7482
rect 22744 6996 22796 7002
rect 22744 6938 22796 6944
rect 22848 6798 22876 8570
rect 22940 8430 22968 10503
rect 23216 10146 23244 14758
rect 23388 13184 23440 13190
rect 23388 13126 23440 13132
rect 23400 12850 23428 13126
rect 23296 12844 23348 12850
rect 23296 12786 23348 12792
rect 23388 12844 23440 12850
rect 23388 12786 23440 12792
rect 23308 11626 23336 12786
rect 23400 12753 23428 12786
rect 23386 12744 23442 12753
rect 23386 12679 23442 12688
rect 23492 12322 23520 14962
rect 23860 13326 23888 16934
rect 23952 16726 23980 17070
rect 23940 16720 23992 16726
rect 23940 16662 23992 16668
rect 24044 16658 24072 17070
rect 24032 16652 24084 16658
rect 24032 16594 24084 16600
rect 23940 16516 23992 16522
rect 23940 16458 23992 16464
rect 23952 15570 23980 16458
rect 24044 15570 24072 16594
rect 24136 15706 24164 17478
rect 24228 15706 24256 19230
rect 24400 19168 24452 19174
rect 24400 19110 24452 19116
rect 24308 16992 24360 16998
rect 24308 16934 24360 16940
rect 24320 16114 24348 16934
rect 24412 16658 24440 19110
rect 24596 19009 24624 25094
rect 24780 24818 24808 28154
rect 25332 26330 25360 29990
rect 25504 29640 25556 29646
rect 25504 29582 25556 29588
rect 25516 27062 25544 29582
rect 25700 29306 25728 30602
rect 25792 30394 25820 30602
rect 25964 30592 26016 30598
rect 25964 30534 26016 30540
rect 25780 30388 25832 30394
rect 25780 30330 25832 30336
rect 25688 29300 25740 29306
rect 25688 29242 25740 29248
rect 25596 28076 25648 28082
rect 25596 28018 25648 28024
rect 25608 27674 25636 28018
rect 25596 27668 25648 27674
rect 25596 27610 25648 27616
rect 25504 27056 25556 27062
rect 25504 26998 25556 27004
rect 25412 26784 25464 26790
rect 25412 26726 25464 26732
rect 25424 26518 25452 26726
rect 25516 26518 25544 26998
rect 25412 26512 25464 26518
rect 25412 26454 25464 26460
rect 25504 26512 25556 26518
rect 25504 26454 25556 26460
rect 25596 26376 25648 26382
rect 25332 26302 25452 26330
rect 25596 26318 25648 26324
rect 25320 26240 25372 26246
rect 25320 26182 25372 26188
rect 24860 25900 24912 25906
rect 24860 25842 24912 25848
rect 24872 25498 24900 25842
rect 25332 25770 25360 26182
rect 25320 25764 25372 25770
rect 25320 25706 25372 25712
rect 25228 25696 25280 25702
rect 25228 25638 25280 25644
rect 24860 25492 24912 25498
rect 24860 25434 24912 25440
rect 24952 25288 25004 25294
rect 24952 25230 25004 25236
rect 24768 24812 24820 24818
rect 24688 24772 24768 24800
rect 24688 23866 24716 24772
rect 24768 24754 24820 24760
rect 24768 24064 24820 24070
rect 24768 24006 24820 24012
rect 24860 24064 24912 24070
rect 24860 24006 24912 24012
rect 24676 23860 24728 23866
rect 24676 23802 24728 23808
rect 24780 23730 24808 24006
rect 24768 23724 24820 23730
rect 24768 23666 24820 23672
rect 24674 21584 24730 21593
rect 24674 21519 24730 21528
rect 24582 19000 24638 19009
rect 24582 18935 24638 18944
rect 24688 18086 24716 21519
rect 24780 18154 24808 23666
rect 24872 23050 24900 24006
rect 24964 23118 24992 25230
rect 25240 25226 25268 25638
rect 25228 25220 25280 25226
rect 25228 25162 25280 25168
rect 25332 25158 25360 25706
rect 25320 25152 25372 25158
rect 25320 25094 25372 25100
rect 25332 24206 25360 25094
rect 25320 24200 25372 24206
rect 25320 24142 25372 24148
rect 24952 23112 25004 23118
rect 24952 23054 25004 23060
rect 24860 23044 24912 23050
rect 24860 22986 24912 22992
rect 24964 22642 24992 23054
rect 24952 22636 25004 22642
rect 24952 22578 25004 22584
rect 24964 21962 24992 22578
rect 25332 21962 25360 24142
rect 24860 21956 24912 21962
rect 24860 21898 24912 21904
rect 24952 21956 25004 21962
rect 24952 21898 25004 21904
rect 25228 21956 25280 21962
rect 25228 21898 25280 21904
rect 25320 21956 25372 21962
rect 25320 21898 25372 21904
rect 24872 21690 24900 21898
rect 24860 21684 24912 21690
rect 24860 21626 24912 21632
rect 25240 20942 25268 21898
rect 25228 20936 25280 20942
rect 25228 20878 25280 20884
rect 24952 20868 25004 20874
rect 24952 20810 25004 20816
rect 25044 20868 25096 20874
rect 25044 20810 25096 20816
rect 24964 20398 24992 20810
rect 24952 20392 25004 20398
rect 24952 20334 25004 20340
rect 24860 20256 24912 20262
rect 25056 20210 25084 20810
rect 25320 20800 25372 20806
rect 25320 20742 25372 20748
rect 25332 20602 25360 20742
rect 25320 20596 25372 20602
rect 25320 20538 25372 20544
rect 25318 20496 25374 20505
rect 25424 20482 25452 26302
rect 25608 25702 25636 26318
rect 25596 25696 25648 25702
rect 25596 25638 25648 25644
rect 25792 25498 25820 30330
rect 25872 29096 25924 29102
rect 25872 29038 25924 29044
rect 25780 25492 25832 25498
rect 25780 25434 25832 25440
rect 25688 25152 25740 25158
rect 25688 25094 25740 25100
rect 25596 24880 25648 24886
rect 25596 24822 25648 24828
rect 25504 22636 25556 22642
rect 25504 22578 25556 22584
rect 25516 22234 25544 22578
rect 25504 22228 25556 22234
rect 25504 22170 25556 22176
rect 25504 21480 25556 21486
rect 25504 21422 25556 21428
rect 25374 20454 25452 20482
rect 25318 20431 25374 20440
rect 24912 20204 25084 20210
rect 24860 20198 25084 20204
rect 24872 20182 25084 20198
rect 24858 20088 24914 20097
rect 24858 20023 24860 20032
rect 24912 20023 24914 20032
rect 24860 19994 24912 20000
rect 24872 19514 24900 19994
rect 24860 19508 24912 19514
rect 24860 19450 24912 19456
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 24872 18154 24900 18226
rect 24768 18148 24820 18154
rect 24768 18090 24820 18096
rect 24860 18148 24912 18154
rect 24860 18090 24912 18096
rect 24584 18080 24636 18086
rect 24584 18022 24636 18028
rect 24676 18080 24728 18086
rect 24676 18022 24728 18028
rect 24596 17270 24624 18022
rect 24584 17264 24636 17270
rect 24584 17206 24636 17212
rect 24584 17128 24636 17134
rect 24584 17070 24636 17076
rect 24400 16652 24452 16658
rect 24400 16594 24452 16600
rect 24492 16584 24544 16590
rect 24492 16526 24544 16532
rect 24308 16108 24360 16114
rect 24308 16050 24360 16056
rect 24124 15700 24176 15706
rect 24124 15642 24176 15648
rect 24216 15700 24268 15706
rect 24216 15642 24268 15648
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 24032 15564 24084 15570
rect 24032 15506 24084 15512
rect 23952 15434 23980 15506
rect 23940 15428 23992 15434
rect 23940 15370 23992 15376
rect 24124 15360 24176 15366
rect 24044 15320 24124 15348
rect 24044 15162 24072 15320
rect 24124 15302 24176 15308
rect 24228 15162 24256 15642
rect 24400 15564 24452 15570
rect 24400 15506 24452 15512
rect 24032 15156 24084 15162
rect 24216 15156 24268 15162
rect 24032 15098 24084 15104
rect 24136 15116 24216 15144
rect 24044 14890 24072 15098
rect 24136 15026 24164 15116
rect 24268 15116 24348 15144
rect 24216 15098 24268 15104
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24032 14884 24084 14890
rect 24032 14826 24084 14832
rect 24124 14272 24176 14278
rect 24124 14214 24176 14220
rect 24136 14074 24164 14214
rect 24124 14068 24176 14074
rect 24124 14010 24176 14016
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 24124 13184 24176 13190
rect 24124 13126 24176 13132
rect 23572 12844 23624 12850
rect 23572 12786 23624 12792
rect 23664 12844 23716 12850
rect 23664 12786 23716 12792
rect 23584 12442 23612 12786
rect 23572 12436 23624 12442
rect 23572 12378 23624 12384
rect 23492 12294 23612 12322
rect 23480 12164 23532 12170
rect 23480 12106 23532 12112
rect 23492 11898 23520 12106
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23296 11620 23348 11626
rect 23296 11562 23348 11568
rect 23308 11150 23336 11562
rect 23296 11144 23348 11150
rect 23296 11086 23348 11092
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 23400 10810 23428 11086
rect 23388 10804 23440 10810
rect 23388 10746 23440 10752
rect 23584 10266 23612 12294
rect 23676 12238 23704 12786
rect 24136 12374 24164 13126
rect 23848 12368 23900 12374
rect 23848 12310 23900 12316
rect 24124 12368 24176 12374
rect 24124 12310 24176 12316
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23860 11898 23888 12310
rect 24030 12200 24086 12209
rect 24030 12135 24086 12144
rect 23848 11892 23900 11898
rect 23848 11834 23900 11840
rect 23664 11824 23716 11830
rect 23664 11766 23716 11772
rect 23572 10260 23624 10266
rect 23572 10202 23624 10208
rect 23216 10118 23428 10146
rect 23020 10056 23072 10062
rect 23020 9998 23072 10004
rect 23296 10056 23348 10062
rect 23296 9998 23348 10004
rect 23032 9586 23060 9998
rect 23204 9920 23256 9926
rect 23204 9862 23256 9868
rect 23216 9586 23244 9862
rect 23308 9722 23336 9998
rect 23296 9716 23348 9722
rect 23296 9658 23348 9664
rect 23020 9580 23072 9586
rect 23020 9522 23072 9528
rect 23204 9580 23256 9586
rect 23204 9522 23256 9528
rect 23112 9444 23164 9450
rect 23112 9386 23164 9392
rect 23124 8634 23152 9386
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 23112 8492 23164 8498
rect 23112 8434 23164 8440
rect 22928 8424 22980 8430
rect 22928 8366 22980 8372
rect 22928 8084 22980 8090
rect 22928 8026 22980 8032
rect 22940 7886 22968 8026
rect 22928 7880 22980 7886
rect 22928 7822 22980 7828
rect 23020 7880 23072 7886
rect 23020 7822 23072 7828
rect 22940 7546 22968 7822
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 23032 7478 23060 7822
rect 23020 7472 23072 7478
rect 23020 7414 23072 7420
rect 23124 7410 23152 8434
rect 23112 7404 23164 7410
rect 23112 7346 23164 7352
rect 22284 6792 22336 6798
rect 22284 6734 22336 6740
rect 22836 6792 22888 6798
rect 22836 6734 22888 6740
rect 22296 6322 22324 6734
rect 23124 6458 23152 7346
rect 23216 6866 23244 9522
rect 23400 8634 23428 10118
rect 23480 10056 23532 10062
rect 23480 9998 23532 10004
rect 23492 9654 23520 9998
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 23572 9580 23624 9586
rect 23572 9522 23624 9528
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 23388 8492 23440 8498
rect 23388 8434 23440 8440
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 23400 8294 23428 8434
rect 23296 8288 23348 8294
rect 23296 8230 23348 8236
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23308 8090 23336 8230
rect 23296 8084 23348 8090
rect 23296 8026 23348 8032
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 23400 7546 23428 7686
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23204 6860 23256 6866
rect 23204 6802 23256 6808
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 22284 6316 22336 6322
rect 22284 6258 22336 6264
rect 22296 5794 22324 6258
rect 22468 6112 22520 6118
rect 22468 6054 22520 6060
rect 22204 5778 22324 5794
rect 22480 5778 22508 6054
rect 22192 5772 22324 5778
rect 22244 5766 22324 5772
rect 22192 5714 22244 5720
rect 22296 5302 22324 5766
rect 22468 5772 22520 5778
rect 22468 5714 22520 5720
rect 23124 5642 23152 6394
rect 23400 6254 23428 6734
rect 23492 6730 23520 8434
rect 23480 6724 23532 6730
rect 23480 6666 23532 6672
rect 23388 6248 23440 6254
rect 23388 6190 23440 6196
rect 23492 5914 23520 6666
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 23400 5778 23520 5794
rect 23388 5772 23520 5778
rect 23440 5766 23520 5772
rect 23388 5714 23440 5720
rect 23112 5636 23164 5642
rect 23112 5578 23164 5584
rect 23204 5636 23256 5642
rect 23204 5578 23256 5584
rect 22284 5296 22336 5302
rect 22284 5238 22336 5244
rect 22296 4690 22324 5238
rect 22284 4684 22336 4690
rect 22284 4626 22336 4632
rect 22744 4548 22796 4554
rect 22744 4490 22796 4496
rect 22756 4282 22784 4490
rect 22744 4276 22796 4282
rect 22744 4218 22796 4224
rect 23216 4078 23244 5578
rect 23296 5160 23348 5166
rect 23296 5102 23348 5108
rect 23308 4146 23336 5102
rect 23492 4690 23520 5766
rect 23584 5234 23612 9522
rect 23676 7546 23704 11766
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 23952 11082 23980 11630
rect 23940 11076 23992 11082
rect 23940 11018 23992 11024
rect 23952 10742 23980 11018
rect 23848 10736 23900 10742
rect 23848 10678 23900 10684
rect 23940 10736 23992 10742
rect 23940 10678 23992 10684
rect 23860 10470 23888 10678
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 24044 9450 24072 12135
rect 24228 9654 24256 14962
rect 24320 9722 24348 15116
rect 24412 13870 24440 15506
rect 24504 14618 24532 16526
rect 24596 16454 24624 17070
rect 24584 16448 24636 16454
rect 24584 16390 24636 16396
rect 24596 15978 24624 16390
rect 24780 16182 24808 18090
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24872 17338 24900 17682
rect 24952 17604 25004 17610
rect 24952 17546 25004 17552
rect 24860 17332 24912 17338
rect 24860 17274 24912 17280
rect 24964 17134 24992 17546
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 25056 16980 25084 20182
rect 25228 19236 25280 19242
rect 25228 19178 25280 19184
rect 25136 18352 25188 18358
rect 25136 18294 25188 18300
rect 25148 17746 25176 18294
rect 25240 18290 25268 19178
rect 25332 18329 25360 20431
rect 25412 19372 25464 19378
rect 25412 19314 25464 19320
rect 25424 18970 25452 19314
rect 25412 18964 25464 18970
rect 25412 18906 25464 18912
rect 25424 18426 25452 18906
rect 25412 18420 25464 18426
rect 25412 18362 25464 18368
rect 25318 18320 25374 18329
rect 25228 18284 25280 18290
rect 25318 18255 25374 18264
rect 25228 18226 25280 18232
rect 25240 17814 25268 18226
rect 25320 18216 25372 18222
rect 25320 18158 25372 18164
rect 25228 17808 25280 17814
rect 25228 17750 25280 17756
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 25332 17542 25360 18158
rect 25424 18154 25452 18362
rect 25412 18148 25464 18154
rect 25412 18090 25464 18096
rect 25424 17882 25452 18090
rect 25412 17876 25464 17882
rect 25412 17818 25464 17824
rect 25136 17536 25188 17542
rect 25136 17478 25188 17484
rect 25320 17536 25372 17542
rect 25320 17478 25372 17484
rect 25148 17202 25176 17478
rect 25136 17196 25188 17202
rect 25136 17138 25188 17144
rect 24964 16952 25084 16980
rect 24676 16176 24728 16182
rect 24676 16118 24728 16124
rect 24768 16176 24820 16182
rect 24768 16118 24820 16124
rect 24584 15972 24636 15978
rect 24584 15914 24636 15920
rect 24688 15502 24716 16118
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24688 15026 24716 15438
rect 24768 15360 24820 15366
rect 24768 15302 24820 15308
rect 24676 15020 24728 15026
rect 24676 14962 24728 14968
rect 24492 14612 24544 14618
rect 24492 14554 24544 14560
rect 24780 14550 24808 15302
rect 24768 14544 24820 14550
rect 24768 14486 24820 14492
rect 24584 14476 24636 14482
rect 24584 14418 24636 14424
rect 24492 14272 24544 14278
rect 24492 14214 24544 14220
rect 24400 13864 24452 13870
rect 24400 13806 24452 13812
rect 24412 13530 24440 13806
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 24504 12434 24532 14214
rect 24596 13530 24624 14418
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 24688 13938 24716 14350
rect 24964 14278 24992 16952
rect 25320 16720 25372 16726
rect 25320 16662 25372 16668
rect 25332 16590 25360 16662
rect 25320 16584 25372 16590
rect 25320 16526 25372 16532
rect 25412 16516 25464 16522
rect 25412 16458 25464 16464
rect 25424 16250 25452 16458
rect 25412 16244 25464 16250
rect 25412 16186 25464 16192
rect 25320 16108 25372 16114
rect 25320 16050 25372 16056
rect 25332 15434 25360 16050
rect 25320 15428 25372 15434
rect 25320 15370 25372 15376
rect 25516 15366 25544 21422
rect 25608 19990 25636 24822
rect 25700 24410 25728 25094
rect 25792 24954 25820 25434
rect 25780 24948 25832 24954
rect 25780 24890 25832 24896
rect 25780 24812 25832 24818
rect 25780 24754 25832 24760
rect 25792 24426 25820 24754
rect 25884 24562 25912 29038
rect 25976 26518 26004 30534
rect 26056 30048 26108 30054
rect 26056 29990 26108 29996
rect 25964 26512 26016 26518
rect 25964 26454 26016 26460
rect 25976 26314 26004 26454
rect 26068 26330 26096 29990
rect 26160 27538 26188 32302
rect 26148 27532 26200 27538
rect 26148 27474 26200 27480
rect 26344 27112 26372 34138
rect 27264 33998 27292 35022
rect 28000 34746 28028 35226
rect 27988 34740 28040 34746
rect 27988 34682 28040 34688
rect 27804 34468 27856 34474
rect 27804 34410 27856 34416
rect 27620 34400 27672 34406
rect 27620 34342 27672 34348
rect 27632 33998 27660 34342
rect 26792 33992 26844 33998
rect 26792 33934 26844 33940
rect 27252 33992 27304 33998
rect 27252 33934 27304 33940
rect 27620 33992 27672 33998
rect 27620 33934 27672 33940
rect 26424 33924 26476 33930
rect 26424 33866 26476 33872
rect 26436 32858 26464 33866
rect 26804 33454 26832 33934
rect 27528 33584 27580 33590
rect 27528 33526 27580 33532
rect 26792 33448 26844 33454
rect 26792 33390 26844 33396
rect 26608 33312 26660 33318
rect 26608 33254 26660 33260
rect 26436 32830 26556 32858
rect 26620 32842 26648 33254
rect 26528 31346 26556 32830
rect 26608 32836 26660 32842
rect 26608 32778 26660 32784
rect 26700 32224 26752 32230
rect 26700 32166 26752 32172
rect 26712 31362 26740 32166
rect 26804 31822 26832 33390
rect 26976 32768 27028 32774
rect 26976 32710 27028 32716
rect 26792 31816 26844 31822
rect 26792 31758 26844 31764
rect 26988 31754 27016 32710
rect 26896 31726 27016 31754
rect 27066 31784 27122 31793
rect 27540 31754 27568 33526
rect 27712 33448 27764 33454
rect 27816 33436 27844 34410
rect 27764 33408 27844 33436
rect 27712 33390 27764 33396
rect 27620 32428 27672 32434
rect 27620 32370 27672 32376
rect 26712 31346 26832 31362
rect 26516 31340 26568 31346
rect 26712 31340 26844 31346
rect 26712 31334 26792 31340
rect 26516 31282 26568 31288
rect 26792 31282 26844 31288
rect 26804 31142 26832 31282
rect 26792 31136 26844 31142
rect 26792 31078 26844 31084
rect 26424 29504 26476 29510
rect 26424 29446 26476 29452
rect 26436 29073 26464 29446
rect 26422 29064 26478 29073
rect 26422 28999 26478 29008
rect 26424 28076 26476 28082
rect 26424 28018 26476 28024
rect 26436 27878 26464 28018
rect 26424 27872 26476 27878
rect 26424 27814 26476 27820
rect 26516 27872 26568 27878
rect 26516 27814 26568 27820
rect 26436 27470 26464 27814
rect 26424 27464 26476 27470
rect 26424 27406 26476 27412
rect 26528 27402 26556 27814
rect 26516 27396 26568 27402
rect 26516 27338 26568 27344
rect 26344 27084 26464 27112
rect 26332 26988 26384 26994
rect 26332 26930 26384 26936
rect 26344 26790 26372 26930
rect 26332 26784 26384 26790
rect 26332 26726 26384 26732
rect 26240 26580 26292 26586
rect 26240 26522 26292 26528
rect 26252 26382 26280 26522
rect 26240 26376 26292 26382
rect 26238 26344 26240 26353
rect 26292 26344 26294 26353
rect 25964 26308 26016 26314
rect 26068 26302 26188 26330
rect 25964 26250 26016 26256
rect 26056 26240 26108 26246
rect 26056 26182 26108 26188
rect 26068 24682 26096 26182
rect 26056 24676 26108 24682
rect 26056 24618 26108 24624
rect 26160 24614 26188 26302
rect 26238 26279 26294 26288
rect 26344 26217 26372 26726
rect 26330 26208 26386 26217
rect 26330 26143 26386 26152
rect 26240 25152 26292 25158
rect 26240 25094 26292 25100
rect 26252 24886 26280 25094
rect 26240 24880 26292 24886
rect 26240 24822 26292 24828
rect 26252 24614 26280 24822
rect 26148 24608 26200 24614
rect 25884 24534 26096 24562
rect 26148 24550 26200 24556
rect 26240 24608 26292 24614
rect 26240 24550 26292 24556
rect 25688 24404 25740 24410
rect 25792 24398 25912 24426
rect 25688 24346 25740 24352
rect 25700 24274 25728 24346
rect 25688 24268 25740 24274
rect 25688 24210 25740 24216
rect 25780 24064 25832 24070
rect 25884 24041 25912 24398
rect 25964 24200 26016 24206
rect 25964 24142 26016 24148
rect 25780 24006 25832 24012
rect 25870 24032 25926 24041
rect 25792 23322 25820 24006
rect 25870 23967 25926 23976
rect 25780 23316 25832 23322
rect 25780 23258 25832 23264
rect 25780 22092 25832 22098
rect 25780 22034 25832 22040
rect 25792 21434 25820 22034
rect 25884 21570 25912 23967
rect 25976 22778 26004 24142
rect 25964 22772 26016 22778
rect 25964 22714 26016 22720
rect 25976 22098 26004 22714
rect 25964 22092 26016 22098
rect 25964 22034 26016 22040
rect 26068 21690 26096 24534
rect 26160 24274 26188 24550
rect 26252 24342 26280 24550
rect 26436 24449 26464 27084
rect 26528 26382 26556 27338
rect 26700 27124 26752 27130
rect 26700 27066 26752 27072
rect 26606 26888 26662 26897
rect 26606 26823 26662 26832
rect 26620 26790 26648 26823
rect 26608 26784 26660 26790
rect 26608 26726 26660 26732
rect 26712 26450 26740 27066
rect 26700 26444 26752 26450
rect 26700 26386 26752 26392
rect 26516 26376 26568 26382
rect 26516 26318 26568 26324
rect 26528 26042 26556 26318
rect 26516 26036 26568 26042
rect 26516 25978 26568 25984
rect 26422 24440 26478 24449
rect 26422 24375 26478 24384
rect 26698 24440 26754 24449
rect 26698 24375 26754 24384
rect 26240 24336 26292 24342
rect 26240 24278 26292 24284
rect 26514 24304 26570 24313
rect 26148 24268 26200 24274
rect 26514 24239 26570 24248
rect 26148 24210 26200 24216
rect 26160 23905 26188 24210
rect 26528 24206 26556 24239
rect 26240 24200 26292 24206
rect 26516 24200 26568 24206
rect 26240 24142 26292 24148
rect 26436 24148 26516 24154
rect 26436 24142 26568 24148
rect 26252 24070 26280 24142
rect 26436 24126 26556 24142
rect 26240 24064 26292 24070
rect 26240 24006 26292 24012
rect 26146 23896 26202 23905
rect 26146 23831 26202 23840
rect 26148 23520 26200 23526
rect 26148 23462 26200 23468
rect 26160 22098 26188 23462
rect 26252 22982 26280 24006
rect 26330 23760 26386 23769
rect 26330 23695 26332 23704
rect 26384 23695 26386 23704
rect 26332 23666 26384 23672
rect 26240 22976 26292 22982
rect 26240 22918 26292 22924
rect 26344 22642 26372 23666
rect 26436 23322 26464 24126
rect 26516 23860 26568 23866
rect 26516 23802 26568 23808
rect 26528 23322 26556 23802
rect 26608 23656 26660 23662
rect 26608 23598 26660 23604
rect 26424 23316 26476 23322
rect 26424 23258 26476 23264
rect 26516 23316 26568 23322
rect 26516 23258 26568 23264
rect 26332 22636 26384 22642
rect 26332 22578 26384 22584
rect 26148 22092 26200 22098
rect 26436 22094 26464 23258
rect 26528 22234 26556 23258
rect 26620 22778 26648 23598
rect 26608 22772 26660 22778
rect 26608 22714 26660 22720
rect 26516 22228 26568 22234
rect 26516 22170 26568 22176
rect 26148 22034 26200 22040
rect 26344 22066 26464 22094
rect 26528 22094 26556 22170
rect 26528 22066 26648 22094
rect 26056 21684 26108 21690
rect 26056 21626 26108 21632
rect 25884 21542 26004 21570
rect 25792 21406 25912 21434
rect 25780 21344 25832 21350
rect 25700 21304 25780 21332
rect 25700 20874 25728 21304
rect 25780 21286 25832 21292
rect 25884 21146 25912 21406
rect 25872 21140 25924 21146
rect 25792 21100 25872 21128
rect 25688 20868 25740 20874
rect 25688 20810 25740 20816
rect 25596 19984 25648 19990
rect 25596 19926 25648 19932
rect 25608 16998 25636 19926
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 25700 18426 25728 19110
rect 25688 18420 25740 18426
rect 25688 18362 25740 18368
rect 25686 18320 25742 18329
rect 25686 18255 25742 18264
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25608 16658 25636 16934
rect 25596 16652 25648 16658
rect 25596 16594 25648 16600
rect 25700 16266 25728 18255
rect 25608 16238 25728 16266
rect 25504 15360 25556 15366
rect 25504 15302 25556 15308
rect 25228 15020 25280 15026
rect 25228 14962 25280 14968
rect 25240 14618 25268 14962
rect 25228 14612 25280 14618
rect 25228 14554 25280 14560
rect 24952 14272 25004 14278
rect 24872 14220 24952 14226
rect 24872 14214 25004 14220
rect 24872 14198 24992 14214
rect 24872 14074 24900 14198
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24872 13938 24900 14010
rect 25412 14000 25464 14006
rect 25412 13942 25464 13948
rect 24676 13932 24728 13938
rect 24676 13874 24728 13880
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 24768 13864 24820 13870
rect 24768 13806 24820 13812
rect 24584 13524 24636 13530
rect 24584 13466 24636 13472
rect 24780 12986 24808 13806
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24676 12912 24728 12918
rect 24676 12854 24728 12860
rect 24412 12406 24532 12434
rect 24412 11626 24440 12406
rect 24492 12368 24544 12374
rect 24492 12310 24544 12316
rect 24400 11620 24452 11626
rect 24400 11562 24452 11568
rect 24400 10056 24452 10062
rect 24400 9998 24452 10004
rect 24308 9716 24360 9722
rect 24308 9658 24360 9664
rect 24216 9648 24268 9654
rect 24216 9590 24268 9596
rect 24412 9586 24440 9998
rect 24124 9580 24176 9586
rect 24124 9522 24176 9528
rect 24400 9580 24452 9586
rect 24400 9522 24452 9528
rect 24032 9444 24084 9450
rect 24032 9386 24084 9392
rect 24136 9382 24164 9522
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 24124 9376 24176 9382
rect 24124 9318 24176 9324
rect 23768 8362 23796 9318
rect 23860 8974 23888 9318
rect 24412 9110 24440 9522
rect 24400 9104 24452 9110
rect 24400 9046 24452 9052
rect 23848 8968 23900 8974
rect 23848 8910 23900 8916
rect 24504 8838 24532 12310
rect 24688 11762 24716 12854
rect 25228 12776 25280 12782
rect 25228 12718 25280 12724
rect 24952 12708 25004 12714
rect 24952 12650 25004 12656
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 24872 12102 24900 12582
rect 24964 12306 24992 12650
rect 24952 12300 25004 12306
rect 24952 12242 25004 12248
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 25044 11892 25096 11898
rect 25044 11834 25096 11840
rect 25056 11762 25084 11834
rect 24676 11756 24728 11762
rect 24676 11698 24728 11704
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 24952 11076 25004 11082
rect 24952 11018 25004 11024
rect 24964 10810 24992 11018
rect 24952 10804 25004 10810
rect 24952 10746 25004 10752
rect 24768 10056 24820 10062
rect 24768 9998 24820 10004
rect 24780 9674 24808 9998
rect 24780 9646 25176 9674
rect 25240 9654 25268 12718
rect 25148 9586 25176 9646
rect 25228 9648 25280 9654
rect 25228 9590 25280 9596
rect 25136 9580 25188 9586
rect 25136 9522 25188 9528
rect 25320 9580 25372 9586
rect 25320 9522 25372 9528
rect 24584 9104 24636 9110
rect 24584 9046 24636 9052
rect 24492 8832 24544 8838
rect 24492 8774 24544 8780
rect 23756 8356 23808 8362
rect 23756 8298 23808 8304
rect 23756 7880 23808 7886
rect 23756 7822 23808 7828
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 23664 7540 23716 7546
rect 23664 7482 23716 7488
rect 23664 6996 23716 7002
rect 23664 6938 23716 6944
rect 23676 6798 23704 6938
rect 23664 6792 23716 6798
rect 23664 6734 23716 6740
rect 23768 6458 23796 7822
rect 23860 7546 23888 7822
rect 23848 7540 23900 7546
rect 23848 7482 23900 7488
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 24320 6780 24348 7346
rect 24400 6792 24452 6798
rect 24320 6752 24400 6780
rect 24400 6734 24452 6740
rect 23756 6452 23808 6458
rect 23756 6394 23808 6400
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23676 6118 23704 6258
rect 23768 6236 23796 6394
rect 23848 6248 23900 6254
rect 23768 6208 23848 6236
rect 23848 6190 23900 6196
rect 23664 6112 23716 6118
rect 23664 6054 23716 6060
rect 23756 6112 23808 6118
rect 23756 6054 23808 6060
rect 23768 5710 23796 6054
rect 23756 5704 23808 5710
rect 23756 5646 23808 5652
rect 23572 5228 23624 5234
rect 23572 5170 23624 5176
rect 23480 4684 23532 4690
rect 23480 4626 23532 4632
rect 23584 4486 23612 5170
rect 23860 5166 23888 6190
rect 24412 5914 24440 6734
rect 24504 6662 24532 7346
rect 24596 6730 24624 9046
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 24780 7410 24808 7482
rect 24768 7404 24820 7410
rect 24768 7346 24820 7352
rect 24780 6798 24808 7346
rect 24768 6792 24820 6798
rect 24768 6734 24820 6740
rect 24584 6724 24636 6730
rect 24584 6666 24636 6672
rect 24492 6656 24544 6662
rect 24492 6598 24544 6604
rect 24504 6322 24532 6598
rect 24596 6458 24624 6666
rect 24584 6452 24636 6458
rect 24584 6394 24636 6400
rect 24596 6322 24624 6394
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 24400 5908 24452 5914
rect 24400 5850 24452 5856
rect 23940 5772 23992 5778
rect 23940 5714 23992 5720
rect 23952 5166 23980 5714
rect 24032 5364 24084 5370
rect 24032 5306 24084 5312
rect 24044 5234 24072 5306
rect 24032 5228 24084 5234
rect 24032 5170 24084 5176
rect 23848 5160 23900 5166
rect 23848 5102 23900 5108
rect 23940 5160 23992 5166
rect 23940 5102 23992 5108
rect 24412 4554 24440 5850
rect 24780 5370 24808 6734
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 24872 5302 24900 8978
rect 25148 8294 25176 9522
rect 25332 9178 25360 9522
rect 25424 9450 25452 13942
rect 25504 13252 25556 13258
rect 25504 13194 25556 13200
rect 25516 12986 25544 13194
rect 25504 12980 25556 12986
rect 25504 12922 25556 12928
rect 25608 12646 25636 16238
rect 25792 15978 25820 21100
rect 25872 21082 25924 21088
rect 25976 19786 26004 21542
rect 26068 21486 26096 21626
rect 26056 21480 26108 21486
rect 26056 21422 26108 21428
rect 26056 20800 26108 20806
rect 26056 20742 26108 20748
rect 26068 20602 26096 20742
rect 26056 20596 26108 20602
rect 26056 20538 26108 20544
rect 26068 20398 26096 20538
rect 26056 20392 26108 20398
rect 26056 20334 26108 20340
rect 26148 19848 26200 19854
rect 26148 19790 26200 19796
rect 25964 19780 26016 19786
rect 25964 19722 26016 19728
rect 25976 19417 26004 19722
rect 25962 19408 26018 19417
rect 25962 19343 26018 19352
rect 25964 19304 26016 19310
rect 25964 19246 26016 19252
rect 25872 19168 25924 19174
rect 25872 19110 25924 19116
rect 25884 18714 25912 19110
rect 25976 18834 26004 19246
rect 25964 18828 26016 18834
rect 25964 18770 26016 18776
rect 25884 18686 26004 18714
rect 25976 18630 26004 18686
rect 26056 18692 26108 18698
rect 26056 18634 26108 18640
rect 25964 18624 26016 18630
rect 25964 18566 26016 18572
rect 25976 18204 26004 18566
rect 26068 18358 26096 18634
rect 26056 18352 26108 18358
rect 26056 18294 26108 18300
rect 25976 18176 26096 18204
rect 25872 18148 25924 18154
rect 25872 18090 25924 18096
rect 25884 17882 25912 18090
rect 25962 17912 26018 17921
rect 25872 17876 25924 17882
rect 25962 17847 25964 17856
rect 25872 17818 25924 17824
rect 26016 17847 26018 17856
rect 25964 17818 26016 17824
rect 26068 17762 26096 18176
rect 26160 17882 26188 19790
rect 26240 19508 26292 19514
rect 26240 19450 26292 19456
rect 26252 18970 26280 19450
rect 26344 19174 26372 22066
rect 26620 22030 26648 22066
rect 26608 22024 26660 22030
rect 26608 21966 26660 21972
rect 26422 21448 26478 21457
rect 26422 21383 26478 21392
rect 26436 20602 26464 21383
rect 26424 20596 26476 20602
rect 26424 20538 26476 20544
rect 26436 20398 26464 20538
rect 26608 20460 26660 20466
rect 26608 20402 26660 20408
rect 26424 20392 26476 20398
rect 26424 20334 26476 20340
rect 26620 20330 26648 20402
rect 26608 20324 26660 20330
rect 26608 20266 26660 20272
rect 26620 20233 26648 20266
rect 26606 20224 26662 20233
rect 26606 20159 26662 20168
rect 26712 19922 26740 24375
rect 26804 24041 26832 31078
rect 26896 28218 26924 31726
rect 27066 31719 27068 31728
rect 27120 31719 27122 31728
rect 27436 31748 27488 31754
rect 27068 31690 27120 31696
rect 27436 31690 27488 31696
rect 27528 31748 27580 31754
rect 27528 31690 27580 31696
rect 27448 31414 27476 31690
rect 27436 31408 27488 31414
rect 27066 31376 27122 31385
rect 27436 31350 27488 31356
rect 27066 31311 27122 31320
rect 27080 31142 27108 31311
rect 27068 31136 27120 31142
rect 27068 31078 27120 31084
rect 27448 30682 27476 31350
rect 27540 30938 27568 31690
rect 27632 31482 27660 32370
rect 27620 31476 27672 31482
rect 27620 31418 27672 31424
rect 27528 30932 27580 30938
rect 27528 30874 27580 30880
rect 27264 30654 27476 30682
rect 27068 30252 27120 30258
rect 27068 30194 27120 30200
rect 27080 29850 27108 30194
rect 27160 30184 27212 30190
rect 27160 30126 27212 30132
rect 27172 29850 27200 30126
rect 27068 29844 27120 29850
rect 27068 29786 27120 29792
rect 27160 29844 27212 29850
rect 27160 29786 27212 29792
rect 27264 29714 27292 30654
rect 27540 30546 27568 30874
rect 27632 30598 27660 31418
rect 27448 30518 27568 30546
rect 27620 30592 27672 30598
rect 27620 30534 27672 30540
rect 27344 30252 27396 30258
rect 27344 30194 27396 30200
rect 27356 29850 27384 30194
rect 27344 29844 27396 29850
rect 27344 29786 27396 29792
rect 27252 29708 27304 29714
rect 27172 29668 27252 29696
rect 26976 29572 27028 29578
rect 26976 29514 27028 29520
rect 26988 29306 27016 29514
rect 26976 29300 27028 29306
rect 26976 29242 27028 29248
rect 27172 28626 27200 29668
rect 27252 29650 27304 29656
rect 27356 29306 27384 29786
rect 27344 29300 27396 29306
rect 27344 29242 27396 29248
rect 27448 29170 27476 30518
rect 27526 30424 27582 30433
rect 27526 30359 27582 30368
rect 27540 30054 27568 30359
rect 27528 30048 27580 30054
rect 27528 29990 27580 29996
rect 27528 29504 27580 29510
rect 27528 29446 27580 29452
rect 27436 29164 27488 29170
rect 27436 29106 27488 29112
rect 27540 29102 27568 29446
rect 27528 29096 27580 29102
rect 27528 29038 27580 29044
rect 27160 28620 27212 28626
rect 27160 28562 27212 28568
rect 27620 28484 27672 28490
rect 27620 28426 27672 28432
rect 27632 28218 27660 28426
rect 26884 28212 26936 28218
rect 26884 28154 26936 28160
rect 27068 28212 27120 28218
rect 27068 28154 27120 28160
rect 27620 28212 27672 28218
rect 27620 28154 27672 28160
rect 26976 27328 27028 27334
rect 26976 27270 27028 27276
rect 26988 27130 27016 27270
rect 26976 27124 27028 27130
rect 26976 27066 27028 27072
rect 26988 26382 27016 27066
rect 26976 26376 27028 26382
rect 26976 26318 27028 26324
rect 26976 25220 27028 25226
rect 26976 25162 27028 25168
rect 26988 24954 27016 25162
rect 26976 24948 27028 24954
rect 26976 24890 27028 24896
rect 26884 24744 26936 24750
rect 26884 24686 26936 24692
rect 26976 24744 27028 24750
rect 26976 24686 27028 24692
rect 26896 24410 26924 24686
rect 26884 24404 26936 24410
rect 26884 24346 26936 24352
rect 26988 24177 27016 24686
rect 27080 24614 27108 28154
rect 27436 27872 27488 27878
rect 27436 27814 27488 27820
rect 27158 27568 27214 27577
rect 27158 27503 27214 27512
rect 27172 27470 27200 27503
rect 27448 27470 27476 27814
rect 27528 27532 27580 27538
rect 27528 27474 27580 27480
rect 27160 27464 27212 27470
rect 27160 27406 27212 27412
rect 27436 27464 27488 27470
rect 27436 27406 27488 27412
rect 27344 26988 27396 26994
rect 27344 26930 27396 26936
rect 27356 26586 27384 26930
rect 27344 26580 27396 26586
rect 27344 26522 27396 26528
rect 27436 26512 27488 26518
rect 27436 26454 27488 26460
rect 27252 25900 27304 25906
rect 27252 25842 27304 25848
rect 27264 25498 27292 25842
rect 27252 25492 27304 25498
rect 27252 25434 27304 25440
rect 27264 24818 27292 25434
rect 27344 25152 27396 25158
rect 27344 25094 27396 25100
rect 27356 24954 27384 25094
rect 27344 24948 27396 24954
rect 27344 24890 27396 24896
rect 27252 24812 27304 24818
rect 27252 24754 27304 24760
rect 27068 24608 27120 24614
rect 27068 24550 27120 24556
rect 27080 24206 27108 24550
rect 27252 24404 27304 24410
rect 27252 24346 27304 24352
rect 27264 24206 27292 24346
rect 27356 24206 27384 24890
rect 27068 24200 27120 24206
rect 26974 24168 27030 24177
rect 27068 24142 27120 24148
rect 27252 24200 27304 24206
rect 27252 24142 27304 24148
rect 27344 24200 27396 24206
rect 27344 24142 27396 24148
rect 26974 24103 27030 24112
rect 27160 24132 27212 24138
rect 27160 24074 27212 24080
rect 26790 24032 26846 24041
rect 26790 23967 26846 23976
rect 27172 23526 27200 24074
rect 27252 23724 27304 23730
rect 27252 23666 27304 23672
rect 27160 23520 27212 23526
rect 27160 23462 27212 23468
rect 27172 23118 27200 23462
rect 27264 23322 27292 23666
rect 27252 23316 27304 23322
rect 27252 23258 27304 23264
rect 27160 23112 27212 23118
rect 27448 23100 27476 26454
rect 27540 24698 27568 27474
rect 27620 27328 27672 27334
rect 27620 27270 27672 27276
rect 27632 26450 27660 27270
rect 27620 26444 27672 26450
rect 27620 26386 27672 26392
rect 27618 25664 27674 25673
rect 27618 25599 27674 25608
rect 27632 24886 27660 25599
rect 27620 24880 27672 24886
rect 27620 24822 27672 24828
rect 27620 24744 27672 24750
rect 27540 24692 27620 24698
rect 27540 24686 27672 24692
rect 27540 24670 27660 24686
rect 27540 23254 27568 24670
rect 27620 24200 27672 24206
rect 27620 24142 27672 24148
rect 27632 23497 27660 24142
rect 27618 23488 27674 23497
rect 27618 23423 27674 23432
rect 27724 23322 27752 33390
rect 27804 32496 27856 32502
rect 27804 32438 27856 32444
rect 27816 31686 27844 32438
rect 28000 32314 28028 34682
rect 28080 34604 28132 34610
rect 28080 34546 28132 34552
rect 28092 34202 28120 34546
rect 28080 34196 28132 34202
rect 28080 34138 28132 34144
rect 28460 33522 28488 35226
rect 28632 34196 28684 34202
rect 28632 34138 28684 34144
rect 28644 33590 28672 34138
rect 34060 33992 34112 33998
rect 34060 33934 34112 33940
rect 29184 33856 29236 33862
rect 29184 33798 29236 33804
rect 32864 33856 32916 33862
rect 32864 33798 32916 33804
rect 28632 33584 28684 33590
rect 28632 33526 28684 33532
rect 28264 33516 28316 33522
rect 28264 33458 28316 33464
rect 28448 33516 28500 33522
rect 28448 33458 28500 33464
rect 28724 33516 28776 33522
rect 28724 33458 28776 33464
rect 28172 32836 28224 32842
rect 28172 32778 28224 32784
rect 28184 32434 28212 32778
rect 28276 32570 28304 33458
rect 28356 33108 28408 33114
rect 28356 33050 28408 33056
rect 28368 32570 28396 33050
rect 28736 32910 28764 33458
rect 29196 33318 29224 33798
rect 29276 33516 29328 33522
rect 29276 33458 29328 33464
rect 29828 33516 29880 33522
rect 29828 33458 29880 33464
rect 29184 33312 29236 33318
rect 29184 33254 29236 33260
rect 28724 32904 28776 32910
rect 28724 32846 28776 32852
rect 28632 32768 28684 32774
rect 28632 32710 28684 32716
rect 28264 32564 28316 32570
rect 28264 32506 28316 32512
rect 28356 32564 28408 32570
rect 28356 32506 28408 32512
rect 28644 32502 28672 32710
rect 28632 32496 28684 32502
rect 28632 32438 28684 32444
rect 28172 32428 28224 32434
rect 28172 32370 28224 32376
rect 28264 32428 28316 32434
rect 28264 32370 28316 32376
rect 28540 32428 28592 32434
rect 28540 32370 28592 32376
rect 28000 32286 28212 32314
rect 27988 32020 28040 32026
rect 27988 31962 28040 31968
rect 27896 31952 27948 31958
rect 27896 31894 27948 31900
rect 27908 31793 27936 31894
rect 27894 31784 27950 31793
rect 27894 31719 27950 31728
rect 27804 31680 27856 31686
rect 27804 31622 27856 31628
rect 28000 30666 28028 31962
rect 28184 31754 28212 32286
rect 28172 31748 28224 31754
rect 28172 31690 28224 31696
rect 28276 31482 28304 32370
rect 28448 32360 28500 32366
rect 28448 32302 28500 32308
rect 28264 31476 28316 31482
rect 28264 31418 28316 31424
rect 28356 31340 28408 31346
rect 28356 31282 28408 31288
rect 28368 30938 28396 31282
rect 28356 30932 28408 30938
rect 28356 30874 28408 30880
rect 27988 30660 28040 30666
rect 27988 30602 28040 30608
rect 27896 30592 27948 30598
rect 27896 30534 27948 30540
rect 27802 24440 27858 24449
rect 27802 24375 27858 24384
rect 27816 24206 27844 24375
rect 27804 24200 27856 24206
rect 27804 24142 27856 24148
rect 27804 24064 27856 24070
rect 27802 24032 27804 24041
rect 27856 24032 27858 24041
rect 27802 23967 27858 23976
rect 27712 23316 27764 23322
rect 27712 23258 27764 23264
rect 27528 23248 27580 23254
rect 27528 23190 27580 23196
rect 27448 23072 27568 23100
rect 27160 23054 27212 23060
rect 27252 22772 27304 22778
rect 27252 22714 27304 22720
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 27068 22024 27120 22030
rect 27068 21966 27120 21972
rect 26884 21412 26936 21418
rect 26884 21354 26936 21360
rect 26790 20360 26846 20369
rect 26790 20295 26792 20304
rect 26844 20295 26846 20304
rect 26792 20266 26844 20272
rect 26700 19916 26752 19922
rect 26700 19858 26752 19864
rect 26712 19718 26740 19858
rect 26700 19712 26752 19718
rect 26700 19654 26752 19660
rect 26424 19440 26476 19446
rect 26476 19417 26556 19428
rect 26476 19408 26570 19417
rect 26476 19400 26514 19408
rect 26424 19382 26476 19388
rect 26792 19372 26844 19378
rect 26514 19343 26570 19352
rect 26608 19346 26660 19352
rect 26332 19168 26384 19174
rect 26332 19110 26384 19116
rect 26424 19168 26476 19174
rect 26424 19110 26476 19116
rect 26240 18964 26292 18970
rect 26240 18906 26292 18912
rect 26332 18964 26384 18970
rect 26332 18906 26384 18912
rect 26252 18698 26280 18906
rect 26240 18692 26292 18698
rect 26240 18634 26292 18640
rect 26344 18426 26372 18906
rect 26436 18834 26464 19110
rect 26424 18828 26476 18834
rect 26424 18770 26476 18776
rect 26528 18714 26556 19343
rect 26792 19314 26844 19320
rect 26608 19288 26660 19294
rect 26436 18686 26556 18714
rect 26332 18420 26384 18426
rect 26332 18362 26384 18368
rect 26148 17876 26200 17882
rect 26148 17818 26200 17824
rect 25976 17734 26096 17762
rect 26344 17746 26372 18362
rect 26332 17740 26384 17746
rect 25872 16448 25924 16454
rect 25872 16390 25924 16396
rect 25884 16182 25912 16390
rect 25872 16176 25924 16182
rect 25872 16118 25924 16124
rect 25780 15972 25832 15978
rect 25780 15914 25832 15920
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 25700 13734 25728 14214
rect 25688 13728 25740 13734
rect 25688 13670 25740 13676
rect 25596 12640 25648 12646
rect 25596 12582 25648 12588
rect 25504 11552 25556 11558
rect 25504 11494 25556 11500
rect 25516 11014 25544 11494
rect 25504 11008 25556 11014
rect 25504 10950 25556 10956
rect 25516 10606 25544 10950
rect 25608 10674 25636 12582
rect 25792 12442 25820 15914
rect 25780 12436 25832 12442
rect 25780 12378 25832 12384
rect 25792 12238 25820 12378
rect 25780 12232 25832 12238
rect 25780 12174 25832 12180
rect 25872 12096 25924 12102
rect 25976 12084 26004 17734
rect 26332 17682 26384 17688
rect 26436 17678 26464 18686
rect 26516 18624 26568 18630
rect 26516 18566 26568 18572
rect 26424 17672 26476 17678
rect 26424 17614 26476 17620
rect 26332 17196 26384 17202
rect 26332 17138 26384 17144
rect 26148 16720 26200 16726
rect 26148 16662 26200 16668
rect 26056 16448 26108 16454
rect 26056 16390 26108 16396
rect 26068 15434 26096 16390
rect 26056 15428 26108 15434
rect 26056 15370 26108 15376
rect 26160 14618 26188 16662
rect 26344 16114 26372 17138
rect 26528 16590 26556 18566
rect 26620 18358 26648 19288
rect 26804 18834 26832 19314
rect 26792 18828 26844 18834
rect 26792 18770 26844 18776
rect 26700 18760 26752 18766
rect 26700 18702 26752 18708
rect 26608 18352 26660 18358
rect 26608 18294 26660 18300
rect 26712 18154 26740 18702
rect 26792 18624 26844 18630
rect 26792 18566 26844 18572
rect 26700 18148 26752 18154
rect 26700 18090 26752 18096
rect 26608 17264 26660 17270
rect 26608 17206 26660 17212
rect 26620 16658 26648 17206
rect 26608 16652 26660 16658
rect 26608 16594 26660 16600
rect 26516 16584 26568 16590
rect 26516 16526 26568 16532
rect 26424 16448 26476 16454
rect 26424 16390 26476 16396
rect 26332 16108 26384 16114
rect 26332 16050 26384 16056
rect 26436 16046 26464 16390
rect 26424 16040 26476 16046
rect 26424 15982 26476 15988
rect 26436 15706 26464 15982
rect 26424 15700 26476 15706
rect 26424 15642 26476 15648
rect 26516 15632 26568 15638
rect 26516 15574 26568 15580
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26148 14612 26200 14618
rect 26068 14572 26148 14600
rect 26068 13938 26096 14572
rect 26148 14554 26200 14560
rect 26148 14476 26200 14482
rect 26148 14418 26200 14424
rect 26160 14278 26188 14418
rect 26252 14414 26280 15098
rect 26528 14822 26556 15574
rect 26332 14816 26384 14822
rect 26332 14758 26384 14764
rect 26516 14816 26568 14822
rect 26516 14758 26568 14764
rect 26240 14408 26292 14414
rect 26240 14350 26292 14356
rect 26148 14272 26200 14278
rect 26148 14214 26200 14220
rect 26160 14006 26188 14214
rect 26148 14000 26200 14006
rect 26148 13942 26200 13948
rect 26056 13932 26108 13938
rect 26056 13874 26108 13880
rect 26160 12782 26188 13942
rect 26344 13530 26372 14758
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 26332 13524 26384 13530
rect 26332 13466 26384 13472
rect 26436 13326 26464 14010
rect 26516 13796 26568 13802
rect 26516 13738 26568 13744
rect 26424 13320 26476 13326
rect 26424 13262 26476 13268
rect 26332 13184 26384 13190
rect 26332 13126 26384 13132
rect 26344 12986 26372 13126
rect 26332 12980 26384 12986
rect 26332 12922 26384 12928
rect 26528 12850 26556 13738
rect 26620 13274 26648 16594
rect 26804 15570 26832 18566
rect 26896 17066 26924 21354
rect 27080 21010 27108 21966
rect 27068 21004 27120 21010
rect 27068 20946 27120 20952
rect 26976 20868 27028 20874
rect 26976 20810 27028 20816
rect 26988 20602 27016 20810
rect 26976 20596 27028 20602
rect 26976 20538 27028 20544
rect 26976 19712 27028 19718
rect 26976 19654 27028 19660
rect 26884 17060 26936 17066
rect 26884 17002 26936 17008
rect 26896 16182 26924 17002
rect 26884 16176 26936 16182
rect 26884 16118 26936 16124
rect 26896 15706 26924 16118
rect 26884 15700 26936 15706
rect 26884 15642 26936 15648
rect 26792 15564 26844 15570
rect 26792 15506 26844 15512
rect 26988 15450 27016 19654
rect 27068 18352 27120 18358
rect 27068 18294 27120 18300
rect 27080 17746 27108 18294
rect 27068 17740 27120 17746
rect 27068 17682 27120 17688
rect 27068 17332 27120 17338
rect 27068 17274 27120 17280
rect 27080 16794 27108 17274
rect 27068 16788 27120 16794
rect 27068 16730 27120 16736
rect 27080 16697 27108 16730
rect 27066 16688 27122 16697
rect 27066 16623 27122 16632
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 26804 15422 27016 15450
rect 26620 13246 26740 13274
rect 26608 13184 26660 13190
rect 26608 13126 26660 13132
rect 26516 12844 26568 12850
rect 26516 12786 26568 12792
rect 26148 12776 26200 12782
rect 26148 12718 26200 12724
rect 26160 12481 26188 12718
rect 26424 12708 26476 12714
rect 26424 12650 26476 12656
rect 26146 12472 26202 12481
rect 26202 12416 26280 12434
rect 26146 12407 26280 12416
rect 26160 12406 26280 12407
rect 26252 12374 26280 12406
rect 26240 12368 26292 12374
rect 26240 12310 26292 12316
rect 26332 12232 26384 12238
rect 26332 12174 26384 12180
rect 25924 12056 26004 12084
rect 25872 12038 25924 12044
rect 25884 11898 25912 12038
rect 25872 11892 25924 11898
rect 25872 11834 25924 11840
rect 26148 11824 26200 11830
rect 26148 11766 26200 11772
rect 26056 11688 26108 11694
rect 26056 11630 26108 11636
rect 26068 11354 26096 11630
rect 26056 11348 26108 11354
rect 26056 11290 26108 11296
rect 26068 10810 26096 11290
rect 26160 11150 26188 11766
rect 26344 11354 26372 12174
rect 26436 12102 26464 12650
rect 26424 12096 26476 12102
rect 26424 12038 26476 12044
rect 26528 11762 26556 12786
rect 26620 12442 26648 13126
rect 26712 12918 26740 13246
rect 26700 12912 26752 12918
rect 26700 12854 26752 12860
rect 26608 12436 26660 12442
rect 26608 12378 26660 12384
rect 26516 11756 26568 11762
rect 26516 11698 26568 11704
rect 26804 11694 26832 15422
rect 27080 15162 27108 16050
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 26882 15056 26938 15065
rect 26882 14991 26884 15000
rect 26936 14991 26938 15000
rect 27068 15020 27120 15026
rect 26884 14962 26936 14968
rect 27068 14962 27120 14968
rect 26976 14952 27028 14958
rect 26976 14894 27028 14900
rect 26988 13938 27016 14894
rect 27080 14618 27108 14962
rect 27068 14612 27120 14618
rect 27068 14554 27120 14560
rect 27066 14104 27122 14113
rect 27066 14039 27068 14048
rect 27120 14039 27122 14048
rect 27068 14010 27120 14016
rect 26976 13932 27028 13938
rect 26976 13874 27028 13880
rect 26884 13456 26936 13462
rect 26884 13398 26936 13404
rect 26896 12986 26924 13398
rect 26884 12980 26936 12986
rect 26884 12922 26936 12928
rect 26988 12850 27016 13874
rect 26976 12844 27028 12850
rect 26976 12786 27028 12792
rect 27068 12436 27120 12442
rect 27068 12378 27120 12384
rect 27080 12170 27108 12378
rect 27068 12164 27120 12170
rect 27068 12106 27120 12112
rect 26792 11688 26844 11694
rect 26792 11630 26844 11636
rect 26516 11552 26568 11558
rect 26516 11494 26568 11500
rect 26700 11552 26752 11558
rect 26700 11494 26752 11500
rect 26528 11354 26556 11494
rect 26332 11348 26384 11354
rect 26332 11290 26384 11296
rect 26516 11348 26568 11354
rect 26516 11290 26568 11296
rect 26148 11144 26200 11150
rect 26148 11086 26200 11092
rect 26056 10804 26108 10810
rect 26056 10746 26108 10752
rect 25596 10668 25648 10674
rect 25596 10610 25648 10616
rect 25504 10600 25556 10606
rect 26712 10577 26740 11494
rect 27172 11082 27200 22578
rect 27264 17270 27292 22714
rect 27540 21690 27568 23072
rect 27908 22001 27936 30534
rect 28172 28484 28224 28490
rect 28172 28426 28224 28432
rect 27988 28416 28040 28422
rect 27988 28358 28040 28364
rect 28000 28218 28028 28358
rect 27988 28212 28040 28218
rect 27988 28154 28040 28160
rect 28184 28014 28212 28426
rect 28172 28008 28224 28014
rect 28172 27950 28224 27956
rect 27988 27328 28040 27334
rect 27986 27296 27988 27305
rect 28040 27296 28042 27305
rect 27986 27231 28042 27240
rect 28184 26042 28212 27950
rect 28172 26036 28224 26042
rect 28224 25996 28304 26024
rect 28172 25978 28224 25984
rect 27988 25288 28040 25294
rect 27988 25230 28040 25236
rect 28000 23798 28028 25230
rect 28080 25220 28132 25226
rect 28080 25162 28132 25168
rect 28092 24954 28120 25162
rect 28080 24948 28132 24954
rect 28080 24890 28132 24896
rect 28080 24608 28132 24614
rect 28080 24550 28132 24556
rect 28172 24608 28224 24614
rect 28172 24550 28224 24556
rect 28092 24410 28120 24550
rect 28080 24404 28132 24410
rect 28080 24346 28132 24352
rect 28184 24274 28212 24550
rect 28172 24268 28224 24274
rect 28172 24210 28224 24216
rect 28080 24200 28132 24206
rect 28080 24142 28132 24148
rect 27988 23792 28040 23798
rect 27988 23734 28040 23740
rect 27986 23624 28042 23633
rect 27986 23559 28042 23568
rect 27710 21992 27766 22001
rect 27620 21956 27672 21962
rect 27710 21927 27766 21936
rect 27894 21992 27950 22001
rect 27894 21927 27950 21936
rect 27620 21898 27672 21904
rect 27632 21690 27660 21898
rect 27528 21684 27580 21690
rect 27528 21626 27580 21632
rect 27620 21684 27672 21690
rect 27620 21626 27672 21632
rect 27436 21616 27488 21622
rect 27436 21558 27488 21564
rect 27448 21146 27476 21558
rect 27540 21418 27568 21626
rect 27528 21412 27580 21418
rect 27528 21354 27580 21360
rect 27436 21140 27488 21146
rect 27436 21082 27488 21088
rect 27448 20602 27476 21082
rect 27528 20800 27580 20806
rect 27528 20742 27580 20748
rect 27436 20596 27488 20602
rect 27436 20538 27488 20544
rect 27434 19408 27490 19417
rect 27434 19343 27490 19352
rect 27344 19168 27396 19174
rect 27344 19110 27396 19116
rect 27356 18970 27384 19110
rect 27448 18970 27476 19343
rect 27344 18964 27396 18970
rect 27344 18906 27396 18912
rect 27436 18964 27488 18970
rect 27436 18906 27488 18912
rect 27356 18834 27384 18906
rect 27344 18828 27396 18834
rect 27344 18770 27396 18776
rect 27356 17746 27384 18770
rect 27436 18760 27488 18766
rect 27436 18702 27488 18708
rect 27448 18358 27476 18702
rect 27436 18352 27488 18358
rect 27436 18294 27488 18300
rect 27344 17740 27396 17746
rect 27344 17682 27396 17688
rect 27252 17264 27304 17270
rect 27252 17206 27304 17212
rect 27344 17128 27396 17134
rect 27344 17070 27396 17076
rect 27356 16590 27384 17070
rect 27344 16584 27396 16590
rect 27344 16526 27396 16532
rect 27436 16448 27488 16454
rect 27342 16416 27398 16425
rect 27436 16390 27488 16396
rect 27342 16351 27398 16360
rect 27252 15972 27304 15978
rect 27252 15914 27304 15920
rect 27264 15570 27292 15914
rect 27252 15564 27304 15570
rect 27252 15506 27304 15512
rect 27356 14362 27384 16351
rect 27448 15570 27476 16390
rect 27436 15564 27488 15570
rect 27436 15506 27488 15512
rect 27448 14482 27476 15506
rect 27436 14476 27488 14482
rect 27436 14418 27488 14424
rect 27356 14334 27476 14362
rect 27252 13864 27304 13870
rect 27252 13806 27304 13812
rect 27264 13530 27292 13806
rect 27252 13524 27304 13530
rect 27252 13466 27304 13472
rect 27264 13326 27292 13466
rect 27342 13424 27398 13433
rect 27342 13359 27398 13368
rect 27356 13326 27384 13359
rect 27252 13320 27304 13326
rect 27252 13262 27304 13268
rect 27344 13320 27396 13326
rect 27344 13262 27396 13268
rect 27356 12918 27384 13262
rect 27344 12912 27396 12918
rect 27344 12854 27396 12860
rect 27252 12844 27304 12850
rect 27252 12786 27304 12792
rect 27264 12442 27292 12786
rect 27252 12436 27304 12442
rect 27252 12378 27304 12384
rect 27252 11892 27304 11898
rect 27252 11834 27304 11840
rect 27160 11076 27212 11082
rect 27160 11018 27212 11024
rect 26976 11008 27028 11014
rect 26976 10950 27028 10956
rect 26988 10810 27016 10950
rect 26976 10804 27028 10810
rect 26976 10746 27028 10752
rect 25504 10542 25556 10548
rect 26698 10568 26754 10577
rect 25516 10198 25544 10542
rect 26698 10503 26754 10512
rect 26792 10260 26844 10266
rect 26792 10202 26844 10208
rect 25504 10192 25556 10198
rect 25504 10134 25556 10140
rect 26804 10130 26832 10202
rect 26792 10124 26844 10130
rect 26792 10066 26844 10072
rect 26988 10062 27016 10746
rect 27172 10441 27200 11018
rect 27158 10432 27214 10441
rect 27158 10367 27214 10376
rect 27160 10260 27212 10266
rect 27160 10202 27212 10208
rect 27172 10062 27200 10202
rect 26976 10056 27028 10062
rect 26976 9998 27028 10004
rect 27160 10056 27212 10062
rect 27160 9998 27212 10004
rect 27264 9926 27292 11834
rect 27448 11150 27476 14334
rect 27540 13530 27568 20742
rect 27620 18284 27672 18290
rect 27620 18226 27672 18232
rect 27632 17746 27660 18226
rect 27620 17740 27672 17746
rect 27620 17682 27672 17688
rect 27724 17678 27752 21927
rect 27896 21480 27948 21486
rect 27896 21422 27948 21428
rect 27804 20868 27856 20874
rect 27804 20810 27856 20816
rect 27816 20602 27844 20810
rect 27804 20596 27856 20602
rect 27804 20538 27856 20544
rect 27908 20534 27936 21422
rect 27896 20528 27948 20534
rect 27896 20470 27948 20476
rect 27804 20256 27856 20262
rect 27804 20198 27856 20204
rect 27816 19242 27844 20198
rect 27804 19236 27856 19242
rect 27804 19178 27856 19184
rect 27896 19168 27948 19174
rect 27896 19110 27948 19116
rect 27908 18698 27936 19110
rect 27896 18692 27948 18698
rect 27896 18634 27948 18640
rect 27712 17672 27764 17678
rect 27712 17614 27764 17620
rect 27712 17536 27764 17542
rect 27712 17478 27764 17484
rect 27724 14249 27752 17478
rect 27804 17128 27856 17134
rect 27804 17070 27856 17076
rect 27816 16046 27844 17070
rect 27804 16040 27856 16046
rect 27804 15982 27856 15988
rect 27816 15502 27844 15982
rect 27804 15496 27856 15502
rect 27804 15438 27856 15444
rect 27710 14240 27766 14249
rect 27710 14175 27766 14184
rect 27816 13938 27844 15438
rect 28000 14906 28028 23559
rect 28092 19514 28120 24142
rect 28172 23316 28224 23322
rect 28172 23258 28224 23264
rect 28184 22642 28212 23258
rect 28172 22636 28224 22642
rect 28172 22578 28224 22584
rect 28184 21486 28212 22578
rect 28172 21480 28224 21486
rect 28172 21422 28224 21428
rect 28276 20806 28304 25996
rect 28460 24954 28488 32302
rect 28552 32026 28580 32370
rect 28540 32020 28592 32026
rect 28540 31962 28592 31968
rect 28552 31822 28580 31962
rect 28540 31816 28592 31822
rect 28540 31758 28592 31764
rect 28736 31754 28764 32846
rect 28644 31726 28764 31754
rect 28908 31748 28960 31754
rect 28540 29572 28592 29578
rect 28540 29514 28592 29520
rect 28552 29306 28580 29514
rect 28540 29300 28592 29306
rect 28540 29242 28592 29248
rect 28448 24948 28500 24954
rect 28448 24890 28500 24896
rect 28540 24812 28592 24818
rect 28540 24754 28592 24760
rect 28356 24608 28408 24614
rect 28356 24550 28408 24556
rect 28368 24070 28396 24550
rect 28552 24449 28580 24754
rect 28538 24440 28594 24449
rect 28448 24404 28500 24410
rect 28538 24375 28540 24384
rect 28448 24346 28500 24352
rect 28592 24375 28594 24384
rect 28540 24346 28592 24352
rect 28356 24064 28408 24070
rect 28354 24032 28356 24041
rect 28408 24032 28410 24041
rect 28354 23967 28410 23976
rect 28356 21344 28408 21350
rect 28356 21286 28408 21292
rect 28368 20913 28396 21286
rect 28354 20904 28410 20913
rect 28354 20839 28410 20848
rect 28264 20800 28316 20806
rect 28264 20742 28316 20748
rect 28356 20392 28408 20398
rect 28356 20334 28408 20340
rect 28368 19718 28396 20334
rect 28356 19712 28408 19718
rect 28356 19654 28408 19660
rect 28080 19508 28132 19514
rect 28080 19450 28132 19456
rect 28264 19440 28316 19446
rect 28264 19382 28316 19388
rect 28276 17814 28304 19382
rect 28264 17808 28316 17814
rect 28264 17750 28316 17756
rect 28264 17604 28316 17610
rect 28264 17546 28316 17552
rect 28080 16584 28132 16590
rect 28080 16526 28132 16532
rect 27908 14878 28028 14906
rect 27908 14618 27936 14878
rect 27988 14816 28040 14822
rect 27988 14758 28040 14764
rect 27896 14612 27948 14618
rect 27896 14554 27948 14560
rect 28000 14414 28028 14758
rect 27988 14408 28040 14414
rect 27894 14376 27950 14385
rect 27988 14350 28040 14356
rect 27894 14311 27950 14320
rect 27908 14074 27936 14311
rect 27988 14272 28040 14278
rect 27988 14214 28040 14220
rect 27896 14068 27948 14074
rect 27896 14010 27948 14016
rect 27804 13932 27856 13938
rect 27804 13874 27856 13880
rect 27528 13524 27580 13530
rect 27528 13466 27580 13472
rect 27540 12306 27568 13466
rect 27896 13320 27948 13326
rect 27896 13262 27948 13268
rect 27804 13252 27856 13258
rect 27804 13194 27856 13200
rect 27816 12986 27844 13194
rect 27804 12980 27856 12986
rect 27804 12922 27856 12928
rect 27816 12730 27844 12922
rect 27908 12866 27936 13262
rect 28000 12968 28028 14214
rect 28092 13394 28120 16526
rect 28172 14884 28224 14890
rect 28172 14826 28224 14832
rect 28184 14346 28212 14826
rect 28276 14482 28304 17546
rect 28368 14906 28396 19654
rect 28460 19394 28488 24346
rect 28644 22030 28672 31726
rect 28908 31690 28960 31696
rect 28816 31476 28868 31482
rect 28816 31418 28868 31424
rect 28828 30734 28856 31418
rect 28920 30802 28948 31690
rect 28908 30796 28960 30802
rect 28908 30738 28960 30744
rect 28816 30728 28868 30734
rect 28816 30670 28868 30676
rect 29000 30660 29052 30666
rect 29000 30602 29052 30608
rect 29012 30122 29040 30602
rect 29000 30116 29052 30122
rect 29000 30058 29052 30064
rect 29092 30048 29144 30054
rect 29092 29990 29144 29996
rect 29104 29510 29132 29990
rect 29092 29504 29144 29510
rect 29092 29446 29144 29452
rect 29104 29102 29132 29446
rect 29092 29096 29144 29102
rect 29092 29038 29144 29044
rect 29000 28076 29052 28082
rect 29000 28018 29052 28024
rect 29012 27878 29040 28018
rect 29000 27872 29052 27878
rect 29000 27814 29052 27820
rect 28724 27532 28776 27538
rect 28724 27474 28776 27480
rect 28736 27334 28764 27474
rect 28724 27328 28776 27334
rect 28724 27270 28776 27276
rect 28736 26382 28764 27270
rect 28906 26480 28962 26489
rect 28906 26415 28908 26424
rect 28960 26415 28962 26424
rect 28908 26386 28960 26392
rect 28724 26376 28776 26382
rect 28724 26318 28776 26324
rect 29012 25770 29040 27814
rect 29092 27464 29144 27470
rect 29092 27406 29144 27412
rect 29000 25764 29052 25770
rect 29000 25706 29052 25712
rect 28724 24744 28776 24750
rect 28724 24686 28776 24692
rect 28908 24744 28960 24750
rect 28908 24686 28960 24692
rect 28736 24410 28764 24686
rect 28816 24608 28868 24614
rect 28816 24550 28868 24556
rect 28724 24404 28776 24410
rect 28724 24346 28776 24352
rect 28724 24200 28776 24206
rect 28724 24142 28776 24148
rect 28736 23633 28764 24142
rect 28828 24138 28856 24550
rect 28920 24206 28948 24686
rect 29000 24336 29052 24342
rect 29000 24278 29052 24284
rect 28908 24200 28960 24206
rect 28908 24142 28960 24148
rect 29012 24138 29040 24278
rect 28816 24132 28868 24138
rect 28816 24074 28868 24080
rect 29000 24132 29052 24138
rect 29000 24074 29052 24080
rect 28908 23724 28960 23730
rect 28908 23666 28960 23672
rect 28722 23624 28778 23633
rect 28722 23559 28778 23568
rect 28920 23322 28948 23666
rect 28908 23316 28960 23322
rect 28908 23258 28960 23264
rect 29012 22137 29040 24074
rect 29104 22506 29132 27406
rect 29196 27282 29224 33254
rect 29288 30734 29316 33458
rect 29552 33380 29604 33386
rect 29552 33322 29604 33328
rect 29564 32298 29592 33322
rect 29840 33114 29868 33458
rect 32128 33448 32180 33454
rect 32128 33390 32180 33396
rect 32404 33448 32456 33454
rect 32404 33390 32456 33396
rect 31024 33380 31076 33386
rect 31024 33322 31076 33328
rect 29828 33108 29880 33114
rect 29828 33050 29880 33056
rect 29840 32994 29868 33050
rect 29840 32966 29960 32994
rect 29644 32904 29696 32910
rect 29644 32846 29696 32852
rect 29656 32502 29684 32846
rect 29828 32836 29880 32842
rect 29828 32778 29880 32784
rect 29644 32496 29696 32502
rect 29644 32438 29696 32444
rect 29552 32292 29604 32298
rect 29552 32234 29604 32240
rect 29460 31816 29512 31822
rect 29460 31758 29512 31764
rect 29276 30728 29328 30734
rect 29276 30670 29328 30676
rect 29288 27538 29316 30670
rect 29368 29776 29420 29782
rect 29368 29718 29420 29724
rect 29380 29306 29408 29718
rect 29368 29300 29420 29306
rect 29368 29242 29420 29248
rect 29368 28620 29420 28626
rect 29368 28562 29420 28568
rect 29380 28422 29408 28562
rect 29368 28416 29420 28422
rect 29366 28384 29368 28393
rect 29420 28384 29422 28393
rect 29366 28319 29422 28328
rect 29276 27532 29328 27538
rect 29276 27474 29328 27480
rect 29196 27254 29316 27282
rect 29184 27124 29236 27130
rect 29184 27066 29236 27072
rect 29196 26382 29224 27066
rect 29184 26376 29236 26382
rect 29184 26318 29236 26324
rect 29184 24948 29236 24954
rect 29184 24890 29236 24896
rect 29196 24290 29224 24890
rect 29288 24410 29316 27254
rect 29276 24404 29328 24410
rect 29276 24346 29328 24352
rect 29196 24262 29316 24290
rect 29288 24138 29316 24262
rect 29276 24132 29328 24138
rect 29276 24074 29328 24080
rect 29288 22982 29316 24074
rect 29472 23186 29500 31758
rect 29656 31346 29684 32438
rect 29840 32026 29868 32778
rect 29828 32020 29880 32026
rect 29828 31962 29880 31968
rect 29932 31890 29960 32966
rect 31036 32842 31064 33322
rect 32140 32910 32168 33390
rect 32416 33114 32444 33390
rect 32404 33108 32456 33114
rect 32404 33050 32456 33056
rect 32772 32972 32824 32978
rect 32772 32914 32824 32920
rect 32128 32904 32180 32910
rect 32128 32846 32180 32852
rect 31024 32836 31076 32842
rect 31024 32778 31076 32784
rect 30288 32292 30340 32298
rect 30288 32234 30340 32240
rect 29920 31884 29972 31890
rect 29920 31826 29972 31832
rect 30104 31884 30156 31890
rect 30104 31826 30156 31832
rect 29644 31340 29696 31346
rect 29644 31282 29696 31288
rect 29920 29844 29972 29850
rect 29920 29786 29972 29792
rect 29552 29640 29604 29646
rect 29552 29582 29604 29588
rect 29460 23180 29512 23186
rect 29460 23122 29512 23128
rect 29564 23118 29592 29582
rect 29932 29578 29960 29786
rect 29828 29572 29880 29578
rect 29828 29514 29880 29520
rect 29920 29572 29972 29578
rect 29920 29514 29972 29520
rect 29840 29306 29868 29514
rect 29828 29300 29880 29306
rect 29828 29242 29880 29248
rect 29736 29164 29788 29170
rect 29736 29106 29788 29112
rect 29748 28762 29776 29106
rect 29736 28756 29788 28762
rect 29736 28698 29788 28704
rect 29840 28558 29868 29242
rect 29828 28552 29880 28558
rect 29828 28494 29880 28500
rect 29932 28098 29960 29514
rect 29840 28070 29960 28098
rect 29644 27328 29696 27334
rect 29644 27270 29696 27276
rect 29656 26994 29684 27270
rect 29644 26988 29696 26994
rect 29644 26930 29696 26936
rect 29736 24812 29788 24818
rect 29840 24800 29868 28070
rect 29920 27940 29972 27946
rect 29920 27882 29972 27888
rect 29932 27334 29960 27882
rect 30116 27538 30144 31826
rect 30300 30802 30328 32234
rect 32784 31890 32812 32914
rect 32772 31884 32824 31890
rect 32772 31826 32824 31832
rect 30380 31680 30432 31686
rect 30380 31622 30432 31628
rect 30840 31680 30892 31686
rect 30840 31622 30892 31628
rect 30392 31414 30420 31622
rect 30852 31482 30880 31622
rect 30840 31476 30892 31482
rect 30840 31418 30892 31424
rect 30380 31408 30432 31414
rect 30380 31350 30432 31356
rect 30288 30796 30340 30802
rect 30288 30738 30340 30744
rect 30852 30734 30880 31418
rect 30840 30728 30892 30734
rect 31208 30728 31260 30734
rect 30840 30670 30892 30676
rect 31128 30688 31208 30716
rect 30196 30048 30248 30054
rect 30196 29990 30248 29996
rect 30104 27532 30156 27538
rect 30104 27474 30156 27480
rect 30116 27402 30144 27474
rect 30104 27396 30156 27402
rect 30104 27338 30156 27344
rect 29920 27328 29972 27334
rect 29920 27270 29972 27276
rect 30012 27328 30064 27334
rect 30012 27270 30064 27276
rect 30024 27130 30052 27270
rect 30012 27124 30064 27130
rect 30012 27066 30064 27072
rect 30104 27056 30156 27062
rect 30104 26998 30156 27004
rect 30116 26450 30144 26998
rect 30104 26444 30156 26450
rect 30104 26386 30156 26392
rect 30104 25832 30156 25838
rect 30104 25774 30156 25780
rect 30116 25158 30144 25774
rect 30208 25362 30236 29990
rect 30380 26988 30432 26994
rect 30380 26930 30432 26936
rect 30288 26784 30340 26790
rect 30288 26726 30340 26732
rect 30196 25356 30248 25362
rect 30196 25298 30248 25304
rect 30104 25152 30156 25158
rect 30104 25094 30156 25100
rect 30116 24954 30144 25094
rect 30104 24948 30156 24954
rect 30104 24890 30156 24896
rect 30300 24818 30328 26726
rect 29788 24772 29868 24800
rect 30012 24812 30064 24818
rect 29736 24754 29788 24760
rect 30012 24754 30064 24760
rect 30288 24812 30340 24818
rect 30288 24754 30340 24760
rect 29748 24614 29776 24754
rect 29736 24608 29788 24614
rect 29736 24550 29788 24556
rect 29644 24200 29696 24206
rect 29644 24142 29696 24148
rect 29656 23866 29684 24142
rect 29644 23860 29696 23866
rect 29644 23802 29696 23808
rect 29644 23520 29696 23526
rect 29644 23462 29696 23468
rect 29552 23112 29604 23118
rect 29552 23054 29604 23060
rect 29276 22976 29328 22982
rect 29276 22918 29328 22924
rect 29288 22778 29316 22918
rect 29276 22772 29328 22778
rect 29276 22714 29328 22720
rect 29184 22704 29236 22710
rect 29184 22646 29236 22652
rect 29092 22500 29144 22506
rect 29092 22442 29144 22448
rect 29092 22228 29144 22234
rect 29196 22216 29224 22646
rect 29288 22438 29316 22714
rect 29564 22642 29592 23054
rect 29552 22636 29604 22642
rect 29552 22578 29604 22584
rect 29276 22432 29328 22438
rect 29274 22400 29276 22409
rect 29460 22432 29512 22438
rect 29328 22400 29330 22409
rect 29460 22374 29512 22380
rect 29274 22335 29330 22344
rect 29144 22188 29224 22216
rect 29092 22170 29144 22176
rect 29368 22160 29420 22166
rect 28998 22128 29054 22137
rect 28998 22063 29054 22072
rect 29196 22120 29368 22148
rect 28540 22024 28592 22030
rect 28540 21966 28592 21972
rect 28632 22024 28684 22030
rect 28684 21984 28948 22012
rect 28632 21966 28684 21972
rect 28552 21690 28580 21966
rect 28920 21894 28948 21984
rect 28816 21888 28868 21894
rect 28816 21830 28868 21836
rect 28908 21888 28960 21894
rect 28908 21830 28960 21836
rect 29000 21888 29052 21894
rect 29196 21876 29224 22120
rect 29368 22102 29420 22108
rect 29472 22098 29500 22374
rect 29460 22092 29512 22098
rect 29460 22034 29512 22040
rect 29276 22024 29328 22030
rect 29276 21966 29328 21972
rect 29368 22024 29420 22030
rect 29368 21966 29420 21972
rect 29552 22024 29604 22030
rect 29552 21966 29604 21972
rect 29052 21848 29224 21876
rect 29288 21865 29316 21966
rect 29274 21856 29330 21865
rect 29000 21830 29052 21836
rect 28828 21690 28856 21830
rect 29274 21791 29330 21800
rect 29182 21720 29238 21729
rect 28540 21684 28592 21690
rect 28540 21626 28592 21632
rect 28816 21684 28868 21690
rect 29182 21655 29238 21664
rect 28816 21626 28868 21632
rect 28816 21548 28868 21554
rect 28816 21490 28868 21496
rect 28908 21548 28960 21554
rect 28908 21490 28960 21496
rect 28724 21480 28776 21486
rect 28724 21422 28776 21428
rect 28736 20534 28764 21422
rect 28724 20528 28776 20534
rect 28724 20470 28776 20476
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 28460 19366 28672 19394
rect 28540 19304 28592 19310
rect 28540 19246 28592 19252
rect 28552 18766 28580 19246
rect 28540 18760 28592 18766
rect 28540 18702 28592 18708
rect 28448 18624 28500 18630
rect 28644 18612 28672 19366
rect 28736 18698 28764 19450
rect 28724 18692 28776 18698
rect 28724 18634 28776 18640
rect 28448 18566 28500 18572
rect 28552 18584 28672 18612
rect 28460 17678 28488 18566
rect 28552 18222 28580 18584
rect 28540 18216 28592 18222
rect 28540 18158 28592 18164
rect 28448 17672 28500 17678
rect 28448 17614 28500 17620
rect 28448 16108 28500 16114
rect 28448 16050 28500 16056
rect 28460 15706 28488 16050
rect 28448 15700 28500 15706
rect 28448 15642 28500 15648
rect 28552 15026 28580 18158
rect 28724 18080 28776 18086
rect 28724 18022 28776 18028
rect 28632 17128 28684 17134
rect 28632 17070 28684 17076
rect 28644 16794 28672 17070
rect 28632 16788 28684 16794
rect 28632 16730 28684 16736
rect 28736 16590 28764 18022
rect 28828 17490 28856 21490
rect 28920 20806 28948 21490
rect 28908 20800 28960 20806
rect 28908 20742 28960 20748
rect 28920 20602 28948 20742
rect 29196 20618 29224 21655
rect 29380 21622 29408 21966
rect 29460 21888 29512 21894
rect 29460 21830 29512 21836
rect 29368 21616 29420 21622
rect 29368 21558 29420 21564
rect 29380 21298 29408 21558
rect 29472 21554 29500 21830
rect 29564 21690 29592 21966
rect 29656 21962 29684 23462
rect 29748 22574 29776 24550
rect 29920 23860 29972 23866
rect 29920 23802 29972 23808
rect 29932 23118 29960 23802
rect 29920 23112 29972 23118
rect 29920 23054 29972 23060
rect 29736 22568 29788 22574
rect 29734 22536 29736 22545
rect 29788 22536 29790 22545
rect 29734 22471 29790 22480
rect 29736 22432 29788 22438
rect 29736 22374 29788 22380
rect 29644 21956 29696 21962
rect 29644 21898 29696 21904
rect 29552 21684 29604 21690
rect 29552 21626 29604 21632
rect 29460 21548 29512 21554
rect 29460 21490 29512 21496
rect 29380 21270 29500 21298
rect 29368 21140 29420 21146
rect 29368 21082 29420 21088
rect 28908 20596 28960 20602
rect 29196 20590 29316 20618
rect 29380 20602 29408 21082
rect 29472 21078 29500 21270
rect 29460 21072 29512 21078
rect 29460 21014 29512 21020
rect 29656 21010 29684 21898
rect 29748 21690 29776 22374
rect 29736 21684 29788 21690
rect 29736 21626 29788 21632
rect 29920 21684 29972 21690
rect 29920 21626 29972 21632
rect 29644 21004 29696 21010
rect 29644 20946 29696 20952
rect 29748 20942 29776 21626
rect 29828 21412 29880 21418
rect 29828 21354 29880 21360
rect 29460 20936 29512 20942
rect 29460 20878 29512 20884
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 28908 20538 28960 20544
rect 29092 19508 29144 19514
rect 29092 19450 29144 19456
rect 29000 19304 29052 19310
rect 29000 19246 29052 19252
rect 29012 18970 29040 19246
rect 29104 19242 29132 19450
rect 29184 19440 29236 19446
rect 29184 19382 29236 19388
rect 29092 19236 29144 19242
rect 29092 19178 29144 19184
rect 29000 18964 29052 18970
rect 29000 18906 29052 18912
rect 28908 18624 28960 18630
rect 29012 18612 29040 18906
rect 29196 18902 29224 19382
rect 29184 18896 29236 18902
rect 29184 18838 29236 18844
rect 29196 18766 29224 18838
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 28960 18584 29040 18612
rect 28908 18566 28960 18572
rect 29092 18420 29144 18426
rect 29196 18408 29224 18702
rect 29144 18380 29224 18408
rect 29092 18362 29144 18368
rect 28920 18290 29132 18306
rect 28908 18284 29144 18290
rect 28960 18278 29092 18284
rect 28908 18226 28960 18232
rect 29092 18226 29144 18232
rect 29196 17882 29224 18380
rect 29288 18086 29316 20590
rect 29368 20596 29420 20602
rect 29368 20538 29420 20544
rect 29368 19168 29420 19174
rect 29368 19110 29420 19116
rect 29380 18698 29408 19110
rect 29368 18692 29420 18698
rect 29368 18634 29420 18640
rect 29276 18080 29328 18086
rect 29276 18022 29328 18028
rect 29184 17876 29236 17882
rect 29184 17818 29236 17824
rect 29000 17536 29052 17542
rect 28828 17484 29000 17490
rect 28828 17478 29052 17484
rect 28828 17462 29040 17478
rect 28920 16590 28948 17462
rect 29276 16992 29328 16998
rect 29276 16934 29328 16940
rect 29000 16652 29052 16658
rect 29000 16594 29052 16600
rect 28724 16584 28776 16590
rect 28724 16526 28776 16532
rect 28908 16584 28960 16590
rect 28908 16526 28960 16532
rect 28920 16182 28948 16526
rect 28908 16176 28960 16182
rect 28908 16118 28960 16124
rect 29012 15910 29040 16594
rect 29288 16454 29316 16934
rect 29092 16448 29144 16454
rect 29092 16390 29144 16396
rect 29276 16448 29328 16454
rect 29276 16390 29328 16396
rect 29104 15978 29132 16390
rect 29288 16182 29316 16390
rect 29276 16176 29328 16182
rect 29276 16118 29328 16124
rect 29472 15978 29500 20878
rect 29840 20466 29868 21354
rect 29932 20942 29960 21626
rect 30024 21146 30052 24754
rect 30104 22636 30156 22642
rect 30104 22578 30156 22584
rect 30012 21140 30064 21146
rect 30012 21082 30064 21088
rect 29920 20936 29972 20942
rect 29920 20878 29972 20884
rect 29828 20460 29880 20466
rect 29828 20402 29880 20408
rect 29920 19508 29972 19514
rect 29920 19450 29972 19456
rect 29644 19372 29696 19378
rect 29644 19314 29696 19320
rect 29656 18834 29684 19314
rect 29828 19304 29880 19310
rect 29828 19246 29880 19252
rect 29644 18828 29696 18834
rect 29644 18770 29696 18776
rect 29552 18624 29604 18630
rect 29552 18566 29604 18572
rect 29564 18358 29592 18566
rect 29656 18426 29684 18770
rect 29644 18420 29696 18426
rect 29644 18362 29696 18368
rect 29552 18352 29604 18358
rect 29552 18294 29604 18300
rect 29564 17746 29592 18294
rect 29840 18086 29868 19246
rect 29644 18080 29696 18086
rect 29644 18022 29696 18028
rect 29828 18080 29880 18086
rect 29828 18022 29880 18028
rect 29552 17740 29604 17746
rect 29552 17682 29604 17688
rect 29656 17678 29684 18022
rect 29840 17678 29868 18022
rect 29644 17672 29696 17678
rect 29644 17614 29696 17620
rect 29828 17672 29880 17678
rect 29828 17614 29880 17620
rect 29552 16584 29604 16590
rect 29552 16526 29604 16532
rect 29564 16250 29592 16526
rect 29552 16244 29604 16250
rect 29552 16186 29604 16192
rect 29092 15972 29144 15978
rect 29092 15914 29144 15920
rect 29460 15972 29512 15978
rect 29460 15914 29512 15920
rect 29000 15904 29052 15910
rect 29000 15846 29052 15852
rect 29184 15904 29236 15910
rect 29184 15846 29236 15852
rect 29092 15564 29144 15570
rect 29092 15506 29144 15512
rect 28908 15088 28960 15094
rect 28908 15030 28960 15036
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 28724 15020 28776 15026
rect 28724 14962 28776 14968
rect 28368 14878 28580 14906
rect 28448 14816 28500 14822
rect 28368 14764 28448 14770
rect 28368 14758 28500 14764
rect 28368 14742 28488 14758
rect 28264 14476 28316 14482
rect 28264 14418 28316 14424
rect 28172 14340 28224 14346
rect 28172 14282 28224 14288
rect 28264 14340 28316 14346
rect 28264 14282 28316 14288
rect 28080 13388 28132 13394
rect 28080 13330 28132 13336
rect 28000 12940 28120 12968
rect 27908 12838 28028 12866
rect 27816 12702 27936 12730
rect 27528 12300 27580 12306
rect 27528 12242 27580 12248
rect 27908 12238 27936 12702
rect 27896 12232 27948 12238
rect 27896 12174 27948 12180
rect 27528 12096 27580 12102
rect 27528 12038 27580 12044
rect 27436 11144 27488 11150
rect 27436 11086 27488 11092
rect 27540 11082 27568 12038
rect 28000 11778 28028 12838
rect 27712 11756 27764 11762
rect 27712 11698 27764 11704
rect 27908 11750 28028 11778
rect 27620 11688 27672 11694
rect 27620 11630 27672 11636
rect 27632 11218 27660 11630
rect 27724 11286 27752 11698
rect 27712 11280 27764 11286
rect 27712 11222 27764 11228
rect 27620 11212 27672 11218
rect 27620 11154 27672 11160
rect 27804 11212 27856 11218
rect 27804 11154 27856 11160
rect 27712 11144 27764 11150
rect 27712 11086 27764 11092
rect 27528 11076 27580 11082
rect 27528 11018 27580 11024
rect 27620 11076 27672 11082
rect 27620 11018 27672 11024
rect 27528 10668 27580 10674
rect 27528 10610 27580 10616
rect 27540 10266 27568 10610
rect 27528 10260 27580 10266
rect 27528 10202 27580 10208
rect 27252 9920 27304 9926
rect 27252 9862 27304 9868
rect 26608 9648 26660 9654
rect 26514 9616 26570 9625
rect 26884 9648 26936 9654
rect 26660 9608 26884 9636
rect 26608 9590 26660 9596
rect 26884 9590 26936 9596
rect 26514 9551 26516 9560
rect 26568 9551 26570 9560
rect 26516 9522 26568 9528
rect 25504 9512 25556 9518
rect 25504 9454 25556 9460
rect 26330 9480 26386 9489
rect 25412 9444 25464 9450
rect 25412 9386 25464 9392
rect 25516 9382 25544 9454
rect 26330 9415 26332 9424
rect 26384 9415 26386 9424
rect 26332 9386 26384 9392
rect 25504 9376 25556 9382
rect 25504 9318 25556 9324
rect 26792 9376 26844 9382
rect 26792 9318 26844 9324
rect 25320 9172 25372 9178
rect 25320 9114 25372 9120
rect 25136 8288 25188 8294
rect 25136 8230 25188 8236
rect 25148 7342 25176 8230
rect 25228 7472 25280 7478
rect 25228 7414 25280 7420
rect 25136 7336 25188 7342
rect 25136 7278 25188 7284
rect 25240 7206 25268 7414
rect 25516 7410 25544 9318
rect 26804 8634 26832 9318
rect 27160 9104 27212 9110
rect 27160 9046 27212 9052
rect 26792 8628 26844 8634
rect 26792 8570 26844 8576
rect 26884 8492 26936 8498
rect 26884 8434 26936 8440
rect 25976 7500 26188 7528
rect 25320 7404 25372 7410
rect 25320 7346 25372 7352
rect 25412 7404 25464 7410
rect 25412 7346 25464 7352
rect 25504 7404 25556 7410
rect 25504 7346 25556 7352
rect 25332 7274 25360 7346
rect 25320 7268 25372 7274
rect 25320 7210 25372 7216
rect 25228 7200 25280 7206
rect 25228 7142 25280 7148
rect 25240 7002 25268 7142
rect 25228 6996 25280 7002
rect 25148 6956 25228 6984
rect 25044 6928 25096 6934
rect 25044 6870 25096 6876
rect 24952 6724 25004 6730
rect 24952 6666 25004 6672
rect 24964 6254 24992 6666
rect 25056 6322 25084 6870
rect 25148 6322 25176 6956
rect 25228 6938 25280 6944
rect 25332 6934 25360 7210
rect 25320 6928 25372 6934
rect 25320 6870 25372 6876
rect 25228 6792 25280 6798
rect 25228 6734 25280 6740
rect 25044 6316 25096 6322
rect 25044 6258 25096 6264
rect 25136 6316 25188 6322
rect 25136 6258 25188 6264
rect 24952 6248 25004 6254
rect 24952 6190 25004 6196
rect 25240 6186 25268 6734
rect 25320 6656 25372 6662
rect 25320 6598 25372 6604
rect 25332 6458 25360 6598
rect 25320 6452 25372 6458
rect 25320 6394 25372 6400
rect 25228 6180 25280 6186
rect 25228 6122 25280 6128
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 25056 5778 25084 6054
rect 25044 5772 25096 5778
rect 25044 5714 25096 5720
rect 25240 5710 25268 6122
rect 25424 5914 25452 7346
rect 25976 6866 26004 7500
rect 26160 7410 26188 7500
rect 26056 7404 26108 7410
rect 26056 7346 26108 7352
rect 26148 7404 26200 7410
rect 26148 7346 26200 7352
rect 26068 7002 26096 7346
rect 26056 6996 26108 7002
rect 26056 6938 26108 6944
rect 26148 6996 26200 7002
rect 26148 6938 26200 6944
rect 25964 6860 26016 6866
rect 25964 6802 26016 6808
rect 26056 6724 26108 6730
rect 26056 6666 26108 6672
rect 25688 6656 25740 6662
rect 25688 6598 25740 6604
rect 25700 6254 25728 6598
rect 25688 6248 25740 6254
rect 25688 6190 25740 6196
rect 25412 5908 25464 5914
rect 25412 5850 25464 5856
rect 25228 5704 25280 5710
rect 25228 5646 25280 5652
rect 26068 5302 26096 6666
rect 26160 6458 26188 6938
rect 26896 6662 26924 8434
rect 27172 7750 27200 9046
rect 27264 9042 27292 9862
rect 27632 9654 27660 11018
rect 27724 10266 27752 11086
rect 27816 10266 27844 11154
rect 27712 10260 27764 10266
rect 27712 10202 27764 10208
rect 27804 10260 27856 10266
rect 27804 10202 27856 10208
rect 27908 9994 27936 11750
rect 27988 11620 28040 11626
rect 27988 11562 28040 11568
rect 28000 11150 28028 11562
rect 28092 11218 28120 12940
rect 28184 12889 28212 14282
rect 28276 14074 28304 14282
rect 28264 14068 28316 14074
rect 28264 14010 28316 14016
rect 28170 12880 28226 12889
rect 28170 12815 28226 12824
rect 28264 12096 28316 12102
rect 28264 12038 28316 12044
rect 28172 11824 28224 11830
rect 28172 11766 28224 11772
rect 28080 11212 28132 11218
rect 28080 11154 28132 11160
rect 27988 11144 28040 11150
rect 27988 11086 28040 11092
rect 28080 11008 28132 11014
rect 28080 10950 28132 10956
rect 28092 10062 28120 10950
rect 28184 10198 28212 11766
rect 28276 11665 28304 12038
rect 28368 11694 28396 14742
rect 28448 14000 28500 14006
rect 28448 13942 28500 13948
rect 28460 13530 28488 13942
rect 28448 13524 28500 13530
rect 28448 13466 28500 13472
rect 28552 12434 28580 14878
rect 28632 14884 28684 14890
rect 28632 14826 28684 14832
rect 28644 14550 28672 14826
rect 28736 14822 28764 14962
rect 28724 14816 28776 14822
rect 28724 14758 28776 14764
rect 28722 14648 28778 14657
rect 28722 14583 28778 14592
rect 28632 14544 28684 14550
rect 28632 14486 28684 14492
rect 28736 14482 28764 14583
rect 28724 14476 28776 14482
rect 28724 14418 28776 14424
rect 28632 14408 28684 14414
rect 28816 14408 28868 14414
rect 28632 14350 28684 14356
rect 28814 14376 28816 14385
rect 28868 14376 28870 14385
rect 28644 14249 28672 14350
rect 28920 14346 28948 15030
rect 28814 14311 28870 14320
rect 28908 14340 28960 14346
rect 28828 14278 28856 14311
rect 28908 14282 28960 14288
rect 28724 14272 28776 14278
rect 28630 14240 28686 14249
rect 28724 14214 28776 14220
rect 28816 14272 28868 14278
rect 28816 14214 28868 14220
rect 28630 14175 28686 14184
rect 28632 13252 28684 13258
rect 28632 13194 28684 13200
rect 28644 12646 28672 13194
rect 28632 12640 28684 12646
rect 28632 12582 28684 12588
rect 28460 12406 28580 12434
rect 28356 11688 28408 11694
rect 28262 11656 28318 11665
rect 28356 11630 28408 11636
rect 28262 11591 28318 11600
rect 28276 11014 28304 11591
rect 28264 11008 28316 11014
rect 28264 10950 28316 10956
rect 28262 10840 28318 10849
rect 28262 10775 28318 10784
rect 28172 10192 28224 10198
rect 28172 10134 28224 10140
rect 28080 10056 28132 10062
rect 28080 9998 28132 10004
rect 27896 9988 27948 9994
rect 27896 9930 27948 9936
rect 28276 9926 28304 10775
rect 28264 9920 28316 9926
rect 28264 9862 28316 9868
rect 27620 9648 27672 9654
rect 27620 9590 27672 9596
rect 28276 9586 28304 9862
rect 28264 9580 28316 9586
rect 28264 9522 28316 9528
rect 27804 9512 27856 9518
rect 27804 9454 27856 9460
rect 27816 9382 27844 9454
rect 28172 9444 28224 9450
rect 28172 9386 28224 9392
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 28080 9376 28132 9382
rect 28080 9318 28132 9324
rect 27816 9042 27844 9318
rect 27252 9036 27304 9042
rect 27252 8978 27304 8984
rect 27804 9036 27856 9042
rect 27804 8978 27856 8984
rect 27264 7886 27292 8978
rect 27816 8566 27844 8978
rect 28092 8974 28120 9318
rect 28080 8968 28132 8974
rect 28080 8910 28132 8916
rect 28092 8634 28120 8910
rect 28184 8906 28212 9386
rect 28460 9217 28488 12406
rect 28540 11348 28592 11354
rect 28540 11290 28592 11296
rect 28552 9926 28580 11290
rect 28644 11218 28672 12582
rect 28736 11762 28764 14214
rect 28816 14068 28868 14074
rect 28816 14010 28868 14016
rect 28828 13326 28856 14010
rect 28816 13320 28868 13326
rect 28816 13262 28868 13268
rect 29104 12434 29132 15506
rect 29196 15434 29224 15846
rect 29184 15428 29236 15434
rect 29184 15370 29236 15376
rect 29196 15026 29224 15370
rect 29276 15360 29328 15366
rect 29276 15302 29328 15308
rect 29184 15020 29236 15026
rect 29184 14962 29236 14968
rect 29288 14550 29316 15302
rect 29368 15020 29420 15026
rect 29368 14962 29420 14968
rect 29460 15020 29512 15026
rect 29460 14962 29512 14968
rect 29552 15020 29604 15026
rect 29552 14962 29604 14968
rect 29380 14890 29408 14962
rect 29368 14884 29420 14890
rect 29368 14826 29420 14832
rect 29276 14544 29328 14550
rect 29276 14486 29328 14492
rect 29276 14408 29328 14414
rect 29276 14350 29328 14356
rect 29288 13530 29316 14350
rect 29276 13524 29328 13530
rect 29276 13466 29328 13472
rect 29380 12434 29408 14826
rect 29472 14414 29500 14962
rect 29460 14408 29512 14414
rect 29460 14350 29512 14356
rect 29564 13938 29592 14962
rect 29552 13932 29604 13938
rect 29552 13874 29604 13880
rect 29012 12406 29132 12434
rect 29288 12406 29408 12434
rect 29460 12436 29512 12442
rect 28724 11756 28776 11762
rect 28724 11698 28776 11704
rect 28632 11212 28684 11218
rect 28632 11154 28684 11160
rect 28644 10266 28672 11154
rect 29012 10810 29040 12406
rect 29092 11756 29144 11762
rect 29092 11698 29144 11704
rect 29104 11354 29132 11698
rect 29092 11348 29144 11354
rect 29092 11290 29144 11296
rect 29000 10804 29052 10810
rect 29000 10746 29052 10752
rect 29092 10736 29144 10742
rect 29092 10678 29144 10684
rect 29000 10668 29052 10674
rect 29000 10610 29052 10616
rect 28722 10432 28778 10441
rect 28722 10367 28778 10376
rect 28632 10260 28684 10266
rect 28632 10202 28684 10208
rect 28540 9920 28592 9926
rect 28540 9862 28592 9868
rect 28446 9208 28502 9217
rect 28446 9143 28502 9152
rect 28736 9110 28764 10367
rect 28814 10160 28870 10169
rect 28814 10095 28870 10104
rect 28828 10062 28856 10095
rect 29012 10062 29040 10610
rect 29104 10266 29132 10678
rect 29288 10674 29316 12406
rect 29460 12378 29512 12384
rect 29276 10668 29328 10674
rect 29276 10610 29328 10616
rect 29184 10464 29236 10470
rect 29184 10406 29236 10412
rect 29092 10260 29144 10266
rect 29092 10202 29144 10208
rect 29196 10062 29224 10406
rect 28816 10056 28868 10062
rect 28816 9998 28868 10004
rect 29000 10056 29052 10062
rect 29000 9998 29052 10004
rect 29184 10056 29236 10062
rect 29184 9998 29236 10004
rect 29276 10056 29328 10062
rect 29276 9998 29328 10004
rect 28908 9988 28960 9994
rect 28908 9930 28960 9936
rect 28920 9654 28948 9930
rect 28908 9648 28960 9654
rect 28908 9590 28960 9596
rect 29288 9178 29316 9998
rect 29276 9172 29328 9178
rect 29276 9114 29328 9120
rect 28724 9104 28776 9110
rect 28724 9046 28776 9052
rect 28172 8900 28224 8906
rect 28172 8842 28224 8848
rect 28184 8634 28212 8842
rect 28356 8832 28408 8838
rect 28356 8774 28408 8780
rect 28080 8628 28132 8634
rect 28080 8570 28132 8576
rect 28172 8628 28224 8634
rect 28172 8570 28224 8576
rect 27436 8560 27488 8566
rect 27436 8502 27488 8508
rect 27804 8560 27856 8566
rect 27804 8502 27856 8508
rect 27448 8090 27476 8502
rect 28368 8362 28396 8774
rect 28356 8356 28408 8362
rect 28356 8298 28408 8304
rect 27436 8084 27488 8090
rect 27436 8026 27488 8032
rect 28368 7886 28396 8298
rect 28736 8090 28764 9046
rect 28724 8084 28776 8090
rect 28724 8026 28776 8032
rect 27252 7880 27304 7886
rect 27252 7822 27304 7828
rect 28356 7880 28408 7886
rect 28356 7822 28408 7828
rect 27160 7744 27212 7750
rect 27160 7686 27212 7692
rect 28724 7404 28776 7410
rect 28724 7346 28776 7352
rect 28736 6934 28764 7346
rect 29368 7200 29420 7206
rect 29368 7142 29420 7148
rect 27804 6928 27856 6934
rect 27804 6870 27856 6876
rect 28724 6928 28776 6934
rect 28724 6870 28776 6876
rect 26884 6656 26936 6662
rect 26884 6598 26936 6604
rect 27344 6656 27396 6662
rect 27344 6598 27396 6604
rect 26148 6452 26200 6458
rect 26148 6394 26200 6400
rect 26240 6452 26292 6458
rect 26240 6394 26292 6400
rect 26252 6118 26280 6394
rect 26240 6112 26292 6118
rect 26240 6054 26292 6060
rect 27356 5778 27384 6598
rect 27816 6186 27844 6870
rect 27896 6860 27948 6866
rect 27896 6802 27948 6808
rect 28816 6860 28868 6866
rect 28816 6802 28868 6808
rect 27908 6662 27936 6802
rect 27896 6656 27948 6662
rect 27896 6598 27948 6604
rect 28828 6458 28856 6802
rect 29000 6792 29052 6798
rect 29000 6734 29052 6740
rect 28816 6452 28868 6458
rect 28816 6394 28868 6400
rect 29012 6322 29040 6734
rect 29092 6384 29144 6390
rect 29092 6326 29144 6332
rect 28816 6316 28868 6322
rect 28816 6258 28868 6264
rect 29000 6316 29052 6322
rect 29000 6258 29052 6264
rect 27804 6180 27856 6186
rect 27804 6122 27856 6128
rect 27436 6112 27488 6118
rect 27436 6054 27488 6060
rect 27344 5772 27396 5778
rect 27344 5714 27396 5720
rect 27448 5642 27476 6054
rect 28828 5914 28856 6258
rect 29104 5914 29132 6326
rect 29380 6254 29408 7142
rect 29472 6458 29500 12378
rect 29656 12374 29684 17614
rect 29828 17128 29880 17134
rect 29828 17070 29880 17076
rect 29736 16788 29788 16794
rect 29736 16730 29788 16736
rect 29748 15162 29776 16730
rect 29736 15156 29788 15162
rect 29736 15098 29788 15104
rect 29736 13864 29788 13870
rect 29736 13806 29788 13812
rect 29644 12368 29696 12374
rect 29644 12310 29696 12316
rect 29748 12306 29776 13806
rect 29840 12442 29868 17070
rect 29932 15094 29960 19450
rect 30116 18630 30144 22578
rect 30392 22030 30420 26930
rect 31128 26382 31156 30688
rect 31208 30670 31260 30676
rect 32772 29640 32824 29646
rect 32772 29582 32824 29588
rect 32784 29238 32812 29582
rect 32772 29232 32824 29238
rect 32772 29174 32824 29180
rect 31852 27600 31904 27606
rect 31852 27542 31904 27548
rect 31760 27532 31812 27538
rect 31760 27474 31812 27480
rect 31484 27464 31536 27470
rect 31536 27424 31616 27452
rect 31484 27406 31536 27412
rect 31116 26376 31168 26382
rect 31116 26318 31168 26324
rect 30472 26308 30524 26314
rect 30472 26250 30524 26256
rect 30484 26042 30512 26250
rect 30472 26036 30524 26042
rect 30472 25978 30524 25984
rect 30748 26036 30800 26042
rect 30748 25978 30800 25984
rect 30656 25832 30708 25838
rect 30656 25774 30708 25780
rect 30668 25498 30696 25774
rect 30656 25492 30708 25498
rect 30656 25434 30708 25440
rect 30564 25356 30616 25362
rect 30564 25298 30616 25304
rect 30576 24410 30604 25298
rect 30760 25294 30788 25978
rect 31024 25696 31076 25702
rect 31024 25638 31076 25644
rect 30932 25492 30984 25498
rect 30932 25434 30984 25440
rect 30748 25288 30800 25294
rect 30748 25230 30800 25236
rect 30840 25152 30892 25158
rect 30840 25094 30892 25100
rect 30852 24818 30880 25094
rect 30840 24812 30892 24818
rect 30840 24754 30892 24760
rect 30564 24404 30616 24410
rect 30564 24346 30616 24352
rect 30656 24132 30708 24138
rect 30656 24074 30708 24080
rect 30668 23866 30696 24074
rect 30944 23866 30972 25434
rect 31036 25294 31064 25638
rect 31024 25288 31076 25294
rect 31024 25230 31076 25236
rect 31036 24562 31064 25230
rect 31128 24750 31156 26318
rect 31484 26240 31536 26246
rect 31484 26182 31536 26188
rect 31496 26042 31524 26182
rect 31484 26036 31536 26042
rect 31484 25978 31536 25984
rect 31300 25424 31352 25430
rect 31300 25366 31352 25372
rect 31312 25158 31340 25366
rect 31300 25152 31352 25158
rect 31300 25094 31352 25100
rect 31116 24744 31168 24750
rect 31116 24686 31168 24692
rect 31036 24534 31156 24562
rect 30656 23860 30708 23866
rect 30656 23802 30708 23808
rect 30932 23860 30984 23866
rect 30932 23802 30984 23808
rect 30656 23724 30708 23730
rect 30656 23666 30708 23672
rect 30564 22636 30616 22642
rect 30564 22578 30616 22584
rect 30576 22234 30604 22578
rect 30564 22228 30616 22234
rect 30564 22170 30616 22176
rect 30380 22024 30432 22030
rect 30380 21966 30432 21972
rect 30288 21412 30340 21418
rect 30288 21354 30340 21360
rect 30300 21146 30328 21354
rect 30288 21140 30340 21146
rect 30288 21082 30340 21088
rect 30300 20466 30328 21082
rect 30288 20460 30340 20466
rect 30288 20402 30340 20408
rect 30380 20256 30432 20262
rect 30380 20198 30432 20204
rect 30392 19922 30420 20198
rect 30380 19916 30432 19922
rect 30380 19858 30432 19864
rect 30472 19712 30524 19718
rect 30472 19654 30524 19660
rect 30484 19310 30512 19654
rect 30472 19304 30524 19310
rect 30472 19246 30524 19252
rect 30196 18964 30248 18970
rect 30196 18906 30248 18912
rect 30012 18624 30064 18630
rect 30012 18566 30064 18572
rect 30104 18624 30156 18630
rect 30104 18566 30156 18572
rect 30024 18290 30052 18566
rect 30012 18284 30064 18290
rect 30012 18226 30064 18232
rect 30024 17746 30052 18226
rect 30104 18216 30156 18222
rect 30104 18158 30156 18164
rect 30012 17740 30064 17746
rect 30012 17682 30064 17688
rect 30116 17338 30144 18158
rect 30208 17678 30236 18906
rect 30380 18896 30432 18902
rect 30380 18838 30432 18844
rect 30288 18624 30340 18630
rect 30288 18566 30340 18572
rect 30196 17672 30248 17678
rect 30196 17614 30248 17620
rect 30104 17332 30156 17338
rect 30104 17274 30156 17280
rect 30196 16788 30248 16794
rect 30196 16730 30248 16736
rect 30012 16584 30064 16590
rect 30010 16552 30012 16561
rect 30064 16552 30066 16561
rect 30010 16487 30066 16496
rect 30024 15162 30052 16487
rect 30208 15706 30236 16730
rect 30196 15700 30248 15706
rect 30196 15642 30248 15648
rect 30012 15156 30064 15162
rect 30012 15098 30064 15104
rect 29920 15088 29972 15094
rect 29920 15030 29972 15036
rect 30024 14822 30052 15098
rect 30208 15026 30236 15642
rect 30196 15020 30248 15026
rect 30196 14962 30248 14968
rect 30012 14816 30064 14822
rect 30012 14758 30064 14764
rect 30300 14482 30328 18566
rect 30392 16810 30420 18838
rect 30484 18766 30512 19246
rect 30564 19236 30616 19242
rect 30564 19178 30616 19184
rect 30472 18760 30524 18766
rect 30472 18702 30524 18708
rect 30576 18154 30604 19178
rect 30564 18148 30616 18154
rect 30564 18090 30616 18096
rect 30392 16782 30512 16810
rect 30380 16584 30432 16590
rect 30380 16526 30432 16532
rect 30392 16046 30420 16526
rect 30380 16040 30432 16046
rect 30380 15982 30432 15988
rect 30392 15502 30420 15982
rect 30380 15496 30432 15502
rect 30380 15438 30432 15444
rect 30380 15360 30432 15366
rect 30380 15302 30432 15308
rect 30288 14476 30340 14482
rect 30288 14418 30340 14424
rect 30012 14272 30064 14278
rect 30012 14214 30064 14220
rect 30024 13938 30052 14214
rect 30012 13932 30064 13938
rect 30012 13874 30064 13880
rect 29828 12436 29880 12442
rect 29828 12378 29880 12384
rect 29736 12300 29788 12306
rect 29736 12242 29788 12248
rect 30104 12164 30156 12170
rect 30104 12106 30156 12112
rect 30116 11898 30144 12106
rect 30104 11892 30156 11898
rect 30104 11834 30156 11840
rect 30288 11756 30340 11762
rect 30288 11698 30340 11704
rect 29828 11688 29880 11694
rect 29828 11630 29880 11636
rect 29552 11552 29604 11558
rect 29552 11494 29604 11500
rect 29564 11150 29592 11494
rect 29552 11144 29604 11150
rect 29552 11086 29604 11092
rect 29644 11144 29696 11150
rect 29644 11086 29696 11092
rect 29564 10713 29592 11086
rect 29656 10810 29684 11086
rect 29644 10804 29696 10810
rect 29644 10746 29696 10752
rect 29550 10704 29606 10713
rect 29550 10639 29606 10648
rect 29840 10606 29868 11630
rect 30196 11144 30248 11150
rect 30196 11086 30248 11092
rect 30208 10742 30236 11086
rect 30300 10810 30328 11698
rect 30288 10804 30340 10810
rect 30288 10746 30340 10752
rect 30196 10736 30248 10742
rect 30196 10678 30248 10684
rect 29828 10600 29880 10606
rect 29828 10542 29880 10548
rect 29840 10266 29868 10542
rect 29828 10260 29880 10266
rect 29828 10202 29880 10208
rect 29642 10160 29698 10169
rect 29642 10095 29698 10104
rect 29656 10062 29684 10095
rect 29840 10062 29868 10202
rect 29644 10056 29696 10062
rect 29644 9998 29696 10004
rect 29828 10056 29880 10062
rect 29828 9998 29880 10004
rect 29656 8430 29684 9998
rect 29736 9920 29788 9926
rect 29736 9862 29788 9868
rect 29748 8945 29776 9862
rect 29840 9586 29868 9998
rect 29828 9580 29880 9586
rect 29828 9522 29880 9528
rect 30300 9518 30328 10746
rect 30288 9512 30340 9518
rect 30288 9454 30340 9460
rect 29734 8936 29790 8945
rect 29734 8871 29790 8880
rect 30392 8498 30420 15302
rect 30484 15094 30512 16782
rect 30668 16402 30696 23666
rect 30932 23656 30984 23662
rect 30932 23598 30984 23604
rect 30748 23180 30800 23186
rect 30748 23122 30800 23128
rect 30760 22001 30788 23122
rect 30746 21992 30802 22001
rect 30746 21927 30802 21936
rect 30760 21350 30788 21927
rect 30944 21418 30972 23598
rect 31024 22092 31076 22098
rect 31024 22034 31076 22040
rect 31036 22001 31064 22034
rect 31022 21992 31078 22001
rect 31022 21927 31078 21936
rect 31024 21888 31076 21894
rect 31024 21830 31076 21836
rect 31036 21457 31064 21830
rect 31022 21448 31078 21457
rect 30932 21412 30984 21418
rect 31022 21383 31078 21392
rect 30932 21354 30984 21360
rect 30748 21344 30800 21350
rect 30746 21312 30748 21321
rect 30800 21312 30802 21321
rect 30746 21247 30802 21256
rect 31128 21185 31156 24534
rect 31312 23730 31340 25094
rect 31392 24608 31444 24614
rect 31392 24550 31444 24556
rect 31484 24608 31536 24614
rect 31484 24550 31536 24556
rect 31404 23730 31432 24550
rect 31300 23724 31352 23730
rect 31300 23666 31352 23672
rect 31392 23724 31444 23730
rect 31392 23666 31444 23672
rect 31392 22636 31444 22642
rect 31392 22578 31444 22584
rect 31404 22030 31432 22578
rect 31392 22024 31444 22030
rect 31392 21966 31444 21972
rect 31208 21412 31260 21418
rect 31208 21354 31260 21360
rect 30838 21176 30894 21185
rect 30838 21111 30894 21120
rect 31114 21176 31170 21185
rect 31220 21146 31248 21354
rect 31114 21111 31170 21120
rect 31208 21140 31260 21146
rect 30748 18760 30800 18766
rect 30748 18702 30800 18708
rect 30760 16590 30788 18702
rect 30852 16794 30880 21111
rect 31208 21082 31260 21088
rect 31116 20868 31168 20874
rect 31116 20810 31168 20816
rect 31024 19168 31076 19174
rect 31024 19110 31076 19116
rect 31036 18834 31064 19110
rect 31024 18828 31076 18834
rect 31024 18770 31076 18776
rect 30932 18352 30984 18358
rect 30932 18294 30984 18300
rect 30944 17678 30972 18294
rect 30932 17672 30984 17678
rect 30932 17614 30984 17620
rect 30944 17338 30972 17614
rect 31024 17536 31076 17542
rect 31024 17478 31076 17484
rect 30932 17332 30984 17338
rect 30932 17274 30984 17280
rect 30840 16788 30892 16794
rect 30840 16730 30892 16736
rect 30748 16584 30800 16590
rect 30748 16526 30800 16532
rect 30932 16516 30984 16522
rect 30932 16458 30984 16464
rect 30668 16374 30788 16402
rect 30564 16040 30616 16046
rect 30564 15982 30616 15988
rect 30576 15366 30604 15982
rect 30656 15904 30708 15910
rect 30656 15846 30708 15852
rect 30668 15502 30696 15846
rect 30656 15496 30708 15502
rect 30656 15438 30708 15444
rect 30564 15360 30616 15366
rect 30564 15302 30616 15308
rect 30562 15192 30618 15201
rect 30562 15127 30564 15136
rect 30616 15127 30618 15136
rect 30564 15098 30616 15104
rect 30472 15088 30524 15094
rect 30472 15030 30524 15036
rect 30564 14476 30616 14482
rect 30564 14418 30616 14424
rect 30576 13462 30604 14418
rect 30564 13456 30616 13462
rect 30564 13398 30616 13404
rect 30656 11688 30708 11694
rect 30656 11630 30708 11636
rect 30668 11354 30696 11630
rect 30656 11348 30708 11354
rect 30656 11290 30708 11296
rect 30760 11218 30788 16374
rect 30840 16108 30892 16114
rect 30840 16050 30892 16056
rect 30852 15434 30880 16050
rect 30840 15428 30892 15434
rect 30840 15370 30892 15376
rect 30852 14550 30880 15370
rect 30944 15162 30972 16458
rect 30932 15156 30984 15162
rect 30932 15098 30984 15104
rect 31036 15094 31064 17478
rect 31128 16046 31156 20810
rect 31496 20346 31524 24550
rect 31588 20874 31616 27424
rect 31772 27062 31800 27474
rect 31760 27056 31812 27062
rect 31760 26998 31812 27004
rect 31864 26382 31892 27542
rect 32784 27538 32812 29174
rect 32772 27532 32824 27538
rect 32772 27474 32824 27480
rect 31852 26376 31904 26382
rect 31852 26318 31904 26324
rect 32784 25838 32812 27474
rect 32772 25832 32824 25838
rect 32772 25774 32824 25780
rect 31760 24812 31812 24818
rect 31760 24754 31812 24760
rect 31772 24410 31800 24754
rect 31760 24404 31812 24410
rect 31760 24346 31812 24352
rect 31772 23866 31800 24346
rect 32784 24206 32812 25774
rect 32772 24200 32824 24206
rect 32772 24142 32824 24148
rect 31760 23860 31812 23866
rect 31760 23802 31812 23808
rect 31576 20868 31628 20874
rect 31576 20810 31628 20816
rect 32220 20528 32272 20534
rect 32220 20470 32272 20476
rect 31404 20318 31524 20346
rect 31404 20262 31432 20318
rect 31392 20256 31444 20262
rect 31392 20198 31444 20204
rect 31208 19508 31260 19514
rect 31208 19450 31260 19456
rect 31220 17814 31248 19450
rect 31300 18080 31352 18086
rect 31300 18022 31352 18028
rect 31208 17808 31260 17814
rect 31208 17750 31260 17756
rect 31312 17610 31340 18022
rect 31300 17604 31352 17610
rect 31300 17546 31352 17552
rect 31300 17332 31352 17338
rect 31300 17274 31352 17280
rect 31208 16176 31260 16182
rect 31208 16118 31260 16124
rect 31116 16040 31168 16046
rect 31116 15982 31168 15988
rect 31220 15434 31248 16118
rect 31208 15428 31260 15434
rect 31208 15370 31260 15376
rect 31024 15088 31076 15094
rect 31024 15030 31076 15036
rect 30840 14544 30892 14550
rect 30840 14486 30892 14492
rect 31116 14408 31168 14414
rect 31116 14350 31168 14356
rect 31128 14074 31156 14350
rect 31116 14068 31168 14074
rect 31116 14010 31168 14016
rect 30932 12096 30984 12102
rect 30932 12038 30984 12044
rect 30944 11762 30972 12038
rect 30932 11756 30984 11762
rect 30932 11698 30984 11704
rect 30748 11212 30800 11218
rect 30748 11154 30800 11160
rect 30470 10024 30526 10033
rect 31220 9994 31248 15370
rect 31312 11762 31340 17274
rect 31404 16538 31432 20198
rect 32036 20052 32088 20058
rect 32036 19994 32088 20000
rect 32048 19786 32076 19994
rect 32232 19786 32260 20470
rect 32496 19848 32548 19854
rect 32496 19790 32548 19796
rect 32036 19780 32088 19786
rect 32036 19722 32088 19728
rect 32220 19780 32272 19786
rect 32220 19722 32272 19728
rect 31760 18624 31812 18630
rect 31760 18566 31812 18572
rect 31772 18358 31800 18566
rect 31760 18352 31812 18358
rect 31760 18294 31812 18300
rect 31668 18284 31720 18290
rect 31668 18226 31720 18232
rect 31576 18148 31628 18154
rect 31576 18090 31628 18096
rect 31588 17678 31616 18090
rect 31576 17672 31628 17678
rect 31576 17614 31628 17620
rect 31484 17536 31536 17542
rect 31484 17478 31536 17484
rect 31496 16658 31524 17478
rect 31484 16652 31536 16658
rect 31484 16594 31536 16600
rect 31404 16510 31524 16538
rect 31392 16108 31444 16114
rect 31392 16050 31444 16056
rect 31404 15706 31432 16050
rect 31496 15910 31524 16510
rect 31680 16454 31708 18226
rect 32048 16574 32076 19722
rect 32128 19372 32180 19378
rect 32128 19314 32180 19320
rect 32140 18426 32168 19314
rect 32232 18834 32260 19722
rect 32508 18970 32536 19790
rect 32876 19310 32904 33798
rect 33508 33516 33560 33522
rect 33508 33458 33560 33464
rect 33416 33380 33468 33386
rect 33416 33322 33468 33328
rect 33140 33312 33192 33318
rect 33140 33254 33192 33260
rect 33152 32842 33180 33254
rect 33428 32978 33456 33322
rect 33416 32972 33468 32978
rect 33416 32914 33468 32920
rect 33520 32842 33548 33458
rect 34072 33318 34100 33934
rect 34336 33924 34388 33930
rect 34336 33866 34388 33872
rect 34348 33561 34376 33866
rect 34428 33856 34480 33862
rect 34428 33798 34480 33804
rect 34334 33552 34390 33561
rect 34152 33516 34204 33522
rect 34440 33522 34468 33798
rect 34532 33658 34560 35634
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34520 33652 34572 33658
rect 34520 33594 34572 33600
rect 34334 33487 34390 33496
rect 34428 33516 34480 33522
rect 34152 33458 34204 33464
rect 34428 33458 34480 33464
rect 34060 33312 34112 33318
rect 34060 33254 34112 33260
rect 33140 32836 33192 32842
rect 33140 32778 33192 32784
rect 33508 32836 33560 32842
rect 33508 32778 33560 32784
rect 33520 31754 33548 32778
rect 34164 32570 34192 33458
rect 34440 32774 34468 33458
rect 34532 33114 34560 33594
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34520 33108 34572 33114
rect 34520 33050 34572 33056
rect 34428 32768 34480 32774
rect 34428 32710 34480 32716
rect 34152 32564 34204 32570
rect 34152 32506 34204 32512
rect 33784 31884 33836 31890
rect 33784 31826 33836 31832
rect 33508 31748 33560 31754
rect 33508 31690 33560 31696
rect 33048 30660 33100 30666
rect 33048 30602 33100 30608
rect 33060 30258 33088 30602
rect 33048 30252 33100 30258
rect 33048 30194 33100 30200
rect 33520 30122 33548 31690
rect 33796 31482 33824 31826
rect 33784 31476 33836 31482
rect 33784 31418 33836 31424
rect 34440 31346 34468 32710
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34520 31680 34572 31686
rect 34520 31622 34572 31628
rect 34794 31648 34850 31657
rect 34532 31346 34560 31622
rect 34794 31583 34850 31592
rect 34808 31414 34836 31583
rect 34796 31408 34848 31414
rect 34796 31350 34848 31356
rect 34428 31340 34480 31346
rect 34428 31282 34480 31288
rect 34520 31340 34572 31346
rect 34520 31282 34572 31288
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34152 30728 34204 30734
rect 34152 30670 34204 30676
rect 34164 30326 34192 30670
rect 34520 30660 34572 30666
rect 34520 30602 34572 30608
rect 34152 30320 34204 30326
rect 34152 30262 34204 30268
rect 33508 30116 33560 30122
rect 33508 30058 33560 30064
rect 33416 30048 33468 30054
rect 33416 29990 33468 29996
rect 33324 27396 33376 27402
rect 33324 27338 33376 27344
rect 33336 27130 33364 27338
rect 33324 27124 33376 27130
rect 33324 27066 33376 27072
rect 33048 24132 33100 24138
rect 33048 24074 33100 24080
rect 33060 23866 33088 24074
rect 33048 23860 33100 23866
rect 33048 23802 33100 23808
rect 33048 22432 33100 22438
rect 33048 22374 33100 22380
rect 33060 22234 33088 22374
rect 33048 22228 33100 22234
rect 33048 22170 33100 22176
rect 33140 22092 33192 22098
rect 33140 22034 33192 22040
rect 33152 20466 33180 22034
rect 33140 20460 33192 20466
rect 33140 20402 33192 20408
rect 33428 20058 33456 29990
rect 33520 29578 33548 30058
rect 33600 30048 33652 30054
rect 33600 29990 33652 29996
rect 33612 29714 33640 29990
rect 34164 29850 34192 30262
rect 34244 30252 34296 30258
rect 34244 30194 34296 30200
rect 34152 29844 34204 29850
rect 34152 29786 34204 29792
rect 33600 29708 33652 29714
rect 33600 29650 33652 29656
rect 33508 29572 33560 29578
rect 33508 29514 33560 29520
rect 34060 27396 34112 27402
rect 34060 27338 34112 27344
rect 33968 26988 34020 26994
rect 33968 26930 34020 26936
rect 33980 26586 34008 26930
rect 33968 26580 34020 26586
rect 33968 26522 34020 26528
rect 33784 26240 33836 26246
rect 34072 26234 34100 27338
rect 34256 26994 34284 30194
rect 34532 29753 34560 30602
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34518 29744 34574 29753
rect 34518 29679 34574 29688
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34520 28076 34572 28082
rect 34520 28018 34572 28024
rect 34532 27674 34560 28018
rect 35348 28008 35400 28014
rect 35348 27950 35400 27956
rect 35360 27849 35388 27950
rect 35346 27840 35402 27849
rect 34934 27772 35242 27781
rect 35346 27775 35402 27784
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34520 27668 34572 27674
rect 34520 27610 34572 27616
rect 34532 27130 34560 27610
rect 34520 27124 34572 27130
rect 34520 27066 34572 27072
rect 34244 26988 34296 26994
rect 34244 26930 34296 26936
rect 34520 26988 34572 26994
rect 34520 26930 34572 26936
rect 34256 26382 34284 26930
rect 34244 26376 34296 26382
rect 34244 26318 34296 26324
rect 33784 26182 33836 26188
rect 33980 26206 34100 26234
rect 33600 26036 33652 26042
rect 33600 25978 33652 25984
rect 33612 25922 33640 25978
rect 33796 25974 33824 26182
rect 33980 25974 34008 26206
rect 33520 25894 33640 25922
rect 33784 25968 33836 25974
rect 33784 25910 33836 25916
rect 33968 25968 34020 25974
rect 33968 25910 34020 25916
rect 33520 24138 33548 25894
rect 33508 24132 33560 24138
rect 33508 24074 33560 24080
rect 33520 21962 33548 24074
rect 34256 23730 34284 26318
rect 34532 26314 34560 26930
rect 34796 26920 34848 26926
rect 34796 26862 34848 26868
rect 34520 26308 34572 26314
rect 34520 26250 34572 26256
rect 34808 25945 34836 26862
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34980 26308 35032 26314
rect 34980 26250 35032 26256
rect 34992 26042 35020 26250
rect 34980 26036 35032 26042
rect 34980 25978 35032 25984
rect 34794 25936 34850 25945
rect 34794 25871 34850 25880
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34520 24064 34572 24070
rect 34520 24006 34572 24012
rect 34794 24032 34850 24041
rect 34532 23730 34560 24006
rect 34794 23967 34850 23976
rect 34808 23798 34836 23967
rect 34796 23792 34848 23798
rect 34796 23734 34848 23740
rect 34244 23724 34296 23730
rect 34244 23666 34296 23672
rect 34520 23724 34572 23730
rect 34520 23666 34572 23672
rect 34256 22642 34284 23666
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34244 22636 34296 22642
rect 34244 22578 34296 22584
rect 34520 22636 34572 22642
rect 34520 22578 34572 22584
rect 33508 21956 33560 21962
rect 33508 21898 33560 21904
rect 33520 20534 33548 21898
rect 33508 20528 33560 20534
rect 33508 20470 33560 20476
rect 33968 20392 34020 20398
rect 33968 20334 34020 20340
rect 33980 20058 34008 20334
rect 33416 20052 33468 20058
rect 33416 19994 33468 20000
rect 33968 20052 34020 20058
rect 33968 19994 34020 20000
rect 34256 19854 34284 22578
rect 34532 22234 34560 22578
rect 34796 22568 34848 22574
rect 34796 22510 34848 22516
rect 34520 22228 34572 22234
rect 34520 22170 34572 22176
rect 34808 22137 34836 22510
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34794 22128 34850 22137
rect 34794 22063 34850 22072
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34704 20936 34756 20942
rect 34704 20878 34756 20884
rect 34716 20262 34744 20878
rect 35348 20868 35400 20874
rect 35348 20810 35400 20816
rect 34704 20256 34756 20262
rect 35360 20233 35388 20810
rect 34704 20198 34756 20204
rect 35346 20224 35402 20233
rect 34244 19848 34296 19854
rect 34244 19790 34296 19796
rect 34716 19786 34744 20198
rect 34934 20156 35242 20165
rect 35346 20159 35402 20168
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34704 19780 34756 19786
rect 34704 19722 34756 19728
rect 34888 19780 34940 19786
rect 34888 19722 34940 19728
rect 34900 19310 34928 19722
rect 32864 19304 32916 19310
rect 32864 19246 32916 19252
rect 34888 19304 34940 19310
rect 34888 19246 34940 19252
rect 32772 19168 32824 19174
rect 32772 19110 32824 19116
rect 32496 18964 32548 18970
rect 32496 18906 32548 18912
rect 32220 18828 32272 18834
rect 32220 18770 32272 18776
rect 32588 18828 32640 18834
rect 32588 18770 32640 18776
rect 32128 18420 32180 18426
rect 32128 18362 32180 18368
rect 32128 17672 32180 17678
rect 32128 17614 32180 17620
rect 31772 16546 32076 16574
rect 31668 16448 31720 16454
rect 31668 16390 31720 16396
rect 31484 15904 31536 15910
rect 31484 15846 31536 15852
rect 31392 15700 31444 15706
rect 31392 15642 31444 15648
rect 31496 15366 31524 15846
rect 31484 15360 31536 15366
rect 31484 15302 31536 15308
rect 31496 14822 31524 15302
rect 31484 14816 31536 14822
rect 31484 14758 31536 14764
rect 31392 12232 31444 12238
rect 31392 12174 31444 12180
rect 31404 11898 31432 12174
rect 31496 11898 31524 14758
rect 31392 11892 31444 11898
rect 31392 11834 31444 11840
rect 31484 11892 31536 11898
rect 31484 11834 31536 11840
rect 31300 11756 31352 11762
rect 31300 11698 31352 11704
rect 31312 10826 31340 11698
rect 31312 10798 31432 10826
rect 30470 9959 30526 9968
rect 31208 9988 31260 9994
rect 30484 9926 30512 9959
rect 31208 9930 31260 9936
rect 30472 9920 30524 9926
rect 30472 9862 30524 9868
rect 30484 9518 30512 9862
rect 31220 9722 31248 9930
rect 31208 9716 31260 9722
rect 31208 9658 31260 9664
rect 30472 9512 30524 9518
rect 30472 9454 30524 9460
rect 30380 8492 30432 8498
rect 30380 8434 30432 8440
rect 29644 8424 29696 8430
rect 29644 8366 29696 8372
rect 31116 8424 31168 8430
rect 31116 8366 31168 8372
rect 29828 8288 29880 8294
rect 29828 8230 29880 8236
rect 29840 7818 29868 8230
rect 31128 7954 31156 8366
rect 29920 7948 29972 7954
rect 29920 7890 29972 7896
rect 31024 7948 31076 7954
rect 31024 7890 31076 7896
rect 31116 7948 31168 7954
rect 31116 7890 31168 7896
rect 29828 7812 29880 7818
rect 29828 7754 29880 7760
rect 29932 6798 29960 7890
rect 30472 7404 30524 7410
rect 30472 7346 30524 7352
rect 30196 6860 30248 6866
rect 30196 6802 30248 6808
rect 29920 6792 29972 6798
rect 29920 6734 29972 6740
rect 29460 6452 29512 6458
rect 29460 6394 29512 6400
rect 29932 6254 29960 6734
rect 30012 6316 30064 6322
rect 30012 6258 30064 6264
rect 29368 6248 29420 6254
rect 29736 6248 29788 6254
rect 29368 6190 29420 6196
rect 29642 6216 29698 6225
rect 29736 6190 29788 6196
rect 29920 6248 29972 6254
rect 29920 6190 29972 6196
rect 29642 6151 29698 6160
rect 28816 5908 28868 5914
rect 28816 5850 28868 5856
rect 29092 5908 29144 5914
rect 29092 5850 29144 5856
rect 29656 5710 29684 6151
rect 29644 5704 29696 5710
rect 29644 5646 29696 5652
rect 27436 5636 27488 5642
rect 27436 5578 27488 5584
rect 28724 5636 28776 5642
rect 28724 5578 28776 5584
rect 24860 5296 24912 5302
rect 24860 5238 24912 5244
rect 26056 5296 26108 5302
rect 26056 5238 26108 5244
rect 24400 4548 24452 4554
rect 24400 4490 24452 4496
rect 23572 4480 23624 4486
rect 23572 4422 23624 4428
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 28736 4078 28764 5578
rect 29000 4684 29052 4690
rect 29000 4626 29052 4632
rect 29012 4146 29040 4626
rect 29092 4548 29144 4554
rect 29092 4490 29144 4496
rect 29104 4146 29132 4490
rect 29748 4434 29776 6190
rect 29828 6180 29880 6186
rect 29828 6122 29880 6128
rect 29840 5642 29868 6122
rect 29828 5636 29880 5642
rect 29828 5578 29880 5584
rect 29932 4554 29960 6190
rect 30024 5642 30052 6258
rect 30208 5710 30236 6802
rect 30484 6254 30512 7346
rect 30840 6656 30892 6662
rect 30840 6598 30892 6604
rect 30748 6316 30800 6322
rect 30748 6258 30800 6264
rect 30472 6248 30524 6254
rect 30472 6190 30524 6196
rect 30288 5840 30340 5846
rect 30288 5782 30340 5788
rect 30196 5704 30248 5710
rect 30196 5646 30248 5652
rect 30012 5636 30064 5642
rect 30012 5578 30064 5584
rect 30208 5574 30236 5646
rect 30196 5568 30248 5574
rect 30196 5510 30248 5516
rect 30300 4690 30328 5782
rect 30380 5704 30432 5710
rect 30380 5646 30432 5652
rect 30392 5370 30420 5646
rect 30380 5364 30432 5370
rect 30380 5306 30432 5312
rect 30484 5234 30512 6190
rect 30656 5840 30708 5846
rect 30656 5782 30708 5788
rect 30668 5710 30696 5782
rect 30760 5778 30788 6258
rect 30852 5817 30880 6598
rect 31036 5896 31064 7890
rect 31128 7206 31156 7890
rect 31116 7200 31168 7206
rect 31116 7142 31168 7148
rect 31116 6792 31168 6798
rect 31116 6734 31168 6740
rect 31128 6322 31156 6734
rect 31220 6458 31248 9658
rect 31300 8492 31352 8498
rect 31300 8434 31352 8440
rect 31312 8090 31340 8434
rect 31404 8242 31432 10798
rect 31772 9081 31800 16546
rect 32140 16046 32168 17614
rect 32600 16454 32628 18770
rect 32784 18766 32812 19110
rect 32772 18760 32824 18766
rect 32772 18702 32824 18708
rect 32784 18426 32812 18702
rect 32772 18420 32824 18426
rect 32772 18362 32824 18368
rect 32680 18080 32732 18086
rect 32680 18022 32732 18028
rect 32692 17678 32720 18022
rect 32680 17672 32732 17678
rect 32680 17614 32732 17620
rect 32876 16590 32904 19246
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34152 18760 34204 18766
rect 34150 18728 34152 18737
rect 34204 18728 34206 18737
rect 34150 18663 34206 18672
rect 33692 18624 33744 18630
rect 33692 18566 33744 18572
rect 33784 18624 33836 18630
rect 33784 18566 33836 18572
rect 34520 18624 34572 18630
rect 34520 18566 34572 18572
rect 33704 18358 33732 18566
rect 33140 18352 33192 18358
rect 33140 18294 33192 18300
rect 33692 18352 33744 18358
rect 33692 18294 33744 18300
rect 33152 17610 33180 18294
rect 33796 17746 33824 18566
rect 34532 18290 34560 18566
rect 34794 18320 34850 18329
rect 34520 18284 34572 18290
rect 34794 18255 34796 18264
rect 34520 18226 34572 18232
rect 34848 18255 34850 18264
rect 34796 18226 34848 18232
rect 34532 17882 34560 18226
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34520 17876 34572 17882
rect 34520 17818 34572 17824
rect 33784 17740 33836 17746
rect 33784 17682 33836 17688
rect 33140 17604 33192 17610
rect 33140 17546 33192 17552
rect 32864 16584 32916 16590
rect 32916 16546 32996 16574
rect 32864 16526 32916 16532
rect 32968 16454 32996 16546
rect 33152 16522 33180 17546
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34060 16584 34112 16590
rect 34060 16526 34112 16532
rect 33140 16516 33192 16522
rect 33140 16458 33192 16464
rect 32588 16448 32640 16454
rect 32588 16390 32640 16396
rect 32956 16448 33008 16454
rect 32956 16390 33008 16396
rect 32128 16040 32180 16046
rect 32128 15982 32180 15988
rect 31852 15904 31904 15910
rect 31852 15846 31904 15852
rect 31944 15904 31996 15910
rect 31944 15846 31996 15852
rect 31864 15026 31892 15846
rect 31852 15020 31904 15026
rect 31852 14962 31904 14968
rect 31758 9072 31814 9081
rect 31758 9007 31814 9016
rect 31404 8214 31892 8242
rect 31300 8084 31352 8090
rect 31300 8026 31352 8032
rect 31312 7478 31340 8026
rect 31576 7744 31628 7750
rect 31576 7686 31628 7692
rect 31588 7546 31616 7686
rect 31576 7540 31628 7546
rect 31576 7482 31628 7488
rect 31300 7472 31352 7478
rect 31352 7420 31432 7426
rect 31300 7414 31432 7420
rect 31312 7398 31432 7414
rect 31300 7336 31352 7342
rect 31300 7278 31352 7284
rect 31312 6458 31340 7278
rect 31404 6662 31432 7398
rect 31864 7274 31892 8214
rect 31956 7546 31984 15846
rect 32140 14890 32168 15982
rect 32600 15026 32628 16390
rect 32680 16040 32732 16046
rect 32680 15982 32732 15988
rect 32692 15162 32720 15982
rect 32680 15156 32732 15162
rect 32680 15098 32732 15104
rect 32588 15020 32640 15026
rect 32588 14962 32640 14968
rect 32036 14884 32088 14890
rect 32036 14826 32088 14832
rect 32128 14884 32180 14890
rect 32128 14826 32180 14832
rect 32048 14618 32076 14826
rect 32036 14612 32088 14618
rect 32036 14554 32088 14560
rect 32140 14006 32168 14826
rect 32128 14000 32180 14006
rect 32128 13942 32180 13948
rect 32140 12850 32168 13942
rect 32128 12844 32180 12850
rect 32128 12786 32180 12792
rect 32404 12776 32456 12782
rect 32404 12718 32456 12724
rect 32416 12442 32444 12718
rect 32404 12436 32456 12442
rect 32404 12378 32456 12384
rect 32864 12368 32916 12374
rect 32864 12310 32916 12316
rect 32876 12170 32904 12310
rect 32864 12164 32916 12170
rect 32864 12106 32916 12112
rect 32772 10600 32824 10606
rect 32772 10542 32824 10548
rect 32784 9994 32812 10542
rect 32772 9988 32824 9994
rect 32772 9930 32824 9936
rect 32784 8974 32812 9930
rect 32772 8968 32824 8974
rect 32772 8910 32824 8916
rect 32968 8922 32996 16390
rect 33152 16182 33180 16458
rect 33140 16176 33192 16182
rect 33140 16118 33192 16124
rect 33048 15428 33100 15434
rect 33048 15370 33100 15376
rect 33060 14890 33088 15370
rect 33152 15162 33180 16118
rect 34072 15910 34100 16526
rect 34336 16516 34388 16522
rect 34336 16458 34388 16464
rect 34348 16425 34376 16458
rect 34334 16416 34390 16425
rect 34334 16351 34390 16360
rect 33416 15904 33468 15910
rect 33416 15846 33468 15852
rect 34060 15904 34112 15910
rect 34060 15846 34112 15852
rect 33140 15156 33192 15162
rect 33140 15098 33192 15104
rect 33048 14884 33100 14890
rect 33048 14826 33100 14832
rect 33152 12918 33180 15098
rect 33428 15094 33456 15846
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34796 15496 34848 15502
rect 34796 15438 34848 15444
rect 34704 15428 34756 15434
rect 34704 15370 34756 15376
rect 33416 15088 33468 15094
rect 33416 15030 33468 15036
rect 33968 14952 34020 14958
rect 33968 14894 34020 14900
rect 33980 14618 34008 14894
rect 33968 14612 34020 14618
rect 33968 14554 34020 14560
rect 34716 14521 34744 15370
rect 34808 14822 34836 15438
rect 34796 14816 34848 14822
rect 34796 14758 34848 14764
rect 34702 14512 34758 14521
rect 34702 14447 34758 14456
rect 34428 14408 34480 14414
rect 34428 14350 34480 14356
rect 33140 12912 33192 12918
rect 33140 12854 33192 12860
rect 33152 12442 33180 12854
rect 33876 12844 33928 12850
rect 33876 12786 33928 12792
rect 33888 12646 33916 12786
rect 33876 12640 33928 12646
rect 33876 12582 33928 12588
rect 33140 12436 33192 12442
rect 33140 12378 33192 12384
rect 33888 12306 33916 12582
rect 33876 12300 33928 12306
rect 33876 12242 33928 12248
rect 34440 12238 34468 14350
rect 34808 14346 34836 14758
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34796 14340 34848 14346
rect 34796 14282 34848 14288
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35348 12776 35400 12782
rect 35348 12718 35400 12724
rect 35360 12617 35388 12718
rect 35346 12608 35402 12617
rect 34934 12540 35242 12549
rect 35346 12543 35402 12552
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34428 12232 34480 12238
rect 34428 12174 34480 12180
rect 34150 11248 34206 11257
rect 34150 11183 34206 11192
rect 34164 11150 34192 11183
rect 34440 11150 34468 12174
rect 34520 11756 34572 11762
rect 34520 11698 34572 11704
rect 34152 11144 34204 11150
rect 34152 11086 34204 11092
rect 34428 11144 34480 11150
rect 34428 11086 34480 11092
rect 33508 11008 33560 11014
rect 33508 10950 33560 10956
rect 33520 10742 33548 10950
rect 33508 10736 33560 10742
rect 33508 10678 33560 10684
rect 34440 9586 34468 11086
rect 34532 11082 34560 11698
rect 34796 11688 34848 11694
rect 34796 11630 34848 11636
rect 34520 11076 34572 11082
rect 34520 11018 34572 11024
rect 34520 10736 34572 10742
rect 34808 10713 34836 11630
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34980 11076 35032 11082
rect 34980 11018 35032 11024
rect 34992 10810 35020 11018
rect 34980 10804 35032 10810
rect 34980 10746 35032 10752
rect 34520 10678 34572 10684
rect 34794 10704 34850 10713
rect 34060 9580 34112 9586
rect 34060 9522 34112 9528
rect 34244 9580 34296 9586
rect 34244 9522 34296 9528
rect 34428 9580 34480 9586
rect 34428 9522 34480 9528
rect 33048 9376 33100 9382
rect 33048 9318 33100 9324
rect 33060 9042 33088 9318
rect 33048 9036 33100 9042
rect 33048 8978 33100 8984
rect 32404 8424 32456 8430
rect 32404 8366 32456 8372
rect 32496 8424 32548 8430
rect 32496 8366 32548 8372
rect 32416 8090 32444 8366
rect 32404 8084 32456 8090
rect 32404 8026 32456 8032
rect 32508 7886 32536 8366
rect 32784 8294 32812 8910
rect 32968 8894 33088 8922
rect 32772 8288 32824 8294
rect 32772 8230 32824 8236
rect 32496 7880 32548 7886
rect 32496 7822 32548 7828
rect 31944 7540 31996 7546
rect 31944 7482 31996 7488
rect 32220 7404 32272 7410
rect 32220 7346 32272 7352
rect 31852 7268 31904 7274
rect 31852 7210 31904 7216
rect 31864 7002 31892 7210
rect 31852 6996 31904 7002
rect 31852 6938 31904 6944
rect 31668 6928 31720 6934
rect 31668 6870 31720 6876
rect 31760 6928 31812 6934
rect 31760 6870 31812 6876
rect 31576 6860 31628 6866
rect 31576 6802 31628 6808
rect 31588 6662 31616 6802
rect 31392 6656 31444 6662
rect 31392 6598 31444 6604
rect 31576 6656 31628 6662
rect 31576 6598 31628 6604
rect 31208 6452 31260 6458
rect 31208 6394 31260 6400
rect 31300 6452 31352 6458
rect 31300 6394 31352 6400
rect 31116 6316 31168 6322
rect 31116 6258 31168 6264
rect 31300 6112 31352 6118
rect 31300 6054 31352 6060
rect 31036 5868 31156 5896
rect 30838 5808 30894 5817
rect 30748 5772 30800 5778
rect 30838 5743 30894 5752
rect 31024 5772 31076 5778
rect 30748 5714 30800 5720
rect 31024 5714 31076 5720
rect 30656 5704 30708 5710
rect 30656 5646 30708 5652
rect 30472 5228 30524 5234
rect 30472 5170 30524 5176
rect 30484 4690 30512 5170
rect 30760 5030 30788 5714
rect 31036 5166 31064 5714
rect 30840 5160 30892 5166
rect 30840 5102 30892 5108
rect 31024 5160 31076 5166
rect 31024 5102 31076 5108
rect 30748 5024 30800 5030
rect 30748 4966 30800 4972
rect 30288 4684 30340 4690
rect 30288 4626 30340 4632
rect 30472 4684 30524 4690
rect 30472 4626 30524 4632
rect 30852 4622 30880 5102
rect 30840 4616 30892 4622
rect 30840 4558 30892 4564
rect 29920 4548 29972 4554
rect 29920 4490 29972 4496
rect 29748 4406 30144 4434
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 29092 4140 29144 4146
rect 29092 4082 29144 4088
rect 30116 4078 30144 4406
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 28724 4072 28776 4078
rect 28724 4014 28776 4020
rect 29828 4072 29880 4078
rect 29828 4014 29880 4020
rect 30104 4072 30156 4078
rect 30104 4014 30156 4020
rect 29000 3936 29052 3942
rect 29000 3878 29052 3884
rect 29012 3602 29040 3878
rect 29840 3738 29868 4014
rect 29828 3732 29880 3738
rect 29828 3674 29880 3680
rect 30116 3670 30144 4014
rect 30852 3942 30880 4558
rect 31128 4486 31156 5868
rect 31312 5642 31340 6054
rect 31404 5914 31432 6598
rect 31680 6322 31708 6870
rect 31772 6798 31800 6870
rect 31864 6798 31892 6938
rect 31760 6792 31812 6798
rect 31760 6734 31812 6740
rect 31852 6792 31904 6798
rect 31852 6734 31904 6740
rect 31944 6792 31996 6798
rect 31944 6734 31996 6740
rect 31484 6316 31536 6322
rect 31484 6258 31536 6264
rect 31668 6316 31720 6322
rect 31668 6258 31720 6264
rect 31496 6202 31524 6258
rect 31772 6202 31800 6734
rect 31956 6662 31984 6734
rect 31944 6656 31996 6662
rect 31944 6598 31996 6604
rect 32232 6458 32260 7346
rect 32404 6928 32456 6934
rect 32508 6914 32536 7822
rect 32588 7812 32640 7818
rect 32588 7754 32640 7760
rect 32600 7546 32628 7754
rect 32680 7744 32732 7750
rect 32680 7686 32732 7692
rect 32588 7540 32640 7546
rect 32588 7482 32640 7488
rect 32692 7410 32720 7686
rect 32680 7404 32732 7410
rect 32680 7346 32732 7352
rect 32784 7342 32812 8230
rect 33060 7750 33088 8894
rect 33140 8900 33192 8906
rect 33140 8842 33192 8848
rect 33152 8566 33180 8842
rect 34072 8809 34100 9522
rect 34256 9178 34284 9522
rect 34244 9172 34296 9178
rect 34244 9114 34296 9120
rect 34058 8800 34114 8809
rect 34058 8735 34114 8744
rect 33140 8560 33192 8566
rect 33140 8502 33192 8508
rect 33152 7954 33180 8502
rect 34256 8498 34284 9114
rect 34244 8492 34296 8498
rect 34244 8434 34296 8440
rect 33140 7948 33192 7954
rect 33140 7890 33192 7896
rect 33048 7744 33100 7750
rect 33048 7686 33100 7692
rect 32864 7540 32916 7546
rect 32864 7482 32916 7488
rect 32772 7336 32824 7342
rect 32772 7278 32824 7284
rect 32456 6886 32536 6914
rect 32404 6870 32456 6876
rect 32416 6730 32444 6870
rect 32876 6798 32904 7482
rect 33060 7206 33088 7686
rect 33152 7546 33180 7890
rect 34336 7880 34388 7886
rect 34256 7828 34336 7834
rect 34256 7822 34388 7828
rect 34256 7806 34376 7822
rect 33140 7540 33192 7546
rect 33140 7482 33192 7488
rect 33140 7404 33192 7410
rect 33140 7346 33192 7352
rect 33048 7200 33100 7206
rect 33048 7142 33100 7148
rect 33060 6934 33088 7142
rect 33048 6928 33100 6934
rect 33048 6870 33100 6876
rect 32588 6792 32640 6798
rect 32588 6734 32640 6740
rect 32864 6792 32916 6798
rect 32864 6734 32916 6740
rect 32312 6724 32364 6730
rect 32312 6666 32364 6672
rect 32404 6724 32456 6730
rect 32404 6666 32456 6672
rect 32324 6458 32352 6666
rect 32220 6452 32272 6458
rect 32220 6394 32272 6400
rect 32312 6452 32364 6458
rect 32312 6394 32364 6400
rect 31496 6174 31800 6202
rect 31392 5908 31444 5914
rect 31392 5850 31444 5856
rect 31496 5710 31524 6174
rect 32496 6112 32548 6118
rect 32496 6054 32548 6060
rect 32036 5840 32088 5846
rect 31666 5808 31722 5817
rect 32036 5782 32088 5788
rect 31666 5743 31668 5752
rect 31720 5743 31722 5752
rect 31668 5714 31720 5720
rect 31484 5704 31536 5710
rect 31484 5646 31536 5652
rect 31300 5636 31352 5642
rect 31300 5578 31352 5584
rect 31116 4480 31168 4486
rect 31116 4422 31168 4428
rect 31128 4282 31156 4422
rect 31116 4276 31168 4282
rect 31116 4218 31168 4224
rect 31312 4214 31340 5578
rect 32048 4622 32076 5782
rect 32508 5574 32536 6054
rect 32600 5778 32628 6734
rect 33048 6384 33100 6390
rect 33048 6326 33100 6332
rect 32864 6316 32916 6322
rect 32864 6258 32916 6264
rect 32876 6225 32904 6258
rect 33060 6254 33088 6326
rect 33048 6248 33100 6254
rect 32862 6216 32918 6225
rect 33048 6190 33100 6196
rect 33152 6186 33180 7346
rect 33508 7336 33560 7342
rect 33508 7278 33560 7284
rect 33520 7002 33548 7278
rect 34256 7206 34284 7806
rect 34244 7200 34296 7206
rect 34244 7142 34296 7148
rect 33508 6996 33560 7002
rect 33508 6938 33560 6944
rect 34058 6896 34114 6905
rect 33416 6860 33468 6866
rect 34058 6831 34114 6840
rect 33416 6802 33468 6808
rect 33428 6730 33456 6802
rect 34072 6798 34100 6831
rect 34256 6798 34284 7142
rect 34440 6798 34468 9522
rect 34532 6914 34560 10678
rect 34794 10639 34850 10648
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34794 8800 34850 8809
rect 34794 8735 34850 8744
rect 34808 8566 34836 8735
rect 34796 8560 34848 8566
rect 34796 8502 34848 8508
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34704 7812 34756 7818
rect 34704 7754 34756 7760
rect 34532 6886 34652 6914
rect 34716 6905 34744 7754
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34060 6792 34112 6798
rect 34060 6734 34112 6740
rect 34244 6792 34296 6798
rect 34244 6734 34296 6740
rect 34428 6792 34480 6798
rect 34428 6734 34480 6740
rect 33416 6724 33468 6730
rect 33416 6666 33468 6672
rect 33428 6458 33456 6666
rect 33416 6452 33468 6458
rect 33416 6394 33468 6400
rect 34428 6316 34480 6322
rect 34428 6258 34480 6264
rect 32862 6151 32918 6160
rect 33140 6180 33192 6186
rect 32876 5914 32904 6151
rect 33140 6122 33192 6128
rect 33232 6112 33284 6118
rect 33232 6054 33284 6060
rect 32864 5908 32916 5914
rect 32864 5850 32916 5856
rect 33244 5846 33272 6054
rect 33232 5840 33284 5846
rect 33232 5782 33284 5788
rect 34152 5840 34204 5846
rect 34152 5782 34204 5788
rect 32588 5772 32640 5778
rect 32588 5714 32640 5720
rect 33140 5636 33192 5642
rect 33140 5578 33192 5584
rect 33968 5636 34020 5642
rect 33968 5578 34020 5584
rect 32496 5568 32548 5574
rect 32496 5510 32548 5516
rect 33152 5370 33180 5578
rect 33140 5364 33192 5370
rect 33140 5306 33192 5312
rect 33152 4826 33180 5306
rect 33980 5234 34008 5578
rect 34164 5234 34192 5782
rect 34440 5710 34468 6258
rect 34428 5704 34480 5710
rect 34428 5646 34480 5652
rect 34440 5234 34468 5646
rect 34624 5574 34652 6886
rect 34702 6896 34758 6905
rect 34702 6831 34758 6840
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34612 5568 34664 5574
rect 34612 5510 34664 5516
rect 33968 5228 34020 5234
rect 33968 5170 34020 5176
rect 34152 5228 34204 5234
rect 34152 5170 34204 5176
rect 34428 5228 34480 5234
rect 34428 5170 34480 5176
rect 34060 5024 34112 5030
rect 34060 4966 34112 4972
rect 33140 4820 33192 4826
rect 33140 4762 33192 4768
rect 32404 4752 32456 4758
rect 32404 4694 32456 4700
rect 31392 4616 31444 4622
rect 31392 4558 31444 4564
rect 32036 4616 32088 4622
rect 32036 4558 32088 4564
rect 31404 4214 31432 4558
rect 32416 4282 32444 4694
rect 33232 4548 33284 4554
rect 33232 4490 33284 4496
rect 33244 4282 33272 4490
rect 32404 4276 32456 4282
rect 32404 4218 32456 4224
rect 33232 4276 33284 4282
rect 33232 4218 33284 4224
rect 31300 4208 31352 4214
rect 31300 4150 31352 4156
rect 31392 4208 31444 4214
rect 31392 4150 31444 4156
rect 30840 3936 30892 3942
rect 30840 3878 30892 3884
rect 30104 3664 30156 3670
rect 30104 3606 30156 3612
rect 29000 3596 29052 3602
rect 29000 3538 29052 3544
rect 30852 3534 30880 3878
rect 34072 3534 34100 4966
rect 34440 4486 34468 5170
rect 35348 5160 35400 5166
rect 35348 5102 35400 5108
rect 35360 5001 35388 5102
rect 35346 4992 35402 5001
rect 34934 4924 35242 4933
rect 35346 4927 35402 4936
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34428 4480 34480 4486
rect 34428 4422 34480 4428
rect 34440 4214 34468 4422
rect 34428 4208 34480 4214
rect 34428 4150 34480 4156
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 30840 3528 30892 3534
rect 30840 3470 30892 3476
rect 34060 3528 34112 3534
rect 34060 3470 34112 3476
rect 34336 3460 34388 3466
rect 34336 3402 34388 3408
rect 21548 3392 21600 3398
rect 21548 3334 21600 3340
rect 34348 3097 34376 3402
rect 34334 3088 34390 3097
rect 34334 3023 34390 3032
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 18142 1184 18198 1193
rect 18142 1119 18198 1128
<< via2 >>
rect 1214 37304 1270 37360
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 1306 35400 1362 35456
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 1306 33496 1362 33552
rect 1398 31592 1454 31648
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 1306 29688 1362 29744
rect 1306 27784 1362 27840
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 1858 26308 1914 26344
rect 1858 26288 1860 26308
rect 1860 26288 1912 26308
rect 1912 26288 1914 26308
rect 1306 25880 1362 25936
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4158 28076 4214 28112
rect 4158 28056 4160 28076
rect 4160 28056 4212 28076
rect 4212 28056 4214 28076
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 1214 23976 1270 24032
rect 1858 22500 1914 22536
rect 1858 22480 1860 22500
rect 1860 22480 1912 22500
rect 1912 22480 1914 22500
rect 1306 22072 1362 22128
rect 1306 20168 1362 20224
rect 1306 18264 1362 18320
rect 1398 16360 1454 16416
rect 1306 14456 1362 14512
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 5722 26580 5778 26616
rect 5722 26560 5724 26580
rect 5724 26560 5776 26580
rect 5776 26560 5778 26580
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 1306 12552 1362 12608
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 1306 10648 1362 10704
rect 3146 10648 3202 10704
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 5078 11076 5134 11112
rect 5078 11056 5080 11076
rect 5080 11056 5132 11076
rect 5132 11056 5134 11076
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 1306 8744 1362 8800
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 9770 33904 9826 33960
rect 9862 33632 9918 33688
rect 8942 28056 8998 28112
rect 10506 33652 10562 33688
rect 10506 33632 10508 33652
rect 10508 33632 10560 33652
rect 10560 33632 10562 33652
rect 10598 26988 10654 27024
rect 10598 26968 10600 26988
rect 10600 26968 10652 26988
rect 10652 26968 10654 26988
rect 10506 26832 10562 26888
rect 10322 26016 10378 26072
rect 10598 25336 10654 25392
rect 8390 21256 8446 21312
rect 5906 10668 5962 10704
rect 5906 10648 5908 10668
rect 5908 10648 5960 10668
rect 5960 10648 5962 10668
rect 5354 9560 5410 9616
rect 6090 9560 6146 9616
rect 11610 34468 11666 34504
rect 11610 34448 11612 34468
rect 11612 34448 11664 34468
rect 11664 34448 11666 34468
rect 13726 33904 13782 33960
rect 12070 32716 12072 32736
rect 12072 32716 12124 32736
rect 12124 32716 12126 32736
rect 12070 32680 12126 32716
rect 11058 30268 11060 30288
rect 11060 30268 11112 30288
rect 11112 30268 11114 30288
rect 11058 30232 11114 30268
rect 11794 26832 11850 26888
rect 10966 25780 10968 25800
rect 10968 25780 11020 25800
rect 11020 25780 11022 25800
rect 10966 25744 11022 25780
rect 10874 25336 10930 25392
rect 11702 26460 11704 26480
rect 11704 26460 11756 26480
rect 11756 26460 11758 26480
rect 11702 26424 11758 26460
rect 10414 19624 10470 19680
rect 10782 19352 10838 19408
rect 9034 15308 9036 15328
rect 9036 15308 9088 15328
rect 9088 15308 9090 15328
rect 9034 15272 9090 15308
rect 6826 8916 6828 8936
rect 6828 8916 6880 8936
rect 6880 8916 6882 8936
rect 6826 8880 6882 8916
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 9770 9968 9826 10024
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 12714 25492 12770 25528
rect 12714 25472 12716 25492
rect 12716 25472 12768 25492
rect 12768 25472 12770 25492
rect 12070 22344 12126 22400
rect 13450 29008 13506 29064
rect 13358 24656 13414 24712
rect 14278 30268 14280 30288
rect 14280 30268 14332 30288
rect 14332 30268 14334 30288
rect 14278 30232 14334 30268
rect 13634 25336 13690 25392
rect 12438 19372 12494 19408
rect 12438 19352 12440 19372
rect 12440 19352 12492 19372
rect 12492 19352 12494 19372
rect 11794 13368 11850 13424
rect 11978 11056 12034 11112
rect 12622 12960 12678 13016
rect 14278 26560 14334 26616
rect 14554 29008 14610 29064
rect 14922 27376 14978 27432
rect 14922 26560 14978 26616
rect 17038 32680 17094 32736
rect 17590 33632 17646 33688
rect 16302 25744 16358 25800
rect 16302 24792 16358 24848
rect 15842 23604 15844 23624
rect 15844 23604 15896 23624
rect 15896 23604 15898 23624
rect 15842 23568 15898 23604
rect 16210 22344 16266 22400
rect 17406 26832 17462 26888
rect 17222 26696 17278 26752
rect 17130 26560 17186 26616
rect 17774 26968 17830 27024
rect 18510 30268 18512 30288
rect 18512 30268 18564 30288
rect 18564 30268 18566 30288
rect 18510 30232 18566 30268
rect 20810 34484 20812 34504
rect 20812 34484 20864 34504
rect 20864 34484 20866 34504
rect 20810 34448 20866 34484
rect 19798 30368 19854 30424
rect 19154 29008 19210 29064
rect 18050 26832 18106 26888
rect 17222 26288 17278 26344
rect 17314 24792 17370 24848
rect 17222 24692 17224 24712
rect 17224 24692 17276 24712
rect 17276 24692 17278 24712
rect 17222 24656 17278 24692
rect 17590 24656 17646 24712
rect 18050 26560 18106 26616
rect 19154 26560 19210 26616
rect 18878 26016 18934 26072
rect 19154 25492 19210 25528
rect 19154 25472 19156 25492
rect 19156 25472 19208 25492
rect 19208 25472 19210 25492
rect 19062 25336 19118 25392
rect 19154 24112 19210 24168
rect 13174 15272 13230 15328
rect 1306 6840 1362 6896
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 12438 10684 12440 10704
rect 12440 10684 12492 10704
rect 12492 10684 12494 10704
rect 12438 10648 12494 10684
rect 14738 16768 14794 16824
rect 15658 19624 15714 19680
rect 14646 12688 14702 12744
rect 12438 6860 12494 6896
rect 12438 6840 12440 6860
rect 12440 6840 12492 6860
rect 12492 6840 12494 6860
rect 15290 16668 15292 16688
rect 15292 16668 15344 16688
rect 15344 16668 15346 16688
rect 15290 16632 15346 16668
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 16026 13640 16082 13696
rect 16394 13640 16450 13696
rect 16670 11636 16672 11656
rect 16672 11636 16724 11656
rect 16724 11636 16726 11656
rect 16670 11600 16726 11636
rect 17222 16532 17224 16552
rect 17224 16532 17276 16552
rect 17276 16532 17278 16552
rect 17222 16496 17278 16532
rect 17682 18692 17738 18728
rect 17682 18672 17684 18692
rect 17684 18672 17736 18692
rect 17736 18672 17738 18692
rect 17130 10684 17132 10704
rect 17132 10684 17184 10704
rect 17184 10684 17186 10704
rect 17130 10648 17186 10684
rect 17590 12844 17646 12880
rect 17590 12824 17592 12844
rect 17592 12824 17644 12844
rect 17644 12824 17646 12844
rect 17590 11620 17646 11656
rect 17590 11600 17592 11620
rect 17592 11600 17644 11620
rect 17644 11600 17646 11620
rect 16946 9968 17002 10024
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 1306 4936 1362 4992
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 1306 3032 1362 3088
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 19246 22480 19302 22536
rect 19246 21392 19302 21448
rect 19982 21256 20038 21312
rect 22926 33804 22928 33824
rect 22928 33804 22980 33824
rect 22980 33804 22982 33824
rect 22926 33768 22982 33804
rect 19062 12960 19118 13016
rect 19154 12552 19210 12608
rect 18326 10668 18382 10704
rect 18326 10648 18328 10668
rect 18328 10648 18380 10668
rect 18380 10648 18382 10668
rect 19338 12300 19394 12336
rect 19338 12280 19340 12300
rect 19340 12280 19392 12300
rect 19392 12280 19394 12300
rect 19706 12588 19708 12608
rect 19708 12588 19760 12608
rect 19760 12588 19762 12608
rect 19706 12552 19762 12588
rect 19522 11192 19578 11248
rect 19614 11076 19670 11112
rect 19614 11056 19616 11076
rect 19616 11056 19668 11076
rect 19668 11056 19670 11076
rect 20534 20868 20590 20904
rect 20994 26868 20996 26888
rect 20996 26868 21048 26888
rect 21048 26868 21050 26888
rect 20994 26832 21050 26868
rect 22098 26696 22154 26752
rect 21914 25744 21970 25800
rect 21730 24284 21732 24304
rect 21732 24284 21784 24304
rect 21784 24284 21786 24304
rect 21730 24248 21786 24284
rect 22466 25744 22522 25800
rect 22650 26696 22706 26752
rect 23018 31320 23074 31376
rect 23662 33768 23718 33824
rect 24122 33804 24124 33824
rect 24124 33804 24176 33824
rect 24176 33804 24178 33824
rect 22466 24248 22522 24304
rect 24122 33768 24178 33804
rect 23570 27512 23626 27568
rect 23662 27412 23664 27432
rect 23664 27412 23716 27432
rect 23716 27412 23718 27432
rect 23662 27376 23718 27412
rect 27434 35436 27436 35456
rect 27436 35436 27488 35456
rect 27488 35436 27490 35456
rect 27434 35400 27490 35436
rect 26238 35128 26294 35184
rect 34334 35572 34336 35592
rect 34336 35572 34388 35592
rect 34388 35572 34390 35592
rect 34334 35536 34390 35572
rect 20534 20848 20536 20868
rect 20536 20848 20588 20868
rect 20588 20848 20590 20868
rect 20994 20168 21050 20224
rect 21546 18572 21548 18592
rect 21548 18572 21600 18592
rect 21600 18572 21602 18592
rect 21546 18536 21602 18572
rect 21822 18964 21878 19000
rect 21822 18944 21824 18964
rect 21824 18944 21876 18964
rect 21876 18944 21878 18964
rect 22098 20576 22154 20632
rect 22466 20440 22522 20496
rect 22098 18264 22154 18320
rect 23386 21936 23442 21992
rect 23202 19660 23204 19680
rect 23204 19660 23256 19680
rect 23256 19660 23258 19680
rect 23202 19624 23258 19660
rect 20350 9596 20352 9616
rect 20352 9596 20404 9616
rect 20404 9596 20406 9616
rect 20350 9560 20406 9596
rect 18602 6840 18658 6896
rect 20626 9016 20682 9072
rect 21730 14612 21786 14648
rect 21730 14592 21732 14612
rect 21732 14592 21784 14612
rect 21784 14592 21786 14612
rect 22190 16108 22246 16144
rect 22190 16088 22192 16108
rect 22192 16088 22244 16108
rect 22244 16088 22246 16108
rect 22466 15580 22468 15600
rect 22468 15580 22520 15600
rect 22520 15580 22522 15600
rect 22466 15544 22522 15580
rect 21362 9152 21418 9208
rect 21638 8608 21694 8664
rect 24122 21120 24178 21176
rect 24306 21528 24362 21584
rect 24398 20304 24454 20360
rect 23938 18264 23994 18320
rect 22006 9036 22062 9072
rect 22466 9424 22522 9480
rect 22006 9016 22008 9036
rect 22008 9016 22060 9036
rect 22060 9016 22062 9036
rect 22282 8780 22284 8800
rect 22284 8780 22336 8800
rect 22336 8780 22338 8800
rect 22282 8744 22338 8780
rect 22466 8608 22522 8664
rect 22650 9596 22652 9616
rect 22652 9596 22704 9616
rect 22704 9596 22706 9616
rect 22650 9560 22706 9596
rect 22742 9016 22798 9072
rect 23110 10784 23166 10840
rect 22926 10512 22982 10568
rect 23386 12688 23442 12744
rect 24674 21528 24730 21584
rect 24582 18944 24638 19000
rect 25318 20440 25374 20496
rect 24858 20052 24914 20088
rect 24858 20032 24860 20052
rect 24860 20032 24912 20052
rect 24912 20032 24914 20052
rect 24030 12144 24086 12200
rect 25318 18264 25374 18320
rect 27066 31748 27122 31784
rect 27066 31728 27068 31748
rect 27068 31728 27120 31748
rect 27120 31728 27122 31748
rect 26422 29008 26478 29064
rect 26238 26324 26240 26344
rect 26240 26324 26292 26344
rect 26292 26324 26294 26344
rect 26238 26288 26294 26324
rect 26330 26152 26386 26208
rect 25870 23976 25926 24032
rect 26606 26832 26662 26888
rect 26422 24384 26478 24440
rect 26698 24384 26754 24440
rect 26514 24248 26570 24304
rect 26146 23840 26202 23896
rect 26330 23724 26386 23760
rect 26330 23704 26332 23724
rect 26332 23704 26384 23724
rect 26384 23704 26386 23724
rect 25686 18264 25742 18320
rect 25962 19352 26018 19408
rect 25962 17876 26018 17912
rect 25962 17856 25964 17876
rect 25964 17856 26016 17876
rect 26016 17856 26018 17876
rect 26422 21392 26478 21448
rect 26606 20168 26662 20224
rect 27066 31320 27122 31376
rect 27526 30368 27582 30424
rect 27158 27512 27214 27568
rect 26974 24112 27030 24168
rect 26790 23976 26846 24032
rect 27618 25608 27674 25664
rect 27618 23432 27674 23488
rect 27894 31728 27950 31784
rect 27802 24384 27858 24440
rect 27802 24012 27804 24032
rect 27804 24012 27856 24032
rect 27856 24012 27858 24032
rect 27802 23976 27858 24012
rect 26790 20324 26846 20360
rect 26790 20304 26792 20324
rect 26792 20304 26844 20324
rect 26844 20304 26846 20324
rect 26514 19352 26570 19408
rect 27066 16632 27122 16688
rect 26146 12416 26202 12472
rect 26882 15020 26938 15056
rect 26882 15000 26884 15020
rect 26884 15000 26936 15020
rect 26936 15000 26938 15020
rect 27066 14068 27122 14104
rect 27066 14048 27068 14068
rect 27068 14048 27120 14068
rect 27120 14048 27122 14068
rect 27986 27276 27988 27296
rect 27988 27276 28040 27296
rect 28040 27276 28042 27296
rect 27986 27240 28042 27276
rect 27986 23568 28042 23624
rect 27710 21936 27766 21992
rect 27894 21936 27950 21992
rect 27434 19352 27490 19408
rect 27342 16360 27398 16416
rect 27342 13368 27398 13424
rect 26698 10512 26754 10568
rect 27158 10376 27214 10432
rect 27710 14184 27766 14240
rect 28538 24404 28594 24440
rect 28538 24384 28540 24404
rect 28540 24384 28592 24404
rect 28592 24384 28594 24404
rect 28354 24012 28356 24032
rect 28356 24012 28408 24032
rect 28408 24012 28410 24032
rect 28354 23976 28410 24012
rect 28354 20848 28410 20904
rect 27894 14320 27950 14376
rect 28906 26444 28962 26480
rect 28906 26424 28908 26444
rect 28908 26424 28960 26444
rect 28960 26424 28962 26444
rect 28722 23568 28778 23624
rect 29366 28364 29368 28384
rect 29368 28364 29420 28384
rect 29420 28364 29422 28384
rect 29366 28328 29422 28364
rect 29274 22380 29276 22400
rect 29276 22380 29328 22400
rect 29328 22380 29330 22400
rect 29274 22344 29330 22380
rect 28998 22072 29054 22128
rect 29274 21800 29330 21856
rect 29182 21664 29238 21720
rect 29734 22516 29736 22536
rect 29736 22516 29788 22536
rect 29788 22516 29790 22536
rect 29734 22480 29790 22516
rect 26514 9580 26570 9616
rect 26514 9560 26516 9580
rect 26516 9560 26568 9580
rect 26568 9560 26570 9580
rect 26330 9444 26386 9480
rect 26330 9424 26332 9444
rect 26332 9424 26384 9444
rect 26384 9424 26386 9444
rect 28170 12824 28226 12880
rect 28722 14592 28778 14648
rect 28814 14356 28816 14376
rect 28816 14356 28868 14376
rect 28868 14356 28870 14376
rect 28814 14320 28870 14356
rect 28630 14184 28686 14240
rect 28262 11600 28318 11656
rect 28262 10784 28318 10840
rect 28722 10376 28778 10432
rect 28446 9152 28502 9208
rect 28814 10104 28870 10160
rect 30010 16532 30012 16552
rect 30012 16532 30064 16552
rect 30064 16532 30066 16552
rect 30010 16496 30066 16532
rect 29550 10648 29606 10704
rect 29642 10104 29698 10160
rect 29734 8880 29790 8936
rect 30746 21936 30802 21992
rect 31022 21936 31078 21992
rect 31022 21392 31078 21448
rect 30746 21292 30748 21312
rect 30748 21292 30800 21312
rect 30800 21292 30802 21312
rect 30746 21256 30802 21292
rect 30838 21120 30894 21176
rect 31114 21120 31170 21176
rect 30562 15156 30618 15192
rect 30562 15136 30564 15156
rect 30564 15136 30616 15156
rect 30616 15136 30618 15156
rect 30470 9968 30526 10024
rect 34334 33496 34390 33552
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34794 31592 34850 31648
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34518 29688 34574 29744
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 35346 27784 35402 27840
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34794 25880 34850 25936
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34794 23976 34850 24032
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34794 22072 34850 22128
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35346 20168 35402 20224
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 29642 6160 29698 6216
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34150 18708 34152 18728
rect 34152 18708 34204 18728
rect 34204 18708 34206 18728
rect 34150 18672 34206 18708
rect 34794 18284 34850 18320
rect 34794 18264 34796 18284
rect 34796 18264 34848 18284
rect 34848 18264 34850 18284
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 31758 9016 31814 9072
rect 34334 16360 34390 16416
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34702 14456 34758 14512
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 35346 12552 35402 12608
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34150 11192 34206 11248
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 30838 5752 30894 5808
rect 34058 8744 34114 8800
rect 31666 5772 31722 5808
rect 31666 5752 31668 5772
rect 31668 5752 31720 5772
rect 31720 5752 31722 5772
rect 32862 6160 32918 6216
rect 34058 6840 34114 6896
rect 34794 10648 34850 10704
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34794 8744 34850 8800
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34702 6840 34758 6896
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35346 4936 35402 4992
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34334 3032 34390 3088
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 18142 1128 18198 1184
<< metal3 >>
rect 0 37362 800 37392
rect 1209 37362 1275 37365
rect 0 37360 1275 37362
rect 0 37304 1214 37360
rect 1270 37304 1275 37360
rect 0 37302 1275 37304
rect 0 37272 800 37302
rect 1209 37299 1275 37302
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 34329 35594 34395 35597
rect 34329 35592 35450 35594
rect 34329 35536 34334 35592
rect 34390 35536 35450 35592
rect 34329 35534 35450 35536
rect 34329 35531 34395 35534
rect 0 35458 800 35488
rect 1301 35458 1367 35461
rect 27429 35460 27495 35461
rect 27429 35458 27476 35460
rect 0 35456 1367 35458
rect 0 35400 1306 35456
rect 1362 35400 1367 35456
rect 0 35398 1367 35400
rect 27384 35456 27476 35458
rect 27384 35400 27434 35456
rect 27384 35398 27476 35400
rect 0 35368 800 35398
rect 1301 35395 1367 35398
rect 27429 35396 27476 35398
rect 27540 35396 27546 35460
rect 35390 35458 35450 35534
rect 35673 35458 36473 35488
rect 35390 35398 36473 35458
rect 27429 35395 27495 35396
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 35673 35368 36473 35398
rect 34930 35327 35246 35328
rect 26233 35186 26299 35189
rect 26550 35186 26556 35188
rect 26233 35184 26556 35186
rect 26233 35128 26238 35184
rect 26294 35128 26556 35184
rect 26233 35126 26556 35128
rect 26233 35123 26299 35126
rect 26550 35124 26556 35126
rect 26620 35124 26626 35188
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 11605 34506 11671 34509
rect 20805 34506 20871 34509
rect 11605 34504 20871 34506
rect 11605 34448 11610 34504
rect 11666 34448 20810 34504
rect 20866 34448 20871 34504
rect 11605 34446 20871 34448
rect 11605 34443 11671 34446
rect 20805 34443 20871 34446
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 9765 33962 9831 33965
rect 13721 33962 13787 33965
rect 9765 33960 13787 33962
rect 9765 33904 9770 33960
rect 9826 33904 13726 33960
rect 13782 33904 13787 33960
rect 9765 33902 13787 33904
rect 9765 33899 9831 33902
rect 13721 33899 13787 33902
rect 22921 33826 22987 33829
rect 23657 33826 23723 33829
rect 24117 33828 24183 33829
rect 24117 33826 24164 33828
rect 22921 33824 24164 33826
rect 22921 33768 22926 33824
rect 22982 33768 23662 33824
rect 23718 33768 24122 33824
rect 22921 33766 24164 33768
rect 22921 33763 22987 33766
rect 23657 33763 23723 33766
rect 24117 33764 24164 33766
rect 24228 33764 24234 33828
rect 24117 33763 24183 33764
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 9857 33690 9923 33693
rect 10501 33690 10567 33693
rect 17585 33690 17651 33693
rect 9857 33688 17651 33690
rect 9857 33632 9862 33688
rect 9918 33632 10506 33688
rect 10562 33632 17590 33688
rect 17646 33632 17651 33688
rect 9857 33630 17651 33632
rect 9857 33627 9923 33630
rect 10501 33627 10567 33630
rect 17585 33627 17651 33630
rect 0 33554 800 33584
rect 1301 33554 1367 33557
rect 0 33552 1367 33554
rect 0 33496 1306 33552
rect 1362 33496 1367 33552
rect 0 33494 1367 33496
rect 0 33464 800 33494
rect 1301 33491 1367 33494
rect 34329 33554 34395 33557
rect 35673 33554 36473 33584
rect 34329 33552 36473 33554
rect 34329 33496 34334 33552
rect 34390 33496 36473 33552
rect 34329 33494 36473 33496
rect 34329 33491 34395 33494
rect 35673 33464 36473 33494
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 12065 32738 12131 32741
rect 17033 32738 17099 32741
rect 12065 32736 17099 32738
rect 12065 32680 12070 32736
rect 12126 32680 17038 32736
rect 17094 32680 17099 32736
rect 12065 32678 17099 32680
rect 12065 32675 12131 32678
rect 17033 32675 17099 32678
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 27061 31786 27127 31789
rect 27889 31786 27955 31789
rect 27061 31784 27955 31786
rect 27061 31728 27066 31784
rect 27122 31728 27894 31784
rect 27950 31728 27955 31784
rect 27061 31726 27955 31728
rect 27061 31723 27127 31726
rect 27889 31723 27955 31726
rect 0 31650 800 31680
rect 1393 31650 1459 31653
rect 0 31648 1459 31650
rect 0 31592 1398 31648
rect 1454 31592 1459 31648
rect 0 31590 1459 31592
rect 0 31560 800 31590
rect 1393 31587 1459 31590
rect 34789 31650 34855 31653
rect 35673 31650 36473 31680
rect 34789 31648 36473 31650
rect 34789 31592 34794 31648
rect 34850 31592 36473 31648
rect 34789 31590 36473 31592
rect 34789 31587 34855 31590
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 35673 31560 36473 31590
rect 4870 31519 5186 31520
rect 23013 31378 23079 31381
rect 27061 31378 27127 31381
rect 23013 31376 27127 31378
rect 23013 31320 23018 31376
rect 23074 31320 27066 31376
rect 27122 31320 27127 31376
rect 23013 31318 27127 31320
rect 23013 31315 23079 31318
rect 27061 31315 27127 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 19793 30426 19859 30429
rect 27521 30426 27587 30429
rect 19793 30424 27587 30426
rect 19793 30368 19798 30424
rect 19854 30368 27526 30424
rect 27582 30368 27587 30424
rect 19793 30366 27587 30368
rect 19793 30363 19859 30366
rect 27521 30363 27587 30366
rect 11053 30290 11119 30293
rect 14273 30290 14339 30293
rect 18505 30290 18571 30293
rect 11053 30288 18571 30290
rect 11053 30232 11058 30288
rect 11114 30232 14278 30288
rect 14334 30232 18510 30288
rect 18566 30232 18571 30288
rect 11053 30230 18571 30232
rect 11053 30227 11119 30230
rect 14273 30227 14339 30230
rect 18505 30227 18571 30230
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 0 29746 800 29776
rect 1301 29746 1367 29749
rect 0 29744 1367 29746
rect 0 29688 1306 29744
rect 1362 29688 1367 29744
rect 0 29686 1367 29688
rect 0 29656 800 29686
rect 1301 29683 1367 29686
rect 34513 29746 34579 29749
rect 35673 29746 36473 29776
rect 34513 29744 36473 29746
rect 34513 29688 34518 29744
rect 34574 29688 36473 29744
rect 34513 29686 36473 29688
rect 34513 29683 34579 29686
rect 35673 29656 36473 29686
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 13445 29066 13511 29069
rect 14549 29066 14615 29069
rect 19149 29066 19215 29069
rect 26417 29068 26483 29069
rect 26366 29066 26372 29068
rect 13445 29064 19215 29066
rect 13445 29008 13450 29064
rect 13506 29008 14554 29064
rect 14610 29008 19154 29064
rect 19210 29008 19215 29064
rect 13445 29006 19215 29008
rect 26326 29006 26372 29066
rect 26436 29064 26483 29068
rect 26478 29008 26483 29064
rect 13445 29003 13511 29006
rect 14549 29003 14615 29006
rect 19149 29003 19215 29006
rect 26366 29004 26372 29006
rect 26436 29004 26483 29008
rect 26417 29003 26483 29004
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 29361 28386 29427 28389
rect 29678 28386 29684 28388
rect 29361 28384 29684 28386
rect 29361 28328 29366 28384
rect 29422 28328 29684 28384
rect 29361 28326 29684 28328
rect 29361 28323 29427 28326
rect 29678 28324 29684 28326
rect 29748 28324 29754 28388
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 4153 28114 4219 28117
rect 8937 28114 9003 28117
rect 4153 28112 9003 28114
rect 4153 28056 4158 28112
rect 4214 28056 8942 28112
rect 8998 28056 9003 28112
rect 4153 28054 9003 28056
rect 4153 28051 4219 28054
rect 8937 28051 9003 28054
rect 0 27842 800 27872
rect 1301 27842 1367 27845
rect 0 27840 1367 27842
rect 0 27784 1306 27840
rect 1362 27784 1367 27840
rect 0 27782 1367 27784
rect 0 27752 800 27782
rect 1301 27779 1367 27782
rect 35341 27842 35407 27845
rect 35673 27842 36473 27872
rect 35341 27840 36473 27842
rect 35341 27784 35346 27840
rect 35402 27784 36473 27840
rect 35341 27782 36473 27784
rect 35341 27779 35407 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 35673 27752 36473 27782
rect 34930 27711 35246 27712
rect 23565 27570 23631 27573
rect 27153 27570 27219 27573
rect 23565 27568 27219 27570
rect 23565 27512 23570 27568
rect 23626 27512 27158 27568
rect 27214 27512 27219 27568
rect 23565 27510 27219 27512
rect 23565 27507 23631 27510
rect 27153 27507 27219 27510
rect 14917 27434 14983 27437
rect 23657 27434 23723 27437
rect 14917 27432 23723 27434
rect 14917 27376 14922 27432
rect 14978 27376 23662 27432
rect 23718 27376 23723 27432
rect 14917 27374 23723 27376
rect 14917 27371 14983 27374
rect 23657 27371 23723 27374
rect 22134 27236 22140 27300
rect 22204 27298 22210 27300
rect 27981 27298 28047 27301
rect 22204 27296 28047 27298
rect 22204 27240 27986 27296
rect 28042 27240 28047 27296
rect 22204 27238 28047 27240
rect 22204 27236 22210 27238
rect 27981 27235 28047 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 10593 27026 10659 27029
rect 17769 27026 17835 27029
rect 10593 27024 17835 27026
rect 10593 26968 10598 27024
rect 10654 26968 17774 27024
rect 17830 26968 17835 27024
rect 10593 26966 17835 26968
rect 10593 26963 10659 26966
rect 17769 26963 17835 26966
rect 10501 26890 10567 26893
rect 11789 26890 11855 26893
rect 17401 26890 17467 26893
rect 18045 26890 18111 26893
rect 10501 26888 18111 26890
rect 10501 26832 10506 26888
rect 10562 26832 11794 26888
rect 11850 26832 17406 26888
rect 17462 26832 18050 26888
rect 18106 26832 18111 26888
rect 10501 26830 18111 26832
rect 10501 26827 10567 26830
rect 11789 26827 11855 26830
rect 17401 26827 17467 26830
rect 18045 26827 18111 26830
rect 20989 26890 21055 26893
rect 26601 26890 26667 26893
rect 20989 26888 26667 26890
rect 20989 26832 20994 26888
rect 21050 26832 26606 26888
rect 26662 26832 26667 26888
rect 20989 26830 26667 26832
rect 20989 26827 21055 26830
rect 26601 26827 26667 26830
rect 17217 26754 17283 26757
rect 22093 26754 22159 26757
rect 22645 26754 22711 26757
rect 17217 26752 22711 26754
rect 17217 26696 17222 26752
rect 17278 26696 22098 26752
rect 22154 26696 22650 26752
rect 22706 26696 22711 26752
rect 17217 26694 22711 26696
rect 17217 26691 17283 26694
rect 22093 26691 22159 26694
rect 22645 26691 22711 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 5717 26618 5783 26621
rect 14273 26618 14339 26621
rect 14917 26618 14983 26621
rect 5717 26616 14983 26618
rect 5717 26560 5722 26616
rect 5778 26560 14278 26616
rect 14334 26560 14922 26616
rect 14978 26560 14983 26616
rect 5717 26558 14983 26560
rect 5717 26555 5783 26558
rect 14273 26555 14339 26558
rect 14917 26555 14983 26558
rect 17125 26618 17191 26621
rect 18045 26618 18111 26621
rect 19149 26618 19215 26621
rect 17125 26616 19215 26618
rect 17125 26560 17130 26616
rect 17186 26560 18050 26616
rect 18106 26560 19154 26616
rect 19210 26560 19215 26616
rect 17125 26558 19215 26560
rect 17125 26555 17191 26558
rect 18045 26555 18111 26558
rect 19149 26555 19215 26558
rect 11697 26482 11763 26485
rect 28901 26482 28967 26485
rect 11697 26480 28967 26482
rect 11697 26424 11702 26480
rect 11758 26424 28906 26480
rect 28962 26424 28967 26480
rect 11697 26422 28967 26424
rect 11697 26419 11763 26422
rect 28901 26419 28967 26422
rect 1853 26346 1919 26349
rect 17217 26346 17283 26349
rect 1853 26344 17283 26346
rect 1853 26288 1858 26344
rect 1914 26288 17222 26344
rect 17278 26288 17283 26344
rect 1853 26286 17283 26288
rect 1853 26283 1919 26286
rect 17217 26283 17283 26286
rect 26233 26346 26299 26349
rect 27102 26346 27108 26348
rect 26233 26344 27108 26346
rect 26233 26288 26238 26344
rect 26294 26288 27108 26344
rect 26233 26286 27108 26288
rect 26233 26283 26299 26286
rect 27102 26284 27108 26286
rect 27172 26284 27178 26348
rect 24342 26148 24348 26212
rect 24412 26210 24418 26212
rect 26325 26210 26391 26213
rect 24412 26208 26391 26210
rect 24412 26152 26330 26208
rect 26386 26152 26391 26208
rect 24412 26150 26391 26152
rect 24412 26148 24418 26150
rect 26325 26147 26391 26150
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 10317 26074 10383 26077
rect 18873 26074 18939 26077
rect 10317 26072 18939 26074
rect 10317 26016 10322 26072
rect 10378 26016 18878 26072
rect 18934 26016 18939 26072
rect 10317 26014 18939 26016
rect 10317 26011 10383 26014
rect 18873 26011 18939 26014
rect 0 25938 800 25968
rect 1301 25938 1367 25941
rect 0 25936 1367 25938
rect 0 25880 1306 25936
rect 1362 25880 1367 25936
rect 0 25878 1367 25880
rect 0 25848 800 25878
rect 1301 25875 1367 25878
rect 34789 25938 34855 25941
rect 35673 25938 36473 25968
rect 34789 25936 36473 25938
rect 34789 25880 34794 25936
rect 34850 25880 36473 25936
rect 34789 25878 36473 25880
rect 34789 25875 34855 25878
rect 35673 25848 36473 25878
rect 10961 25802 11027 25805
rect 16297 25802 16363 25805
rect 10961 25800 16363 25802
rect 10961 25744 10966 25800
rect 11022 25744 16302 25800
rect 16358 25744 16363 25800
rect 10961 25742 16363 25744
rect 10961 25739 11027 25742
rect 16297 25739 16363 25742
rect 21909 25802 21975 25805
rect 22461 25802 22527 25805
rect 21909 25800 22527 25802
rect 21909 25744 21914 25800
rect 21970 25744 22466 25800
rect 22522 25744 22527 25800
rect 21909 25742 22527 25744
rect 21909 25739 21975 25742
rect 22461 25739 22527 25742
rect 27470 25604 27476 25668
rect 27540 25666 27546 25668
rect 27613 25666 27679 25669
rect 27540 25664 27679 25666
rect 27540 25608 27618 25664
rect 27674 25608 27679 25664
rect 27540 25606 27679 25608
rect 27540 25604 27546 25606
rect 27613 25603 27679 25606
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 12709 25530 12775 25533
rect 19149 25530 19215 25533
rect 12709 25528 19215 25530
rect 12709 25472 12714 25528
rect 12770 25472 19154 25528
rect 19210 25472 19215 25528
rect 12709 25470 19215 25472
rect 12709 25467 12775 25470
rect 19149 25467 19215 25470
rect 10593 25394 10659 25397
rect 10869 25394 10935 25397
rect 13629 25394 13695 25397
rect 19057 25394 19123 25397
rect 10593 25392 19123 25394
rect 10593 25336 10598 25392
rect 10654 25336 10874 25392
rect 10930 25336 13634 25392
rect 13690 25336 19062 25392
rect 19118 25336 19123 25392
rect 10593 25334 19123 25336
rect 10593 25331 10659 25334
rect 10869 25331 10935 25334
rect 13629 25331 13695 25334
rect 19057 25331 19123 25334
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 16297 24850 16363 24853
rect 17309 24850 17375 24853
rect 16297 24848 17375 24850
rect 16297 24792 16302 24848
rect 16358 24792 17314 24848
rect 17370 24792 17375 24848
rect 16297 24790 17375 24792
rect 16297 24787 16363 24790
rect 17309 24787 17375 24790
rect 13353 24714 13419 24717
rect 17217 24714 17283 24717
rect 17585 24714 17651 24717
rect 13353 24712 17651 24714
rect 13353 24656 13358 24712
rect 13414 24656 17222 24712
rect 17278 24656 17590 24712
rect 17646 24656 17651 24712
rect 13353 24654 17651 24656
rect 13353 24651 13419 24654
rect 17217 24651 17283 24654
rect 17585 24651 17651 24654
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 26417 24442 26483 24445
rect 26693 24442 26759 24445
rect 27797 24442 27863 24445
rect 28533 24442 28599 24445
rect 26417 24440 28599 24442
rect 26417 24384 26422 24440
rect 26478 24384 26698 24440
rect 26754 24384 27802 24440
rect 27858 24384 28538 24440
rect 28594 24384 28599 24440
rect 26417 24382 28599 24384
rect 26417 24379 26483 24382
rect 26693 24379 26759 24382
rect 27797 24379 27863 24382
rect 28533 24379 28599 24382
rect 21725 24306 21791 24309
rect 22461 24306 22527 24309
rect 26509 24308 26575 24309
rect 26509 24306 26556 24308
rect 21725 24304 22527 24306
rect 21725 24248 21730 24304
rect 21786 24248 22466 24304
rect 22522 24248 22527 24304
rect 21725 24246 22527 24248
rect 26464 24304 26556 24306
rect 26464 24248 26514 24304
rect 26464 24246 26556 24248
rect 21725 24243 21791 24246
rect 22461 24243 22527 24246
rect 26509 24244 26556 24246
rect 26620 24244 26626 24308
rect 26509 24243 26575 24244
rect 19149 24170 19215 24173
rect 26969 24170 27035 24173
rect 19149 24168 27035 24170
rect 19149 24112 19154 24168
rect 19210 24112 26974 24168
rect 27030 24112 27035 24168
rect 19149 24110 27035 24112
rect 19149 24107 19215 24110
rect 26969 24107 27035 24110
rect 0 24034 800 24064
rect 1209 24034 1275 24037
rect 0 24032 1275 24034
rect 0 23976 1214 24032
rect 1270 23976 1275 24032
rect 0 23974 1275 23976
rect 0 23944 800 23974
rect 1209 23971 1275 23974
rect 25865 24034 25931 24037
rect 26785 24034 26851 24037
rect 27797 24034 27863 24037
rect 28349 24034 28415 24037
rect 25865 24032 28415 24034
rect 25865 23976 25870 24032
rect 25926 23976 26790 24032
rect 26846 23976 27802 24032
rect 27858 23976 28354 24032
rect 28410 23976 28415 24032
rect 25865 23974 28415 23976
rect 25865 23971 25931 23974
rect 26785 23971 26851 23974
rect 27797 23971 27863 23974
rect 28349 23971 28415 23974
rect 34789 24034 34855 24037
rect 35673 24034 36473 24064
rect 34789 24032 36473 24034
rect 34789 23976 34794 24032
rect 34850 23976 36473 24032
rect 34789 23974 36473 23976
rect 34789 23971 34855 23974
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 35673 23944 36473 23974
rect 4870 23903 5186 23904
rect 24894 23836 24900 23900
rect 24964 23898 24970 23900
rect 26141 23898 26207 23901
rect 24964 23896 26207 23898
rect 24964 23840 26146 23896
rect 26202 23840 26207 23896
rect 24964 23838 26207 23840
rect 24964 23836 24970 23838
rect 26141 23835 26207 23838
rect 26325 23764 26391 23765
rect 26325 23762 26372 23764
rect 26280 23760 26372 23762
rect 26280 23704 26330 23760
rect 26280 23702 26372 23704
rect 26325 23700 26372 23702
rect 26436 23700 26442 23764
rect 26325 23699 26391 23700
rect 15837 23626 15903 23629
rect 27981 23626 28047 23629
rect 28717 23626 28783 23629
rect 15837 23624 28783 23626
rect 15837 23568 15842 23624
rect 15898 23568 27986 23624
rect 28042 23568 28722 23624
rect 28778 23568 28783 23624
rect 15837 23566 28783 23568
rect 15837 23563 15903 23566
rect 27981 23563 28047 23566
rect 28717 23563 28783 23566
rect 27613 23492 27679 23493
rect 27613 23488 27660 23492
rect 27724 23490 27730 23492
rect 27613 23432 27618 23488
rect 27613 23428 27660 23432
rect 27724 23430 27770 23490
rect 27724 23428 27730 23430
rect 27613 23427 27679 23428
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 1853 22538 1919 22541
rect 19241 22538 19307 22541
rect 1853 22536 19307 22538
rect 1853 22480 1858 22536
rect 1914 22480 19246 22536
rect 19302 22480 19307 22536
rect 1853 22478 19307 22480
rect 1853 22475 1919 22478
rect 19241 22475 19307 22478
rect 29729 22538 29795 22541
rect 30230 22538 30236 22540
rect 29729 22536 30236 22538
rect 29729 22480 29734 22536
rect 29790 22480 30236 22536
rect 29729 22478 30236 22480
rect 29729 22475 29795 22478
rect 30230 22476 30236 22478
rect 30300 22476 30306 22540
rect 12065 22402 12131 22405
rect 16205 22402 16271 22405
rect 12065 22400 16271 22402
rect 12065 22344 12070 22400
rect 12126 22344 16210 22400
rect 16266 22344 16271 22400
rect 12065 22342 16271 22344
rect 12065 22339 12131 22342
rect 16205 22339 16271 22342
rect 29126 22340 29132 22404
rect 29196 22402 29202 22404
rect 29269 22402 29335 22405
rect 29196 22400 29335 22402
rect 29196 22344 29274 22400
rect 29330 22344 29335 22400
rect 29196 22342 29335 22344
rect 29196 22340 29202 22342
rect 29269 22339 29335 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 0 22130 800 22160
rect 1301 22130 1367 22133
rect 28993 22130 29059 22133
rect 0 22128 1367 22130
rect 0 22072 1306 22128
rect 1362 22072 1367 22128
rect 0 22070 1367 22072
rect 0 22040 800 22070
rect 1301 22067 1367 22070
rect 28950 22128 29059 22130
rect 28950 22072 28998 22128
rect 29054 22072 29059 22128
rect 28950 22067 29059 22072
rect 34789 22130 34855 22133
rect 35673 22130 36473 22160
rect 34789 22128 36473 22130
rect 34789 22072 34794 22128
rect 34850 22072 36473 22128
rect 34789 22070 36473 22072
rect 34789 22067 34855 22070
rect 23381 21994 23447 21997
rect 27705 21994 27771 21997
rect 27889 21994 27955 21997
rect 23381 21992 27955 21994
rect 23381 21936 23386 21992
rect 23442 21936 27710 21992
rect 27766 21936 27894 21992
rect 27950 21936 27955 21992
rect 23381 21934 27955 21936
rect 23381 21931 23447 21934
rect 27705 21931 27771 21934
rect 27889 21931 27955 21934
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 28950 21722 29010 22067
rect 35673 22040 36473 22070
rect 30741 21994 30807 21997
rect 31017 21994 31083 21997
rect 30741 21992 31083 21994
rect 30741 21936 30746 21992
rect 30802 21936 31022 21992
rect 31078 21936 31083 21992
rect 30741 21934 31083 21936
rect 30741 21931 30807 21934
rect 31017 21931 31083 21934
rect 29126 21796 29132 21860
rect 29196 21858 29202 21860
rect 29269 21858 29335 21861
rect 29196 21856 29335 21858
rect 29196 21800 29274 21856
rect 29330 21800 29335 21856
rect 29196 21798 29335 21800
rect 29196 21796 29202 21798
rect 29269 21795 29335 21798
rect 29177 21722 29243 21725
rect 28950 21720 29243 21722
rect 28950 21664 29182 21720
rect 29238 21664 29243 21720
rect 28950 21662 29243 21664
rect 29177 21659 29243 21662
rect 24301 21586 24367 21589
rect 24669 21586 24735 21589
rect 24301 21584 24735 21586
rect 24301 21528 24306 21584
rect 24362 21528 24674 21584
rect 24730 21528 24735 21584
rect 24301 21526 24735 21528
rect 24301 21523 24367 21526
rect 24669 21523 24735 21526
rect 19241 21450 19307 21453
rect 26417 21450 26483 21453
rect 31017 21450 31083 21453
rect 19241 21448 31083 21450
rect 19241 21392 19246 21448
rect 19302 21392 26422 21448
rect 26478 21392 31022 21448
rect 31078 21392 31083 21448
rect 19241 21390 31083 21392
rect 19241 21387 19307 21390
rect 26417 21387 26483 21390
rect 31017 21387 31083 21390
rect 8385 21314 8451 21317
rect 19977 21314 20043 21317
rect 8385 21312 20043 21314
rect 8385 21256 8390 21312
rect 8446 21256 19982 21312
rect 20038 21256 20043 21312
rect 8385 21254 20043 21256
rect 8385 21251 8451 21254
rect 19977 21251 20043 21254
rect 30598 21252 30604 21316
rect 30668 21314 30674 21316
rect 30741 21314 30807 21317
rect 30668 21312 30807 21314
rect 30668 21256 30746 21312
rect 30802 21256 30807 21312
rect 30668 21254 30807 21256
rect 30668 21252 30674 21254
rect 30741 21251 30807 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 24117 21178 24183 21181
rect 30833 21178 30899 21181
rect 31109 21178 31175 21181
rect 24117 21176 31175 21178
rect 24117 21120 24122 21176
rect 24178 21120 30838 21176
rect 30894 21120 31114 21176
rect 31170 21120 31175 21176
rect 24117 21118 31175 21120
rect 24117 21115 24183 21118
rect 30833 21115 30899 21118
rect 31109 21115 31175 21118
rect 20529 20906 20595 20909
rect 28349 20906 28415 20909
rect 20529 20904 28415 20906
rect 20529 20848 20534 20904
rect 20590 20848 28354 20904
rect 28410 20848 28415 20904
rect 20529 20846 28415 20848
rect 20529 20843 20595 20846
rect 28349 20843 28415 20846
rect 28758 20708 28764 20772
rect 28828 20770 28834 20772
rect 29126 20770 29132 20772
rect 28828 20710 29132 20770
rect 28828 20708 28834 20710
rect 29126 20708 29132 20710
rect 29196 20708 29202 20772
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 22093 20636 22159 20637
rect 22093 20632 22140 20636
rect 22204 20634 22210 20636
rect 22093 20576 22098 20632
rect 22093 20572 22140 20576
rect 22204 20574 22250 20634
rect 22204 20572 22210 20574
rect 22093 20571 22159 20572
rect 22461 20498 22527 20501
rect 25313 20498 25379 20501
rect 22461 20496 25379 20498
rect 22461 20440 22466 20496
rect 22522 20440 25318 20496
rect 25374 20440 25379 20496
rect 22461 20438 25379 20440
rect 22461 20435 22527 20438
rect 25313 20435 25379 20438
rect 24393 20362 24459 20365
rect 26785 20362 26851 20365
rect 24393 20360 26851 20362
rect 24393 20304 24398 20360
rect 24454 20304 26790 20360
rect 26846 20304 26851 20360
rect 24393 20302 26851 20304
rect 24393 20299 24459 20302
rect 26785 20299 26851 20302
rect 0 20226 800 20256
rect 1301 20226 1367 20229
rect 0 20224 1367 20226
rect 0 20168 1306 20224
rect 1362 20168 1367 20224
rect 0 20166 1367 20168
rect 0 20136 800 20166
rect 1301 20163 1367 20166
rect 20989 20226 21055 20229
rect 26601 20226 26667 20229
rect 20989 20224 26667 20226
rect 20989 20168 20994 20224
rect 21050 20168 26606 20224
rect 26662 20168 26667 20224
rect 20989 20166 26667 20168
rect 20989 20163 21055 20166
rect 26601 20163 26667 20166
rect 35341 20226 35407 20229
rect 35673 20226 36473 20256
rect 35341 20224 36473 20226
rect 35341 20168 35346 20224
rect 35402 20168 36473 20224
rect 35341 20166 36473 20168
rect 35341 20163 35407 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 35673 20136 36473 20166
rect 34930 20095 35246 20096
rect 24853 20092 24919 20093
rect 24853 20090 24900 20092
rect 24808 20088 24900 20090
rect 24808 20032 24858 20088
rect 24808 20030 24900 20032
rect 24853 20028 24900 20030
rect 24964 20028 24970 20092
rect 24853 20027 24919 20028
rect 10409 19682 10475 19685
rect 15653 19682 15719 19685
rect 23197 19684 23263 19685
rect 23197 19682 23244 19684
rect 10409 19680 15719 19682
rect 10409 19624 10414 19680
rect 10470 19624 15658 19680
rect 15714 19624 15719 19680
rect 10409 19622 15719 19624
rect 23152 19680 23244 19682
rect 23152 19624 23202 19680
rect 23152 19622 23244 19624
rect 10409 19619 10475 19622
rect 15653 19619 15719 19622
rect 23197 19620 23244 19622
rect 23308 19620 23314 19684
rect 23197 19619 23263 19620
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 10777 19410 10843 19413
rect 12433 19410 12499 19413
rect 10777 19408 12499 19410
rect 10777 19352 10782 19408
rect 10838 19352 12438 19408
rect 12494 19352 12499 19408
rect 10777 19350 12499 19352
rect 10777 19347 10843 19350
rect 12433 19347 12499 19350
rect 25957 19410 26023 19413
rect 26182 19410 26188 19412
rect 25957 19408 26188 19410
rect 25957 19352 25962 19408
rect 26018 19352 26188 19408
rect 25957 19350 26188 19352
rect 25957 19347 26023 19350
rect 26182 19348 26188 19350
rect 26252 19348 26258 19412
rect 26509 19410 26575 19413
rect 27429 19410 27495 19413
rect 26509 19408 27495 19410
rect 26509 19352 26514 19408
rect 26570 19352 27434 19408
rect 27490 19352 27495 19408
rect 26509 19350 27495 19352
rect 26509 19347 26575 19350
rect 27429 19347 27495 19350
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 21817 19002 21883 19005
rect 24577 19002 24643 19005
rect 21817 19000 24643 19002
rect 21817 18944 21822 19000
rect 21878 18944 24582 19000
rect 24638 18944 24643 19000
rect 21817 18942 24643 18944
rect 21817 18939 21883 18942
rect 24577 18939 24643 18942
rect 17677 18730 17743 18733
rect 34145 18730 34211 18733
rect 17677 18728 34211 18730
rect 17677 18672 17682 18728
rect 17738 18672 34150 18728
rect 34206 18672 34211 18728
rect 17677 18670 34211 18672
rect 17677 18667 17743 18670
rect 34145 18667 34211 18670
rect 21541 18594 21607 18597
rect 24342 18594 24348 18596
rect 21541 18592 24348 18594
rect 21541 18536 21546 18592
rect 21602 18536 24348 18592
rect 21541 18534 24348 18536
rect 21541 18531 21607 18534
rect 24342 18532 24348 18534
rect 24412 18532 24418 18596
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 0 18322 800 18352
rect 1301 18322 1367 18325
rect 0 18320 1367 18322
rect 0 18264 1306 18320
rect 1362 18264 1367 18320
rect 0 18262 1367 18264
rect 0 18232 800 18262
rect 1301 18259 1367 18262
rect 22093 18322 22159 18325
rect 23933 18322 23999 18325
rect 22093 18320 23999 18322
rect 22093 18264 22098 18320
rect 22154 18264 23938 18320
rect 23994 18264 23999 18320
rect 22093 18262 23999 18264
rect 22093 18259 22159 18262
rect 23933 18259 23999 18262
rect 25313 18322 25379 18325
rect 25681 18322 25747 18325
rect 25313 18320 25747 18322
rect 25313 18264 25318 18320
rect 25374 18264 25686 18320
rect 25742 18264 25747 18320
rect 25313 18262 25747 18264
rect 25313 18259 25379 18262
rect 25681 18259 25747 18262
rect 34789 18322 34855 18325
rect 35673 18322 36473 18352
rect 34789 18320 36473 18322
rect 34789 18264 34794 18320
rect 34850 18264 36473 18320
rect 34789 18262 36473 18264
rect 34789 18259 34855 18262
rect 35673 18232 36473 18262
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 25957 17914 26023 17917
rect 27654 17914 27660 17916
rect 25957 17912 27660 17914
rect 25957 17856 25962 17912
rect 26018 17856 27660 17912
rect 25957 17854 27660 17856
rect 25957 17851 26023 17854
rect 27654 17852 27660 17854
rect 27724 17852 27730 17916
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 14733 16826 14799 16829
rect 14733 16824 15210 16826
rect 14733 16768 14738 16824
rect 14794 16768 15210 16824
rect 14733 16766 15210 16768
rect 14733 16763 14799 16766
rect 15150 16690 15210 16766
rect 15285 16690 15351 16693
rect 15510 16690 15516 16692
rect 15150 16688 15516 16690
rect 15150 16632 15290 16688
rect 15346 16632 15516 16688
rect 15150 16630 15516 16632
rect 15285 16627 15351 16630
rect 15510 16628 15516 16630
rect 15580 16628 15586 16692
rect 26918 16628 26924 16692
rect 26988 16690 26994 16692
rect 27061 16690 27127 16693
rect 26988 16688 27127 16690
rect 26988 16632 27066 16688
rect 27122 16632 27127 16688
rect 26988 16630 27127 16632
rect 26988 16628 26994 16630
rect 27061 16627 27127 16630
rect 17217 16554 17283 16557
rect 24158 16554 24164 16556
rect 17217 16552 24164 16554
rect 17217 16496 17222 16552
rect 17278 16496 24164 16552
rect 17217 16494 24164 16496
rect 17217 16491 17283 16494
rect 24158 16492 24164 16494
rect 24228 16554 24234 16556
rect 30005 16554 30071 16557
rect 24228 16552 30071 16554
rect 24228 16496 30010 16552
rect 30066 16496 30071 16552
rect 24228 16494 30071 16496
rect 24228 16492 24234 16494
rect 30005 16491 30071 16494
rect 0 16418 800 16448
rect 1393 16418 1459 16421
rect 0 16416 1459 16418
rect 0 16360 1398 16416
rect 1454 16360 1459 16416
rect 0 16358 1459 16360
rect 0 16328 800 16358
rect 1393 16355 1459 16358
rect 26182 16356 26188 16420
rect 26252 16418 26258 16420
rect 27337 16418 27403 16421
rect 26252 16416 27403 16418
rect 26252 16360 27342 16416
rect 27398 16360 27403 16416
rect 26252 16358 27403 16360
rect 26252 16356 26258 16358
rect 27337 16355 27403 16358
rect 34329 16418 34395 16421
rect 35673 16418 36473 16448
rect 34329 16416 36473 16418
rect 34329 16360 34334 16416
rect 34390 16360 36473 16416
rect 34329 16358 36473 16360
rect 34329 16355 34395 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 35673 16328 36473 16358
rect 4870 16287 5186 16288
rect 22185 16148 22251 16149
rect 22134 16084 22140 16148
rect 22204 16146 22251 16148
rect 22204 16144 22296 16146
rect 22246 16088 22296 16144
rect 22204 16086 22296 16088
rect 22204 16084 22251 16086
rect 22185 16083 22251 16084
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 22461 15602 22527 15605
rect 23054 15602 23060 15604
rect 22461 15600 23060 15602
rect 22461 15544 22466 15600
rect 22522 15544 23060 15600
rect 22461 15542 23060 15544
rect 22461 15539 22527 15542
rect 23054 15540 23060 15542
rect 23124 15540 23130 15604
rect 9029 15330 9095 15333
rect 13169 15330 13235 15333
rect 9029 15328 13235 15330
rect 9029 15272 9034 15328
rect 9090 15272 13174 15328
rect 13230 15272 13235 15328
rect 9029 15270 13235 15272
rect 9029 15267 9095 15270
rect 13169 15267 13235 15270
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 30230 15132 30236 15196
rect 30300 15194 30306 15196
rect 30557 15194 30623 15197
rect 30300 15192 30623 15194
rect 30300 15136 30562 15192
rect 30618 15136 30623 15192
rect 30300 15134 30623 15136
rect 30300 15132 30306 15134
rect 30557 15131 30623 15134
rect 26877 15060 26943 15061
rect 26877 15058 26924 15060
rect 26832 15056 26924 15058
rect 26832 15000 26882 15056
rect 26832 14998 26924 15000
rect 26877 14996 26924 14998
rect 26988 14996 26994 15060
rect 26877 14995 26943 14996
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 21725 14650 21791 14653
rect 28717 14650 28783 14653
rect 21725 14648 28783 14650
rect 21725 14592 21730 14648
rect 21786 14592 28722 14648
rect 28778 14592 28783 14648
rect 21725 14590 28783 14592
rect 21725 14587 21791 14590
rect 28717 14587 28783 14590
rect 0 14514 800 14544
rect 1301 14514 1367 14517
rect 0 14512 1367 14514
rect 0 14456 1306 14512
rect 1362 14456 1367 14512
rect 0 14454 1367 14456
rect 0 14424 800 14454
rect 1301 14451 1367 14454
rect 34697 14514 34763 14517
rect 35673 14514 36473 14544
rect 34697 14512 36473 14514
rect 34697 14456 34702 14512
rect 34758 14456 36473 14512
rect 34697 14454 36473 14456
rect 34697 14451 34763 14454
rect 35673 14424 36473 14454
rect 15510 14316 15516 14380
rect 15580 14378 15586 14380
rect 27889 14378 27955 14381
rect 28809 14378 28875 14381
rect 15580 14376 28875 14378
rect 15580 14320 27894 14376
rect 27950 14320 28814 14376
rect 28870 14320 28875 14376
rect 15580 14318 28875 14320
rect 15580 14316 15586 14318
rect 27889 14315 27955 14318
rect 28809 14315 28875 14318
rect 27705 14242 27771 14245
rect 28625 14242 28691 14245
rect 27705 14240 28691 14242
rect 27705 14184 27710 14240
rect 27766 14184 28630 14240
rect 28686 14184 28691 14240
rect 27705 14182 28691 14184
rect 27705 14179 27771 14182
rect 28625 14179 28691 14182
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 27061 14108 27127 14109
rect 27061 14106 27108 14108
rect 27016 14104 27108 14106
rect 27016 14048 27066 14104
rect 27016 14046 27108 14048
rect 27061 14044 27108 14046
rect 27172 14044 27178 14108
rect 27061 14043 27127 14044
rect 16021 13698 16087 13701
rect 16389 13698 16455 13701
rect 16021 13696 16455 13698
rect 16021 13640 16026 13696
rect 16082 13640 16394 13696
rect 16450 13640 16455 13696
rect 16021 13638 16455 13640
rect 16021 13635 16087 13638
rect 16389 13635 16455 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 11789 13426 11855 13429
rect 27337 13426 27403 13429
rect 11789 13424 27403 13426
rect 11789 13368 11794 13424
rect 11850 13368 27342 13424
rect 27398 13368 27403 13424
rect 11789 13366 27403 13368
rect 11789 13363 11855 13366
rect 27337 13363 27403 13366
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 12617 13018 12683 13021
rect 19057 13018 19123 13021
rect 12617 13016 19123 13018
rect 12617 12960 12622 13016
rect 12678 12960 19062 13016
rect 19118 12960 19123 13016
rect 12617 12958 19123 12960
rect 12617 12955 12683 12958
rect 19057 12955 19123 12958
rect 17585 12882 17651 12885
rect 28165 12882 28231 12885
rect 17585 12880 28231 12882
rect 17585 12824 17590 12880
rect 17646 12824 28170 12880
rect 28226 12824 28231 12880
rect 17585 12822 28231 12824
rect 17585 12819 17651 12822
rect 28165 12819 28231 12822
rect 14641 12746 14707 12749
rect 23381 12746 23447 12749
rect 14641 12744 23447 12746
rect 14641 12688 14646 12744
rect 14702 12688 23386 12744
rect 23442 12688 23447 12744
rect 14641 12686 23447 12688
rect 14641 12683 14707 12686
rect 23381 12683 23447 12686
rect 0 12610 800 12640
rect 1301 12610 1367 12613
rect 0 12608 1367 12610
rect 0 12552 1306 12608
rect 1362 12552 1367 12608
rect 0 12550 1367 12552
rect 0 12520 800 12550
rect 1301 12547 1367 12550
rect 19149 12610 19215 12613
rect 19701 12610 19767 12613
rect 19149 12608 19767 12610
rect 19149 12552 19154 12608
rect 19210 12552 19706 12608
rect 19762 12552 19767 12608
rect 19149 12550 19767 12552
rect 19149 12547 19215 12550
rect 19701 12547 19767 12550
rect 35341 12610 35407 12613
rect 35673 12610 36473 12640
rect 35341 12608 36473 12610
rect 35341 12552 35346 12608
rect 35402 12552 36473 12608
rect 35341 12550 36473 12552
rect 35341 12547 35407 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 35673 12520 36473 12550
rect 34930 12479 35246 12480
rect 26141 12474 26207 12477
rect 25270 12472 26207 12474
rect 25270 12416 26146 12472
rect 26202 12416 26207 12472
rect 25270 12414 26207 12416
rect 19333 12338 19399 12341
rect 25270 12338 25330 12414
rect 26141 12411 26207 12414
rect 19333 12336 25330 12338
rect 19333 12280 19338 12336
rect 19394 12280 25330 12336
rect 19333 12278 25330 12280
rect 19333 12275 19399 12278
rect 24025 12202 24091 12205
rect 24342 12202 24348 12204
rect 24025 12200 24348 12202
rect 24025 12144 24030 12200
rect 24086 12144 24348 12200
rect 24025 12142 24348 12144
rect 24025 12139 24091 12142
rect 24342 12140 24348 12142
rect 24412 12140 24418 12204
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 15142 11596 15148 11660
rect 15212 11658 15218 11660
rect 16665 11658 16731 11661
rect 15212 11656 16731 11658
rect 15212 11600 16670 11656
rect 16726 11600 16731 11656
rect 15212 11598 16731 11600
rect 15212 11596 15218 11598
rect 16665 11595 16731 11598
rect 17585 11658 17651 11661
rect 23238 11658 23244 11660
rect 17585 11656 23244 11658
rect 17585 11600 17590 11656
rect 17646 11600 23244 11656
rect 17585 11598 23244 11600
rect 17585 11595 17651 11598
rect 23238 11596 23244 11598
rect 23308 11658 23314 11660
rect 28257 11658 28323 11661
rect 23308 11656 28323 11658
rect 23308 11600 28262 11656
rect 28318 11600 28323 11656
rect 23308 11598 28323 11600
rect 23308 11596 23314 11598
rect 28257 11595 28323 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19517 11250 19583 11253
rect 34145 11250 34211 11253
rect 19517 11248 34211 11250
rect 19517 11192 19522 11248
rect 19578 11192 34150 11248
rect 34206 11192 34211 11248
rect 19517 11190 34211 11192
rect 19517 11187 19583 11190
rect 34145 11187 34211 11190
rect 5073 11114 5139 11117
rect 11973 11114 12039 11117
rect 19609 11114 19675 11117
rect 5073 11112 19675 11114
rect 5073 11056 5078 11112
rect 5134 11056 11978 11112
rect 12034 11056 19614 11112
rect 19670 11056 19675 11112
rect 5073 11054 19675 11056
rect 5073 11051 5139 11054
rect 11973 11051 12039 11054
rect 19609 11051 19675 11054
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 23105 10842 23171 10845
rect 28257 10842 28323 10845
rect 23105 10840 28323 10842
rect 23105 10784 23110 10840
rect 23166 10784 28262 10840
rect 28318 10784 28323 10840
rect 23105 10782 28323 10784
rect 23105 10779 23171 10782
rect 28257 10779 28323 10782
rect 0 10706 800 10736
rect 1301 10706 1367 10709
rect 0 10704 1367 10706
rect 0 10648 1306 10704
rect 1362 10648 1367 10704
rect 0 10646 1367 10648
rect 0 10616 800 10646
rect 1301 10643 1367 10646
rect 3141 10706 3207 10709
rect 5901 10706 5967 10709
rect 3141 10704 5967 10706
rect 3141 10648 3146 10704
rect 3202 10648 5906 10704
rect 5962 10648 5967 10704
rect 3141 10646 5967 10648
rect 3141 10643 3207 10646
rect 5901 10643 5967 10646
rect 12433 10706 12499 10709
rect 17125 10706 17191 10709
rect 12433 10704 17191 10706
rect 12433 10648 12438 10704
rect 12494 10648 17130 10704
rect 17186 10648 17191 10704
rect 12433 10646 17191 10648
rect 12433 10643 12499 10646
rect 17125 10643 17191 10646
rect 18321 10706 18387 10709
rect 29545 10706 29611 10709
rect 18321 10704 29611 10706
rect 18321 10648 18326 10704
rect 18382 10648 29550 10704
rect 29606 10648 29611 10704
rect 18321 10646 29611 10648
rect 18321 10643 18387 10646
rect 29545 10643 29611 10646
rect 34789 10706 34855 10709
rect 35673 10706 36473 10736
rect 34789 10704 36473 10706
rect 34789 10648 34794 10704
rect 34850 10648 36473 10704
rect 34789 10646 36473 10648
rect 34789 10643 34855 10646
rect 35673 10616 36473 10646
rect 22921 10570 22987 10573
rect 26693 10570 26759 10573
rect 22921 10568 26759 10570
rect 22921 10512 22926 10568
rect 22982 10512 26698 10568
rect 26754 10512 26759 10568
rect 22921 10510 26759 10512
rect 22921 10507 22987 10510
rect 26693 10507 26759 10510
rect 27153 10434 27219 10437
rect 28717 10434 28783 10437
rect 27153 10432 28783 10434
rect 27153 10376 27158 10432
rect 27214 10376 28722 10432
rect 28778 10376 28783 10432
rect 27153 10374 28783 10376
rect 27153 10371 27219 10374
rect 28717 10371 28783 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 28809 10164 28875 10165
rect 28758 10100 28764 10164
rect 28828 10162 28875 10164
rect 29637 10164 29703 10165
rect 29637 10162 29684 10164
rect 28828 10160 28920 10162
rect 28870 10104 28920 10160
rect 28828 10102 28920 10104
rect 29592 10160 29684 10162
rect 29592 10104 29642 10160
rect 29592 10102 29684 10104
rect 28828 10100 28875 10102
rect 28809 10099 28875 10100
rect 29637 10100 29684 10102
rect 29748 10100 29754 10164
rect 29637 10099 29703 10100
rect 9765 10026 9831 10029
rect 16941 10026 17007 10029
rect 9765 10024 17007 10026
rect 9765 9968 9770 10024
rect 9826 9968 16946 10024
rect 17002 9968 17007 10024
rect 9765 9966 17007 9968
rect 9765 9963 9831 9966
rect 16941 9963 17007 9966
rect 30465 10026 30531 10029
rect 30598 10026 30604 10028
rect 30465 10024 30604 10026
rect 30465 9968 30470 10024
rect 30526 9968 30604 10024
rect 30465 9966 30604 9968
rect 30465 9963 30531 9966
rect 30598 9964 30604 9966
rect 30668 9964 30674 10028
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 5349 9618 5415 9621
rect 6085 9618 6151 9621
rect 5349 9616 6151 9618
rect 5349 9560 5354 9616
rect 5410 9560 6090 9616
rect 6146 9560 6151 9616
rect 5349 9558 6151 9560
rect 5349 9555 5415 9558
rect 6085 9555 6151 9558
rect 20345 9618 20411 9621
rect 22645 9618 22711 9621
rect 20345 9616 22711 9618
rect 20345 9560 20350 9616
rect 20406 9560 22650 9616
rect 22706 9560 22711 9616
rect 20345 9558 22711 9560
rect 20345 9555 20411 9558
rect 22645 9555 22711 9558
rect 23054 9556 23060 9620
rect 23124 9618 23130 9620
rect 26509 9618 26575 9621
rect 23124 9616 26575 9618
rect 23124 9560 26514 9616
rect 26570 9560 26575 9616
rect 23124 9558 26575 9560
rect 23124 9556 23130 9558
rect 26509 9555 26575 9558
rect 22461 9482 22527 9485
rect 26325 9482 26391 9485
rect 22461 9480 26391 9482
rect 22461 9424 22466 9480
rect 22522 9424 26330 9480
rect 26386 9424 26391 9480
rect 22461 9422 26391 9424
rect 22461 9419 22527 9422
rect 26325 9419 26391 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 21357 9210 21423 9213
rect 28441 9210 28507 9213
rect 21357 9208 28507 9210
rect 21357 9152 21362 9208
rect 21418 9152 28446 9208
rect 28502 9152 28507 9208
rect 21357 9150 28507 9152
rect 21357 9147 21423 9150
rect 28441 9147 28507 9150
rect 20621 9074 20687 9077
rect 22001 9074 22067 9077
rect 20621 9072 22067 9074
rect 20621 9016 20626 9072
rect 20682 9016 22006 9072
rect 22062 9016 22067 9072
rect 20621 9014 22067 9016
rect 20621 9011 20687 9014
rect 22001 9011 22067 9014
rect 22737 9074 22803 9077
rect 31753 9074 31819 9077
rect 22737 9072 31819 9074
rect 22737 9016 22742 9072
rect 22798 9016 31758 9072
rect 31814 9016 31819 9072
rect 22737 9014 31819 9016
rect 22737 9011 22803 9014
rect 31753 9011 31819 9014
rect 6821 8938 6887 8941
rect 29729 8938 29795 8941
rect 6821 8936 29795 8938
rect 6821 8880 6826 8936
rect 6882 8880 29734 8936
rect 29790 8880 29795 8936
rect 6821 8878 29795 8880
rect 6821 8875 6887 8878
rect 29729 8875 29795 8878
rect 0 8802 800 8832
rect 1301 8802 1367 8805
rect 0 8800 1367 8802
rect 0 8744 1306 8800
rect 1362 8744 1367 8800
rect 0 8742 1367 8744
rect 0 8712 800 8742
rect 1301 8739 1367 8742
rect 22277 8802 22343 8805
rect 34053 8802 34119 8805
rect 22277 8800 34119 8802
rect 22277 8744 22282 8800
rect 22338 8744 34058 8800
rect 34114 8744 34119 8800
rect 22277 8742 34119 8744
rect 22277 8739 22343 8742
rect 34053 8739 34119 8742
rect 34789 8802 34855 8805
rect 35673 8802 36473 8832
rect 34789 8800 36473 8802
rect 34789 8744 34794 8800
rect 34850 8744 36473 8800
rect 34789 8742 36473 8744
rect 34789 8739 34855 8742
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 35673 8712 36473 8742
rect 4870 8671 5186 8672
rect 21633 8666 21699 8669
rect 22461 8666 22527 8669
rect 21633 8664 22527 8666
rect 21633 8608 21638 8664
rect 21694 8608 22466 8664
rect 22522 8608 22527 8664
rect 21633 8606 22527 8608
rect 21633 8603 21699 8606
rect 22461 8603 22527 8606
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6898 800 6928
rect 1301 6898 1367 6901
rect 0 6896 1367 6898
rect 0 6840 1306 6896
rect 1362 6840 1367 6896
rect 0 6838 1367 6840
rect 0 6808 800 6838
rect 1301 6835 1367 6838
rect 12433 6898 12499 6901
rect 15142 6898 15148 6900
rect 12433 6896 15148 6898
rect 12433 6840 12438 6896
rect 12494 6840 15148 6896
rect 12433 6838 15148 6840
rect 12433 6835 12499 6838
rect 15142 6836 15148 6838
rect 15212 6836 15218 6900
rect 18597 6898 18663 6901
rect 34053 6898 34119 6901
rect 18597 6896 34119 6898
rect 18597 6840 18602 6896
rect 18658 6840 34058 6896
rect 34114 6840 34119 6896
rect 18597 6838 34119 6840
rect 18597 6835 18663 6838
rect 34053 6835 34119 6838
rect 34697 6898 34763 6901
rect 35673 6898 36473 6928
rect 34697 6896 36473 6898
rect 34697 6840 34702 6896
rect 34758 6840 36473 6896
rect 34697 6838 36473 6840
rect 34697 6835 34763 6838
rect 35673 6808 36473 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 29637 6218 29703 6221
rect 32857 6218 32923 6221
rect 29637 6216 32923 6218
rect 29637 6160 29642 6216
rect 29698 6160 32862 6216
rect 32918 6160 32923 6216
rect 29637 6158 32923 6160
rect 29637 6155 29703 6158
rect 32857 6155 32923 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 30833 5810 30899 5813
rect 31661 5810 31727 5813
rect 30833 5808 31727 5810
rect 30833 5752 30838 5808
rect 30894 5752 31666 5808
rect 31722 5752 31727 5808
rect 30833 5750 31727 5752
rect 30833 5747 30899 5750
rect 31661 5747 31727 5750
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 0 4994 800 5024
rect 1301 4994 1367 4997
rect 0 4992 1367 4994
rect 0 4936 1306 4992
rect 1362 4936 1367 4992
rect 0 4934 1367 4936
rect 0 4904 800 4934
rect 1301 4931 1367 4934
rect 35341 4994 35407 4997
rect 35673 4994 36473 5024
rect 35341 4992 36473 4994
rect 35341 4936 35346 4992
rect 35402 4936 36473 4992
rect 35341 4934 36473 4936
rect 35341 4931 35407 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 35673 4904 36473 4934
rect 34930 4863 35246 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 0 3090 800 3120
rect 1301 3090 1367 3093
rect 0 3088 1367 3090
rect 0 3032 1306 3088
rect 1362 3032 1367 3088
rect 0 3030 1367 3032
rect 0 3000 800 3030
rect 1301 3027 1367 3030
rect 34329 3090 34395 3093
rect 35673 3090 36473 3120
rect 34329 3088 36473 3090
rect 34329 3032 34334 3088
rect 34390 3032 36473 3088
rect 34329 3030 36473 3032
rect 34329 3027 34395 3030
rect 35673 3000 36473 3030
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 0 1186 800 1216
rect 18137 1186 18203 1189
rect 0 1184 18203 1186
rect 0 1128 18142 1184
rect 18198 1128 18203 1184
rect 0 1126 18203 1128
rect 0 1096 800 1126
rect 18137 1123 18203 1126
<< via3 >>
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 27476 35456 27540 35460
rect 27476 35400 27490 35456
rect 27490 35400 27540 35456
rect 27476 35396 27540 35400
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 26556 35124 26620 35188
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 24164 33824 24228 33828
rect 24164 33768 24178 33824
rect 24178 33768 24228 33824
rect 24164 33764 24228 33768
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 26372 29064 26436 29068
rect 26372 29008 26422 29064
rect 26422 29008 26436 29064
rect 26372 29004 26436 29008
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 29684 28324 29748 28388
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 22140 27236 22204 27300
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 27108 26284 27172 26348
rect 24348 26148 24412 26212
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 27476 25604 27540 25668
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 26556 24304 26620 24308
rect 26556 24248 26570 24304
rect 26570 24248 26620 24304
rect 26556 24244 26620 24248
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 24900 23836 24964 23900
rect 26372 23760 26436 23764
rect 26372 23704 26386 23760
rect 26386 23704 26436 23760
rect 26372 23700 26436 23704
rect 27660 23488 27724 23492
rect 27660 23432 27674 23488
rect 27674 23432 27724 23488
rect 27660 23428 27724 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 30236 22476 30300 22540
rect 29132 22340 29196 22404
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 29132 21796 29196 21860
rect 30604 21252 30668 21316
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 28764 20708 28828 20772
rect 29132 20708 29196 20772
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 22140 20632 22204 20636
rect 22140 20576 22154 20632
rect 22154 20576 22204 20632
rect 22140 20572 22204 20576
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 24900 20088 24964 20092
rect 24900 20032 24914 20088
rect 24914 20032 24964 20088
rect 24900 20028 24964 20032
rect 23244 19680 23308 19684
rect 23244 19624 23258 19680
rect 23258 19624 23308 19680
rect 23244 19620 23308 19624
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 26188 19348 26252 19412
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 24348 18532 24412 18596
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 27660 17852 27724 17916
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 15516 16628 15580 16692
rect 26924 16628 26988 16692
rect 24164 16492 24228 16556
rect 26188 16356 26252 16420
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 22140 16144 22204 16148
rect 22140 16088 22190 16144
rect 22190 16088 22204 16144
rect 22140 16084 22204 16088
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 23060 15540 23124 15604
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 30236 15132 30300 15196
rect 26924 15056 26988 15060
rect 26924 15000 26938 15056
rect 26938 15000 26988 15056
rect 26924 14996 26988 15000
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 15516 14316 15580 14380
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 27108 14104 27172 14108
rect 27108 14048 27122 14104
rect 27122 14048 27172 14104
rect 27108 14044 27172 14048
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 24348 12140 24412 12204
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 15148 11596 15212 11660
rect 23244 11596 23308 11660
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 28764 10160 28828 10164
rect 28764 10104 28814 10160
rect 28814 10104 28828 10160
rect 28764 10100 28828 10104
rect 29684 10160 29748 10164
rect 29684 10104 29698 10160
rect 29698 10104 29748 10160
rect 29684 10100 29748 10104
rect 30604 9964 30668 10028
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 23060 9556 23124 9620
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 15148 6836 15212 6900
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 35392 4528 35952
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 35936 5188 35952
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 27475 35460 27541 35461
rect 27475 35396 27476 35460
rect 27540 35396 27541 35460
rect 27475 35395 27541 35396
rect 26555 35188 26621 35189
rect 26555 35124 26556 35188
rect 26620 35124 26621 35188
rect 26555 35123 26621 35124
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 24163 33828 24229 33829
rect 24163 33764 24164 33828
rect 24228 33764 24229 33828
rect 24163 33763 24229 33764
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 22139 27300 22205 27301
rect 22139 27236 22140 27300
rect 22204 27236 22205 27300
rect 22139 27235 22205 27236
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 22142 20637 22202 27235
rect 22139 20636 22205 20637
rect 22139 20572 22140 20636
rect 22204 20572 22205 20636
rect 22139 20571 22205 20572
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 15515 16692 15581 16693
rect 15515 16628 15516 16692
rect 15580 16628 15581 16692
rect 15515 16627 15581 16628
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 15518 14381 15578 16627
rect 22142 16149 22202 20571
rect 23243 19684 23309 19685
rect 23243 19620 23244 19684
rect 23308 19620 23309 19684
rect 23243 19619 23309 19620
rect 22139 16148 22205 16149
rect 22139 16084 22140 16148
rect 22204 16084 22205 16148
rect 22139 16083 22205 16084
rect 23059 15604 23125 15605
rect 23059 15540 23060 15604
rect 23124 15540 23125 15604
rect 23059 15539 23125 15540
rect 15515 14380 15581 14381
rect 15515 14316 15516 14380
rect 15580 14316 15581 14380
rect 15515 14315 15581 14316
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 15147 11660 15213 11661
rect 15147 11596 15148 11660
rect 15212 11596 15213 11660
rect 15147 11595 15213 11596
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 15150 6901 15210 11595
rect 23062 9621 23122 15539
rect 23246 11661 23306 19619
rect 24166 16557 24226 33763
rect 26371 29068 26437 29069
rect 26371 29004 26372 29068
rect 26436 29004 26437 29068
rect 26371 29003 26437 29004
rect 24347 26212 24413 26213
rect 24347 26148 24348 26212
rect 24412 26148 24413 26212
rect 24347 26147 24413 26148
rect 24350 18597 24410 26147
rect 24899 23900 24965 23901
rect 24899 23836 24900 23900
rect 24964 23836 24965 23900
rect 24899 23835 24965 23836
rect 24902 20093 24962 23835
rect 26374 23765 26434 29003
rect 26558 24309 26618 35123
rect 27107 26348 27173 26349
rect 27107 26284 27108 26348
rect 27172 26284 27173 26348
rect 27107 26283 27173 26284
rect 26555 24308 26621 24309
rect 26555 24244 26556 24308
rect 26620 24244 26621 24308
rect 26555 24243 26621 24244
rect 26371 23764 26437 23765
rect 26371 23700 26372 23764
rect 26436 23700 26437 23764
rect 26371 23699 26437 23700
rect 24899 20092 24965 20093
rect 24899 20028 24900 20092
rect 24964 20028 24965 20092
rect 24899 20027 24965 20028
rect 26187 19412 26253 19413
rect 26187 19348 26188 19412
rect 26252 19348 26253 19412
rect 26187 19347 26253 19348
rect 24347 18596 24413 18597
rect 24347 18532 24348 18596
rect 24412 18532 24413 18596
rect 24347 18531 24413 18532
rect 24163 16556 24229 16557
rect 24163 16492 24164 16556
rect 24228 16492 24229 16556
rect 24163 16491 24229 16492
rect 24350 12205 24410 18531
rect 26190 16421 26250 19347
rect 26923 16692 26989 16693
rect 26923 16628 26924 16692
rect 26988 16628 26989 16692
rect 26923 16627 26989 16628
rect 26187 16420 26253 16421
rect 26187 16356 26188 16420
rect 26252 16356 26253 16420
rect 26187 16355 26253 16356
rect 26926 15061 26986 16627
rect 26923 15060 26989 15061
rect 26923 14996 26924 15060
rect 26988 14996 26989 15060
rect 26923 14995 26989 14996
rect 27110 14109 27170 26283
rect 27478 25669 27538 35395
rect 34928 35392 35248 35952
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 29683 28388 29749 28389
rect 29683 28324 29684 28388
rect 29748 28324 29749 28388
rect 29683 28323 29749 28324
rect 27475 25668 27541 25669
rect 27475 25604 27476 25668
rect 27540 25604 27541 25668
rect 27475 25603 27541 25604
rect 27659 23492 27725 23493
rect 27659 23428 27660 23492
rect 27724 23428 27725 23492
rect 27659 23427 27725 23428
rect 27662 17917 27722 23427
rect 29131 22404 29197 22405
rect 29131 22340 29132 22404
rect 29196 22340 29197 22404
rect 29131 22339 29197 22340
rect 29134 21861 29194 22339
rect 29131 21860 29197 21861
rect 29131 21796 29132 21860
rect 29196 21796 29197 21860
rect 29131 21795 29197 21796
rect 29134 20773 29194 21795
rect 28763 20772 28829 20773
rect 28763 20708 28764 20772
rect 28828 20708 28829 20772
rect 28763 20707 28829 20708
rect 29131 20772 29197 20773
rect 29131 20708 29132 20772
rect 29196 20708 29197 20772
rect 29131 20707 29197 20708
rect 27659 17916 27725 17917
rect 27659 17852 27660 17916
rect 27724 17852 27725 17916
rect 27659 17851 27725 17852
rect 27107 14108 27173 14109
rect 27107 14044 27108 14108
rect 27172 14044 27173 14108
rect 27107 14043 27173 14044
rect 24347 12204 24413 12205
rect 24347 12140 24348 12204
rect 24412 12140 24413 12204
rect 24347 12139 24413 12140
rect 23243 11660 23309 11661
rect 23243 11596 23244 11660
rect 23308 11596 23309 11660
rect 23243 11595 23309 11596
rect 28766 10165 28826 20707
rect 29686 10165 29746 28323
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 30235 22540 30301 22541
rect 30235 22476 30236 22540
rect 30300 22476 30301 22540
rect 30235 22475 30301 22476
rect 30238 15197 30298 22475
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 30603 21316 30669 21317
rect 30603 21252 30604 21316
rect 30668 21252 30669 21316
rect 30603 21251 30669 21252
rect 30235 15196 30301 15197
rect 30235 15132 30236 15196
rect 30300 15132 30301 15196
rect 30235 15131 30301 15132
rect 28763 10164 28829 10165
rect 28763 10100 28764 10164
rect 28828 10100 28829 10164
rect 28763 10099 28829 10100
rect 29683 10164 29749 10165
rect 29683 10100 29684 10164
rect 29748 10100 29749 10164
rect 29683 10099 29749 10100
rect 30606 10029 30666 21251
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 30603 10028 30669 10029
rect 30603 9964 30604 10028
rect 30668 9964 30669 10028
rect 30603 9963 30669 9964
rect 23059 9620 23125 9621
rect 23059 9556 23060 9620
rect 23124 9556 23125 9620
rect 23059 9555 23125 9556
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 15147 6900 15213 6901
rect 15147 6836 15148 6900
rect 15212 6836 15213 6900
rect 15147 6835 15213 6836
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__inv_2  _0519_
timestamp -25199
transform -1 0 34500 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp -25199
transform 1 0 26312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0521_
timestamp -25199
transform -1 0 29348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0522_
timestamp -25199
transform 1 0 30912 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0523_
timestamp -25199
transform 1 0 34224 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0524_
timestamp -25199
transform -1 0 34224 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0525_
timestamp -25199
transform 1 0 32108 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0526_
timestamp -25199
transform -1 0 33396 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _0527_
timestamp -25199
transform 1 0 33212 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0528_
timestamp -25199
transform -1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0529_
timestamp -25199
transform -1 0 32936 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0530_
timestamp -25199
transform 1 0 28704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0531_
timestamp -25199
transform 1 0 29072 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0532_
timestamp -25199
transform -1 0 30912 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0533_
timestamp -25199
transform 1 0 31464 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0534_
timestamp -25199
transform -1 0 32476 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0535_
timestamp -25199
transform -1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0536_
timestamp -25199
transform -1 0 31464 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0537_
timestamp -25199
transform 1 0 31004 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0538_
timestamp -25199
transform -1 0 32660 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0539_
timestamp -25199
transform -1 0 30820 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0540_
timestamp -25199
transform 1 0 30820 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0541_
timestamp -25199
transform -1 0 29256 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0542_
timestamp -25199
transform 1 0 28336 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0543_
timestamp -25199
transform -1 0 30912 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0544_
timestamp -25199
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0545_
timestamp -25199
transform 1 0 28428 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0546_
timestamp -25199
transform 1 0 29808 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0547_
timestamp -25199
transform 1 0 30452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0548_
timestamp -25199
transform -1 0 30912 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0549_
timestamp -25199
transform 1 0 31188 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0550_
timestamp -25199
transform 1 0 31832 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0551_
timestamp -25199
transform -1 0 33304 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _0552_
timestamp -25199
transform 1 0 25668 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_1  _0553_
timestamp -25199
transform 1 0 26404 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _0554_
timestamp -25199
transform -1 0 26036 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0555_
timestamp -25199
transform 1 0 29900 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0556_
timestamp -25199
transform 1 0 27048 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0557_
timestamp -25199
transform -1 0 25944 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _0558_
timestamp -25199
transform -1 0 25576 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_2  _0559_
timestamp -25199
transform -1 0 30452 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _0560_
timestamp -25199
transform 1 0 28704 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0561_
timestamp -25199
transform -1 0 27876 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0562_
timestamp -25199
transform -1 0 26956 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _0563_
timestamp -25199
transform 1 0 26036 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0564_
timestamp -25199
transform 1 0 26956 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0565_
timestamp -25199
transform -1 0 25024 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0566_
timestamp -25199
transform 1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0567_
timestamp -25199
transform 1 0 27876 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0568_
timestamp -25199
transform -1 0 25668 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _0569_
timestamp -25199
transform 1 0 25944 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0570_
timestamp -25199
transform 1 0 6072 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0571_
timestamp -25199
transform 1 0 7636 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0572_
timestamp -25199
transform 1 0 8004 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0573_
timestamp -25199
transform 1 0 17204 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0574_
timestamp -25199
transform 1 0 17296 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0575_
timestamp -25199
transform 1 0 9844 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0576_
timestamp -25199
transform -1 0 10764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0577_
timestamp -25199
transform 1 0 10212 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0578_
timestamp -25199
transform 1 0 9936 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0579_
timestamp -25199
transform 1 0 17848 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0580_
timestamp -25199
transform 1 0 33856 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0581_
timestamp -25199
transform -1 0 21712 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0582_
timestamp -25199
transform 1 0 4140 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0583_
timestamp -25199
transform 1 0 13340 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0584_
timestamp -25199
transform 1 0 20424 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0585_
timestamp -25199
transform 1 0 4876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0586_
timestamp -25199
transform 1 0 12696 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0587_
timestamp -25199
transform 1 0 14260 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0588_
timestamp -25199
transform -1 0 15272 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0589_
timestamp -25199
transform 1 0 14812 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0590_
timestamp -25199
transform 1 0 21528 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0591_
timestamp -25199
transform 1 0 33856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0592_
timestamp -25199
transform 1 0 4324 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0593_
timestamp -25199
transform 1 0 16836 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0594_
timestamp -25199
transform 1 0 12420 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0595_
timestamp -25199
transform 1 0 18032 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0596_
timestamp -25199
transform 1 0 13800 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0597_
timestamp -25199
transform 1 0 7176 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0598_
timestamp -25199
transform 1 0 10764 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0599_
timestamp -25199
transform -1 0 9292 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0600_
timestamp -25199
transform 1 0 12236 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0601_
timestamp -25199
transform 1 0 18768 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0602_
timestamp -25199
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0603_
timestamp -25199
transform 1 0 21068 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0604_
timestamp -25199
transform 1 0 24656 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0605_
timestamp -25199
transform 1 0 23184 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0606_
timestamp -25199
transform 1 0 26404 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0607_
timestamp -25199
transform 1 0 27968 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0608_
timestamp -25199
transform -1 0 29348 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0609_
timestamp -25199
transform 1 0 25944 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0610_
timestamp -25199
transform 1 0 26312 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0611_
timestamp -25199
transform 1 0 26404 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0612_
timestamp -25199
transform -1 0 31464 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0613_
timestamp -25199
transform 1 0 31648 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0614_
timestamp -25199
transform 1 0 7176 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0615_
timestamp -25199
transform 1 0 5244 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0616_
timestamp -25199
transform 1 0 14536 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0617_
timestamp -25199
transform 1 0 15548 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0618_
timestamp -25199
transform 1 0 10856 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0619_
timestamp -25199
transform 1 0 7176 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0620_
timestamp -25199
transform 1 0 10764 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0621_
timestamp -25199
transform 1 0 8832 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0622_
timestamp -25199
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0623_
timestamp -25199
transform 1 0 15640 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0624_
timestamp -25199
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0625_
timestamp -25199
transform 1 0 21804 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0626_
timestamp -25199
transform 1 0 18584 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0627_
timestamp -25199
transform 1 0 20792 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0628_
timestamp -25199
transform -1 0 22448 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0629_
timestamp -25199
transform 1 0 27968 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0630_
timestamp -25199
transform 1 0 29072 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0631_
timestamp -25199
transform 1 0 25300 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0632_
timestamp -25199
transform 1 0 26956 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0633_
timestamp -25199
transform 1 0 29532 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0634_
timestamp -25199
transform -1 0 31924 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0635_
timestamp -25199
transform 1 0 32108 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0636_
timestamp -25199
transform 1 0 14536 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0637_
timestamp -25199
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0638_
timestamp -25199
transform 1 0 9660 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0639_
timestamp -25199
transform 1 0 8832 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0640_
timestamp -25199
transform 1 0 4600 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0641_
timestamp -25199
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0642_
timestamp -25199
transform -1 0 13524 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0643_
timestamp -25199
transform 1 0 10580 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0644_
timestamp -25199
transform 1 0 10028 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0645_
timestamp -25199
transform 1 0 16928 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0646_
timestamp -25199
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0647_
timestamp -25199
transform 1 0 28520 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0648_
timestamp -25199
transform 1 0 20516 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0649_
timestamp -25199
transform -1 0 29164 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0650_
timestamp -25199
transform 1 0 22356 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0651_
timestamp -25199
transform -1 0 24288 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0652_
timestamp -25199
transform 1 0 23460 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0653_
timestamp -25199
transform 1 0 19228 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0654_
timestamp -25199
transform -1 0 21988 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0655_
timestamp -25199
transform 1 0 24012 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0656_
timestamp -25199
transform 1 0 29624 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0657_
timestamp -25199
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0658_
timestamp -25199
transform 1 0 13524 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0659_
timestamp -25199
transform 1 0 15732 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0660_
timestamp -25199
transform 1 0 7176 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0661_
timestamp -25199
transform 1 0 8004 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0662_
timestamp -25199
transform 1 0 4784 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0663_
timestamp -25199
transform 1 0 4600 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0664_
timestamp -25199
transform 1 0 11040 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0665_
timestamp -25199
transform 1 0 9936 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0666_
timestamp -25199
transform 1 0 7912 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0667_
timestamp -25199
transform 1 0 16652 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0668_
timestamp -25199
transform 1 0 33948 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0669_
timestamp -25199
transform 1 0 29532 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0670_
timestamp -25199
transform 1 0 30360 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0671_
timestamp -25199
transform 1 0 25760 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0672_
timestamp -25199
transform -1 0 27600 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0673_
timestamp -25199
transform 1 0 23276 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0674_
timestamp -25199
transform 1 0 25392 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0675_
timestamp -25199
transform 1 0 22080 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0676_
timestamp -25199
transform 1 0 23920 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0677_
timestamp -25199
transform 1 0 26404 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0678_
timestamp -25199
transform 1 0 30636 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0679_
timestamp -25199
transform 1 0 33948 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0680_
timestamp -25199
transform 1 0 15456 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0681_
timestamp -25199
transform 1 0 7176 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0682_
timestamp -25199
transform 1 0 19228 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0683_
timestamp -25199
transform 1 0 19596 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0684_
timestamp -25199
transform 1 0 16744 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0685_
timestamp -25199
transform 1 0 16008 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0686_
timestamp -25199
transform 1 0 17112 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0687_
timestamp -25199
transform -1 0 9568 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0688_
timestamp -25199
transform 1 0 17480 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0689_
timestamp -25199
transform 1 0 19964 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0690_
timestamp -25199
transform 1 0 33764 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0691_
timestamp -25199
transform 1 0 26956 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0692_
timestamp -25199
transform -1 0 27692 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0693_
timestamp -25199
transform -1 0 12144 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0694_
timestamp -25199
transform -1 0 13156 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0695_
timestamp -25199
transform 1 0 4232 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0696_
timestamp -25199
transform 1 0 4784 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0697_
timestamp -25199
transform 1 0 8924 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0698_
timestamp -25199
transform 1 0 9936 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0699_
timestamp -25199
transform 1 0 11224 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0700_
timestamp -25199
transform 1 0 28612 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0701_
timestamp -25199
transform 1 0 33764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0702_
timestamp -25199
transform -1 0 30176 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0703_
timestamp -25199
transform 1 0 26956 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0704_
timestamp -25199
transform 1 0 23092 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0705_
timestamp -25199
transform 1 0 24380 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0706_
timestamp -25199
transform 1 0 25300 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0707_
timestamp -25199
transform 1 0 25852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0708_
timestamp -25199
transform 1 0 23184 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0709_
timestamp -25199
transform 1 0 26036 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0710_
timestamp -25199
transform 1 0 25852 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0711_
timestamp -25199
transform 1 0 30360 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0712_
timestamp -25199
transform 1 0 33580 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0713_
timestamp -25199
transform 1 0 14628 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0714_
timestamp -25199
transform 1 0 15456 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0715_
timestamp -25199
transform 1 0 10304 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0716_
timestamp -25199
transform -1 0 12236 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0717_
timestamp -25199
transform 1 0 9660 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0718_
timestamp -25199
transform 1 0 10488 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0719_
timestamp -25199
transform 1 0 4232 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0720_
timestamp -25199
transform 1 0 4784 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0721_
timestamp -25199
transform 1 0 10856 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0722_
timestamp -25199
transform 1 0 16652 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0723_
timestamp -25199
transform 1 0 33948 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0724_
timestamp -25199
transform 1 0 20424 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0725_
timestamp -25199
transform -1 0 28612 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0726_
timestamp -25199
transform 1 0 28244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0727_
timestamp -25199
transform 1 0 20516 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0728_
timestamp -25199
transform 1 0 18032 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0729_
timestamp -25199
transform 1 0 18676 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0730_
timestamp -25199
transform 1 0 20700 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0731_
timestamp -25199
transform 1 0 20976 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0732_
timestamp -25199
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0733_
timestamp -25199
transform 1 0 29256 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0734_
timestamp -25199
transform 1 0 32200 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0735_
timestamp -25199
transform 1 0 14352 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0736_
timestamp -25199
transform 1 0 14996 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0737_
timestamp -25199
transform -1 0 8188 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0738_
timestamp -25199
transform 1 0 7360 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0739_
timestamp -25199
transform 1 0 8188 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0740_
timestamp -25199
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0741_
timestamp -25199
transform -1 0 14260 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0742_
timestamp -25199
transform 1 0 12696 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0743_
timestamp -25199
transform 1 0 10028 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0744_
timestamp -25199
transform 1 0 17204 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0745_
timestamp -25199
transform 1 0 33948 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0746_
timestamp -25199
transform 1 0 32568 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0747_
timestamp -25199
transform -1 0 31464 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0748_
timestamp -25199
transform -1 0 31372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0749_
timestamp -25199
transform 1 0 31372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0750_
timestamp -25199
transform 1 0 29808 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0751_
timestamp -25199
transform 1 0 28704 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0752_
timestamp -25199
transform 1 0 28428 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0753_
timestamp -25199
transform -1 0 23092 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0754_
timestamp -25199
transform 1 0 21068 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0755_
timestamp -25199
transform 1 0 23092 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0756_
timestamp -25199
transform 1 0 24380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0757_
timestamp -25199
transform -1 0 24012 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0758_
timestamp -25199
transform 1 0 25116 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0759_
timestamp -25199
transform 1 0 23828 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0760_
timestamp -25199
transform 1 0 25208 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0761_
timestamp -25199
transform -1 0 24472 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0762_
timestamp -25199
transform 1 0 24840 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0763_
timestamp -25199
transform -1 0 23920 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0764_
timestamp -25199
transform 1 0 17848 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0765_
timestamp -25199
transform 1 0 20792 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0766_
timestamp -25199
transform 1 0 19228 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0767_
timestamp -25199
transform 1 0 30084 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp -25199
transform 1 0 16652 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0769_
timestamp -25199
transform 1 0 30544 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0770_
timestamp -25199
transform 1 0 16836 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0771_
timestamp -25199
transform 1 0 29900 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0772_
timestamp -25199
transform 1 0 16652 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0773_
timestamp -25199
transform 1 0 30636 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0774_
timestamp -25199
transform 1 0 19688 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0775_
timestamp -25199
transform 1 0 29532 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0776_
timestamp -25199
transform 1 0 30360 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0777_
timestamp -25199
transform 1 0 16652 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0778_
timestamp -25199
transform 1 0 29532 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0779_
timestamp -25199
transform -1 0 16560 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _0780_
timestamp -25199
transform -1 0 24840 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _0781_
timestamp -25199
transform 1 0 22632 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0782_
timestamp -25199
transform 1 0 17756 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0783_
timestamp -25199
transform 1 0 12328 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0784_
timestamp -25199
transform 1 0 11500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp -25199
transform 1 0 27048 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0786_
timestamp -25199
transform 1 0 11776 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0787_
timestamp -25199
transform 1 0 19872 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0788_
timestamp -25199
transform 1 0 12052 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp -25199
transform 1 0 23276 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0790_
timestamp -25199
transform 1 0 11500 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp -25199
transform 1 0 25484 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0792_
timestamp -25199
transform -1 0 17204 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp -25199
transform 1 0 12144 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0794_
timestamp -25199
transform 1 0 26956 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0795_
timestamp -25199
transform 1 0 11592 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0796_
timestamp -25199
transform 1 0 20792 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0797_
timestamp -25199
transform 1 0 12788 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _0798_
timestamp -25199
transform -1 0 23000 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_2  _0799_
timestamp -25199
transform -1 0 23276 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0800_
timestamp -25199
transform 1 0 16652 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0801_
timestamp -25199
transform 1 0 20332 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0802_
timestamp -25199
transform 1 0 2944 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0803_
timestamp -25199
transform 1 0 20332 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0804_
timestamp -25199
transform 1 0 4140 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp -25199
transform 1 0 23460 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0806_
timestamp -25199
transform 1 0 3772 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0807_
timestamp -25199
transform 1 0 18124 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp -25199
transform 1 0 3772 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0809_
timestamp -25199
transform 1 0 21436 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0810_
timestamp -25199
transform 1 0 17940 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0811_
timestamp -25199
transform 1 0 3864 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0812_
timestamp -25199
transform 1 0 21988 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0813_
timestamp -25199
transform 1 0 8924 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0814_
timestamp -25199
transform -1 0 19780 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0815_
timestamp -25199
transform 1 0 12788 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _0816_
timestamp -25199
transform 1 0 23184 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0817_
timestamp -25199
transform 1 0 16468 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0818_
timestamp -25199
transform 1 0 14168 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0819_
timestamp -25199
transform 1 0 14076 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0820_
timestamp -25199
transform 1 0 24932 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0821_
timestamp -25199
transform 1 0 12144 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0822_
timestamp -25199
transform 1 0 22264 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0823_
timestamp -25199
transform 1 0 14076 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0824_
timestamp -25199
transform 1 0 20792 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0825_
timestamp -25199
transform 1 0 12788 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0826_
timestamp -25199
transform 1 0 24840 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0827_
timestamp -25199
transform 1 0 16652 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0828_
timestamp -25199
transform 1 0 12512 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0829_
timestamp -25199
transform -1 0 26128 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0830_
timestamp -25199
transform 1 0 11684 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0831_
timestamp -25199
transform 1 0 19228 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0832_
timestamp -25199
transform 1 0 15548 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__nand4_2  _0833_
timestamp -25199
transform -1 0 25392 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0834_
timestamp -25199
transform 1 0 25116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0835_
timestamp -25199
transform 1 0 7360 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0836_
timestamp -25199
transform 1 0 15732 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0837_
timestamp -25199
transform 1 0 8924 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0838_
timestamp -25199
transform 1 0 23460 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0839_
timestamp -25199
transform 1 0 7912 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0840_
timestamp -25199
transform 1 0 26036 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0841_
timestamp -25199
transform 1 0 16652 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0842_
timestamp -25199
transform 1 0 27600 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0843_
timestamp -25199
transform 1 0 9016 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0844_
timestamp -25199
transform -1 0 21712 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0845_
timestamp -25199
transform 1 0 14628 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0846_
timestamp -25199
transform 1 0 10120 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0847_
timestamp -25199
transform 1 0 26956 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0848_
timestamp -25199
transform 1 0 15732 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0849_
timestamp -25199
transform 1 0 27692 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0850_
timestamp -25199
transform 1 0 7360 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0851_
timestamp -25199
transform -1 0 24656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0852_
timestamp -25199
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0853_
timestamp -25199
transform 1 0 20240 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0854_
timestamp -25199
transform 1 0 6348 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0855_
timestamp -25199
transform 1 0 29900 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0856_
timestamp -25199
transform -1 0 6900 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0857_
timestamp -25199
transform 1 0 28428 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0858_
timestamp -25199
transform 1 0 15456 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0859_
timestamp -25199
transform 1 0 19596 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0860_
timestamp -25199
transform 1 0 5796 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0861_
timestamp -25199
transform 1 0 29532 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0862_
timestamp -25199
transform 1 0 6348 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0863_
timestamp -25199
transform 1 0 8832 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0864_
timestamp -25199
transform 1 0 28520 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0865_
timestamp -25199
transform 1 0 8832 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0866_
timestamp -25199
transform 1 0 17756 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0867_
timestamp -25199
transform 1 0 13156 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0868_
timestamp -25199
transform -1 0 23828 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0869_
timestamp -25199
transform -1 0 11224 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0870_
timestamp -25199
transform 1 0 4876 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0871_
timestamp -25199
transform 1 0 9844 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0872_
timestamp -25199
transform 1 0 27232 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0873_
timestamp -25199
transform 1 0 15732 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0874_
timestamp -25199
transform 1 0 29992 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0875_
timestamp -25199
transform 1 0 10304 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0876_
timestamp -25199
transform 1 0 24932 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0877_
timestamp -25199
transform 1 0 5336 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0878_
timestamp -25199
transform 1 0 30268 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0879_
timestamp -25199
transform 1 0 18308 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0880_
timestamp -25199
transform 1 0 27600 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0881_
timestamp -25199
transform 1 0 22080 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0882_
timestamp -25199
transform 1 0 9568 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0883_
timestamp -25199
transform 1 0 20148 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0884_
timestamp -25199
transform 1 0 5428 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0885_
timestamp -25199
transform -1 0 23276 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0886_
timestamp -25199
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0887_
timestamp -25199
transform 1 0 20700 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0888_
timestamp -25199
transform 1 0 12788 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0889_
timestamp -25199
transform 1 0 22172 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0890_
timestamp -25199
transform 1 0 8004 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0891_
timestamp -25199
transform 1 0 18032 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0892_
timestamp -25199
transform 1 0 12420 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0893_
timestamp -25199
transform 1 0 27784 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0894_
timestamp -25199
transform 1 0 12696 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0895_
timestamp -25199
transform 1 0 26956 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0896_
timestamp -25199
transform 1 0 8004 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0897_
timestamp -25199
transform 1 0 7544 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0898_
timestamp -25199
transform 1 0 24564 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0899_
timestamp -25199
transform 1 0 8096 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0900_
timestamp -25199
transform 1 0 27508 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0901_
timestamp -25199
transform 1 0 9200 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_2  _0902_
timestamp -25199
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0903_
timestamp -25199
transform 1 0 24840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0904_
timestamp -25199
transform 1 0 8924 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0905_
timestamp -25199
transform 1 0 3772 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0906_
timestamp -25199
transform 1 0 18032 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0907_
timestamp -25199
transform 1 0 25484 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0908_
timestamp -25199
transform 1 0 9844 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0909_
timestamp -25199
transform 1 0 25208 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0910_
timestamp -25199
transform 1 0 5336 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0911_
timestamp -25199
transform 1 0 26956 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0912_
timestamp -25199
transform 1 0 14812 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0913_
timestamp -25199
transform 1 0 24564 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0914_
timestamp -25199
transform 1 0 15180 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0915_
timestamp -25199
transform 1 0 3588 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0916_
timestamp -25199
transform 1 0 23092 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0917_
timestamp -25199
transform 1 0 3956 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0918_
timestamp -25199
transform 1 0 21436 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0919_
timestamp -25199
transform 1 0 14444 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0920_
timestamp -25199
transform 1 0 24380 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0921_
timestamp -25199
transform 1 0 7268 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0922_
timestamp -25199
transform 1 0 14168 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0923_
timestamp -25199
transform 1 0 12328 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0924_
timestamp -25199
transform 1 0 27140 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0925_
timestamp -25199
transform 1 0 14536 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0926_
timestamp -25199
transform 1 0 21804 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0927_
timestamp -25199
transform 1 0 8924 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0928_
timestamp -25199
transform -1 0 20792 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0929_
timestamp -25199
transform 1 0 7912 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0930_
timestamp -25199
transform 1 0 24840 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0931_
timestamp -25199
transform 1 0 19688 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0932_
timestamp -25199
transform -1 0 27416 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0933_
timestamp -25199
transform 1 0 23276 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0934_
timestamp -25199
transform 1 0 14444 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0935_
timestamp -25199
transform 1 0 20240 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0936_
timestamp -25199
transform 1 0 7360 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0937_
timestamp -25199
transform 1 0 22908 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0938_
timestamp -25199
transform 1 0 5428 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0939_
timestamp -25199
transform 1 0 3312 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0940_
timestamp -25199
transform 1 0 3956 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0941_
timestamp -25199
transform 1 0 29900 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0942_
timestamp -25199
transform 1 0 4048 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0943_
timestamp -25199
transform 1 0 20056 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0944_
timestamp -25199
transform 1 0 3772 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0945_
timestamp -25199
transform 1 0 30544 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0946_
timestamp -25199
transform 1 0 3772 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0947_
timestamp -25199
transform 1 0 29532 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0948_
timestamp -25199
transform 1 0 6808 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0949_
timestamp -25199
transform 1 0 6348 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0950_
timestamp -25199
transform 1 0 29716 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0951_
timestamp -25199
transform 1 0 4968 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0952_
timestamp -25199
transform 1 0 28152 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0953_
timestamp -25199
transform 1 0 6716 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0954_
timestamp -25199
transform -1 0 23000 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0955_
timestamp -25199
transform 1 0 6992 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0956_
timestamp -25199
transform 1 0 14076 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0957_
timestamp -25199
transform 1 0 10948 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0958_
timestamp -25199
transform 1 0 21804 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0959_
timestamp -25199
transform 1 0 9936 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0960_
timestamp -25199
transform 1 0 17940 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0961_
timestamp -25199
transform 1 0 7084 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0962_
timestamp -25199
transform 1 0 22264 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0963_
timestamp -25199
transform 1 0 7176 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0964_
timestamp -25199
transform 1 0 21804 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0965_
timestamp -25199
transform -1 0 13984 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0966_
timestamp -25199
transform -1 0 12236 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0967_
timestamp -25199
transform 1 0 23276 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0968_
timestamp -25199
transform 1 0 11500 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0969_
timestamp -25199
transform 1 0 17940 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0970_
timestamp -25199
transform 1 0 14076 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__nand4_2  _0971_
timestamp -25199
transform -1 0 26312 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0972_
timestamp -25199
transform -1 0 25668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0973_
timestamp -25199
transform 1 0 10028 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0974_
timestamp -25199
transform 1 0 11500 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0975_
timestamp -25199
transform 1 0 16652 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0976_
timestamp -25199
transform -1 0 27508 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0977_
timestamp -25199
transform 1 0 14628 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0978_
timestamp -25199
transform 1 0 26956 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0979_
timestamp -25199
transform 1 0 10304 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0980_
timestamp -25199
transform 1 0 22356 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0981_
timestamp -25199
transform 1 0 14812 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0982_
timestamp -25199
transform 1 0 27140 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0983_
timestamp -25199
transform -1 0 19044 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0984_
timestamp -25199
transform 1 0 25576 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0985_
timestamp -25199
transform 1 0 24380 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0986_
timestamp -25199
transform 1 0 14536 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0987_
timestamp -25199
transform 1 0 19596 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0988_
timestamp -25199
transform 1 0 12788 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0989_
timestamp -25199
transform 1 0 24104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0990_
timestamp -25199
transform 1 0 4508 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0991_
timestamp -25199
transform 1 0 3772 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0992_
timestamp -25199
transform 1 0 17296 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0993_
timestamp -25199
transform 1 0 24380 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0994_
timestamp -25199
transform 1 0 2852 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0995_
timestamp -25199
transform 1 0 19964 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0996_
timestamp -25199
transform 1 0 8924 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0997_
timestamp -25199
transform 1 0 24748 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0998_
timestamp -25199
transform 1 0 10396 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0999_
timestamp -25199
transform 1 0 23092 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1000_
timestamp -25199
transform 1 0 16744 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1001_
timestamp -25199
transform 1 0 2576 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1002_
timestamp -25199
transform 1 0 24656 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1003_
timestamp -25199
transform 1 0 3036 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1004_
timestamp -25199
transform 1 0 17388 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1005_
timestamp -25199
transform 1 0 6348 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1006_
timestamp -25199
transform -1 0 23276 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1007_
timestamp -25199
transform 1 0 7636 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1008_
timestamp -25199
transform 1 0 20608 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1009_
timestamp -25199
transform 1 0 6348 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1010_
timestamp -25199
transform -1 0 29164 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1011_
timestamp -25199
transform -1 0 14720 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1012_
timestamp -25199
transform 1 0 28428 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1013_
timestamp -25199
transform 1 0 13616 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1014_
timestamp -25199
transform -1 0 23092 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1015_
timestamp -25199
transform 1 0 4140 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1016_
timestamp -25199
transform 1 0 22816 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1017_
timestamp -25199
transform 1 0 15088 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1018_
timestamp -25199
transform 1 0 4508 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1019_
timestamp -25199
transform 1 0 25116 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1020_
timestamp -25199
transform 1 0 4232 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1021_
timestamp -25199
transform 1 0 28428 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1022_
timestamp -25199
transform 1 0 9568 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1023_
timestamp -25199
transform -1 0 23552 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1024_
timestamp -25199
transform 1 0 9384 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1025_
timestamp -25199
transform 1 0 11684 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1026_
timestamp -25199
transform 1 0 15640 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1027_
timestamp -25199
transform 1 0 23828 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1028_
timestamp -25199
transform 1 0 6348 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1029_
timestamp -25199
transform 1 0 24288 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1030_
timestamp -25199
transform 1 0 7912 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1031_
timestamp -25199
transform 1 0 18216 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1032_
timestamp -25199
transform 1 0 6072 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1033_
timestamp -25199
transform 1 0 23000 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1034_
timestamp -25199
transform 1 0 19320 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1035_
timestamp -25199
transform 1 0 10120 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1036_
timestamp -25199
transform 1 0 22816 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1037_
timestamp -25199
transform 1 0 10120 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1038_
timestamp -25199
transform 1 0 19228 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1039_
timestamp -25199
transform 1 0 6256 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _1040_
timestamp -25199
transform 1 0 29532 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1041_
timestamp -25199
transform 1 0 32108 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1042_
timestamp -25199
transform 1 0 27048 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1043_
timestamp -25199
transform 1 0 29072 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1044_
timestamp -25199
transform 1 0 32660 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1045_
timestamp -25199
transform 1 0 33212 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1046_
timestamp -25199
transform 1 0 32752 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1047_
timestamp -25199
transform 1 0 33212 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1048_
timestamp -25199
transform 1 0 32108 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1049_
timestamp -25199
transform 1 0 33212 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1050_
timestamp -25199
transform 1 0 32384 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1051_
timestamp -25199
transform 1 0 32752 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1052_
timestamp -25199
transform 1 0 33212 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1053_
timestamp -25199
transform 1 0 32752 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1054_
timestamp -25199
transform 1 0 32752 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1055_
timestamp -25199
transform 1 0 33212 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1056_
timestamp -25199
transform 1 0 32752 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1057_
timestamp -25199
transform 1 0 32752 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1058_
timestamp -25199
transform 1 0 32752 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1059_
timestamp -25199
transform 1 0 32108 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1060_
timestamp -25199
transform 1 0 32752 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1061_
timestamp -25199
transform -1 0 34040 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1062_
timestamp -25199
transform 1 0 30728 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1063_
timestamp -25199
transform 1 0 30728 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1064_
timestamp -25199
transform 1 0 28336 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1065_
timestamp -25199
transform 1 0 22448 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1066_
timestamp -25199
transform 1 0 21160 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1067_
timestamp -25199
transform 1 0 24472 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1068_
timestamp -25199
transform -1 0 27876 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp -25199
transform 1 0 17388 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp -25199
transform 1 0 20332 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp -25199
transform 1 0 18308 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp -25199
transform 1 0 29808 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp -25199
transform -1 0 17112 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp -25199
transform 1 0 30360 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp -25199
transform 1 0 16652 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp -25199
transform 1 0 29624 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1077_
timestamp -25199
transform 1 0 16100 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp -25199
transform 1 0 30360 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp -25199
transform 1 0 19228 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp -25199
transform -1 0 29992 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp -25199
transform 1 0 29992 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp -25199
transform 1 0 15272 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp -25199
transform 1 0 29532 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp -25199
transform 1 0 16652 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp -25199
transform 1 0 17388 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp -25199
transform 1 0 11776 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp -25199
transform 1 0 10488 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp -25199
transform 1 0 26956 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp -25199
transform 1 0 11500 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp -25199
transform 1 0 19320 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp -25199
transform 1 0 11500 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp -25199
transform 1 0 22632 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp -25199
transform 1 0 9936 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp -25199
transform 1 0 24932 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp -25199
transform -1 0 18124 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp -25199
transform 1 0 11592 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1097_
timestamp -25199
transform 1 0 26036 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1098_
timestamp -25199
transform 1 0 10120 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp -25199
transform 1 0 20424 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp -25199
transform 1 0 12236 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp -25199
transform 1 0 15088 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp -25199
transform 1 0 18860 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp -25199
transform 1 0 2208 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1104_
timestamp -25199
transform 1 0 19780 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1105_
timestamp -25199
transform 1 0 3772 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1106_
timestamp -25199
transform 1 0 22264 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1107_
timestamp -25199
transform 1 0 2300 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1108_
timestamp -25199
transform 1 0 17572 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1109_
timestamp -25199
transform 1 0 2392 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1110_
timestamp -25199
transform 1 0 20884 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1111_
timestamp -25199
transform 1 0 17388 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1112_
timestamp -25199
transform 1 0 3404 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1113_
timestamp -25199
transform 1 0 21804 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1114_
timestamp -25199
transform 1 0 8372 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp -25199
transform 1 0 19228 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1116_
timestamp -25199
transform 1 0 11316 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1117_
timestamp -25199
transform 1 0 15916 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1118_
timestamp -25199
transform 1 0 14076 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1119_
timestamp -25199
transform 1 0 13708 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1120_
timestamp -25199
transform 1 0 24380 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1121_
timestamp -25199
transform -1 0 13156 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1122_
timestamp -25199
transform 1 0 20792 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1123_
timestamp -25199
transform 1 0 13524 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1124_
timestamp -25199
transform 1 0 19872 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1125_
timestamp -25199
transform 1 0 12144 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1126_
timestamp -25199
transform 1 0 24380 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1127_
timestamp -25199
transform 1 0 15916 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1128_
timestamp -25199
transform -1 0 13524 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1129_
timestamp -25199
transform -1 0 27324 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1130_
timestamp -25199
transform 1 0 11500 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1131_
timestamp -25199
transform 1 0 17664 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1132_
timestamp -25199
transform 1 0 15088 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1133_
timestamp -25199
transform 1 0 6808 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1134_
timestamp -25199
transform -1 0 15916 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1135_
timestamp -25199
transform 1 0 7360 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1136_
timestamp -25199
transform 1 0 22816 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1137_
timestamp -25199
transform 1 0 7360 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1138_
timestamp -25199
transform 1 0 25392 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1139_
timestamp -25199
transform 1 0 15732 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1140_
timestamp -25199
transform 1 0 27048 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1141_
timestamp -25199
transform 1 0 8464 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1142_
timestamp -25199
transform 1 0 21436 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1143_
timestamp -25199
transform 1 0 14076 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1144_
timestamp -25199
transform 1 0 9660 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1145_
timestamp -25199
transform -1 0 26864 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1146_
timestamp -25199
transform 1 0 15364 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1147_
timestamp -25199
transform 1 0 27324 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1148_
timestamp -25199
transform 1 0 6256 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1149_
timestamp -25199
transform 1 0 15732 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1150_
timestamp -25199
transform -1 0 20240 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1151_
timestamp -25199
transform 1 0 5336 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1152_
timestamp -25199
transform -1 0 29900 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1153_
timestamp -25199
transform 1 0 6348 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1154_
timestamp -25199
transform 1 0 27784 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1155_
timestamp -25199
transform 1 0 14904 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1156_
timestamp -25199
transform 1 0 19044 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1157_
timestamp -25199
transform 1 0 4784 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1158_
timestamp -25199
transform 1 0 27968 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1159_
timestamp -25199
transform 1 0 4692 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1160_
timestamp -25199
transform 1 0 8280 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1161_
timestamp -25199
transform 1 0 27968 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1162_
timestamp -25199
transform 1 0 8924 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1163_
timestamp -25199
transform 1 0 17204 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1164_
timestamp -25199
transform 1 0 11960 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1165_
timestamp -25199
transform -1 0 11408 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1166_
timestamp -25199
transform 1 0 4324 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1167_
timestamp -25199
transform 1 0 9292 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1168_
timestamp -25199
transform 1 0 26956 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1169_
timestamp -25199
transform 1 0 15088 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1170_
timestamp -25199
transform 1 0 29716 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1171_
timestamp -25199
transform 1 0 9752 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1172_
timestamp -25199
transform 1 0 24564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1173_
timestamp -25199
transform 1 0 3864 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1174_
timestamp -25199
transform 1 0 30084 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1175_
timestamp -25199
transform 1 0 17664 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1176_
timestamp -25199
transform 1 0 27140 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1177_
timestamp -25199
transform 1 0 21804 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1178_
timestamp -25199
transform 1 0 9476 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1179_
timestamp -25199
transform 1 0 19596 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1180_
timestamp -25199
transform 1 0 4784 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1181_
timestamp -25199
transform 1 0 7912 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1182_
timestamp -25199
transform 1 0 19228 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1183_
timestamp -25199
transform 1 0 12328 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1184_
timestamp -25199
transform 1 0 21804 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1185_
timestamp -25199
transform 1 0 7360 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1186_
timestamp -25199
transform 1 0 17480 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1187_
timestamp -25199
transform 1 0 11592 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1188_
timestamp -25199
transform 1 0 27508 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1189_
timestamp -25199
transform 1 0 12144 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1190_
timestamp -25199
transform 1 0 26312 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1191_
timestamp -25199
transform 1 0 7912 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1192_
timestamp -25199
transform 1 0 6808 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1193_
timestamp -25199
transform 1 0 24380 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1194_
timestamp -25199
transform 1 0 7360 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1195_
timestamp -25199
transform 1 0 27324 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1196_
timestamp -25199
transform 1 0 7728 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1197_
timestamp -25199
transform 1 0 8372 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1198_
timestamp -25199
transform 1 0 2852 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1199_
timestamp -25199
transform 1 0 17572 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1200_
timestamp -25199
transform 1 0 24932 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1201_
timestamp -25199
transform 1 0 9292 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1202_
timestamp -25199
transform 1 0 24656 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1203_
timestamp -25199
transform 1 0 4784 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1204_
timestamp -25199
transform 1 0 26036 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1205_
timestamp -25199
transform 1 0 14260 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1206_
timestamp -25199
transform 1 0 24012 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1207_
timestamp -25199
transform 1 0 13708 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1208_
timestamp -25199
transform 1 0 2852 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1209_
timestamp -25199
transform 1 0 22540 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1210_
timestamp -25199
transform 1 0 3404 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1211_
timestamp -25199
transform 1 0 21068 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1212_
timestamp -25199
transform 1 0 14076 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1213_
timestamp -25199
transform 1 0 6440 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1214_
timestamp -25199
transform 1 0 13616 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1215_
timestamp -25199
transform 1 0 11776 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1216_
timestamp -25199
transform 1 0 25668 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1217_
timestamp -25199
transform 1 0 13064 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1218_
timestamp -25199
transform 1 0 21252 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1219_
timestamp -25199
transform 1 0 7728 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1220_
timestamp -25199
transform -1 0 20700 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1221_
timestamp -25199
transform -1 0 7912 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1222_
timestamp -25199
transform 1 0 24288 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1223_
timestamp -25199
transform 1 0 19320 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1224_
timestamp -25199
transform -1 0 28428 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1225_
timestamp -25199
transform 1 0 22724 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1226_
timestamp -25199
transform 1 0 12972 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1227_
timestamp -25199
transform 1 0 19688 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1228_
timestamp -25199
transform 1 0 6716 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1229_
timestamp -25199
transform 1 0 5244 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1230_
timestamp -25199
transform -1 0 3312 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1231_
timestamp -25199
transform 1 0 3772 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1232_
timestamp -25199
transform -1 0 29900 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1233_
timestamp -25199
transform 1 0 3496 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1234_
timestamp -25199
transform 1 0 19504 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1235_
timestamp -25199
transform 1 0 3772 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1236_
timestamp -25199
transform -1 0 30912 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1237_
timestamp -25199
transform -1 0 3312 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1238_
timestamp -25199
transform 1 0 28612 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1239_
timestamp -25199
transform 1 0 6164 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1240_
timestamp -25199
transform 1 0 5336 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1241_
timestamp -25199
transform 1 0 29440 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1242_
timestamp -25199
transform -1 0 4048 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1243_
timestamp -25199
transform 1 0 26680 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1244_
timestamp -25199
transform 1 0 5244 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1245_
timestamp -25199
transform 1 0 6072 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1246_
timestamp -25199
transform 1 0 12512 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1247_
timestamp -25199
transform 1 0 9936 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1248_
timestamp -25199
transform 1 0 20424 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1249_
timestamp -25199
transform 1 0 9384 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1250_
timestamp -25199
transform 1 0 17480 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1251_
timestamp -25199
transform 1 0 5612 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1252_
timestamp -25199
transform 1 0 20792 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1253_
timestamp -25199
transform 1 0 6624 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1254_
timestamp -25199
transform 1 0 20884 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1255_
timestamp -25199
transform 1 0 13340 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1256_
timestamp -25199
transform -1 0 12972 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1257_
timestamp -25199
transform 1 0 22172 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1258_
timestamp -25199
transform 1 0 11040 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1259_
timestamp -25199
transform 1 0 17388 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1260_
timestamp -25199
transform 1 0 13432 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1261_
timestamp -25199
transform 1 0 9384 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1262_
timestamp -25199
transform 1 0 11500 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1263_
timestamp -25199
transform 1 0 15916 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1264_
timestamp -25199
transform -1 0 28428 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1265_
timestamp -25199
transform 1 0 14076 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1266_
timestamp -25199
transform 1 0 26956 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1267_
timestamp -25199
transform 1 0 9752 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1268_
timestamp -25199
transform 1 0 21804 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1269_
timestamp -25199
transform 1 0 14260 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1270_
timestamp -25199
transform 1 0 26956 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1271_
timestamp -25199
transform -1 0 19136 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1272_
timestamp -25199
transform 1 0 25024 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1273_
timestamp -25199
transform 1 0 24380 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1274_
timestamp -25199
transform 1 0 14076 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1275_
timestamp -25199
transform 1 0 19228 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1276_
timestamp -25199
transform 1 0 12328 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1277_
timestamp -25199
transform 1 0 3772 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1278_
timestamp -25199
transform -1 0 3956 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1279_
timestamp -25199
transform 1 0 16744 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1280_
timestamp -25199
transform 1 0 22816 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1281_
timestamp -25199
transform 1 0 2208 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1282_
timestamp -25199
transform 1 0 19412 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1283_
timestamp -25199
transform 1 0 8096 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1284_
timestamp -25199
transform 1 0 23276 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1285_
timestamp -25199
transform 1 0 9844 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1286_
timestamp -25199
transform 1 0 22540 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1287_
timestamp -25199
transform 1 0 16652 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1288_
timestamp -25199
transform 1 0 2208 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1289_
timestamp -25199
transform 1 0 24380 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1290_
timestamp -25199
transform 1 0 2208 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1291_
timestamp -25199
transform 1 0 16928 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1292_
timestamp -25199
transform 1 0 5244 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1293_
timestamp -25199
transform 1 0 6992 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1294_
timestamp -25199
transform 1 0 20332 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1295_
timestamp -25199
transform 1 0 5520 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1296_
timestamp -25199
transform -1 0 29440 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1297_
timestamp -25199
transform 1 0 14076 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1298_
timestamp -25199
transform 1 0 28152 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1299_
timestamp -25199
transform 1 0 13064 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1300_
timestamp -25199
transform -1 0 23276 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1301_
timestamp -25199
transform 1 0 3312 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1302_
timestamp -25199
transform 1 0 22264 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1303_
timestamp -25199
transform 1 0 14536 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1304_
timestamp -25199
transform 1 0 3864 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1305_
timestamp -25199
transform 1 0 24564 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1306_
timestamp -25199
transform 1 0 3772 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1307_
timestamp -25199
transform 1 0 28060 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1308_
timestamp -25199
transform 1 0 8096 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1309_
timestamp -25199
transform 1 0 8464 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1310_
timestamp -25199
transform 1 0 11592 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1311_
timestamp -25199
transform 1 0 15088 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1312_
timestamp -25199
transform 1 0 22356 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1313_
timestamp -25199
transform 1 0 5336 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1314_
timestamp -25199
transform 1 0 23276 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1315_
timestamp -25199
transform 1 0 7360 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1316_
timestamp -25199
transform 1 0 17664 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1317_
timestamp -25199
transform 1 0 5428 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1318_
timestamp -25199
transform 1 0 22540 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1319_
timestamp -25199
transform 1 0 18952 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1320_
timestamp -25199
transform 1 0 9568 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1321_
timestamp -25199
transform 1 0 22264 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1322_
timestamp -25199
transform 1 0 9568 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1323_
timestamp -25199
transform 1 0 18584 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1324_
timestamp -25199
transform -1 0 7820 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -25199
transform 1 0 8372 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0525__B1
timestamp -25199
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0526__B1
timestamp -25199
transform -1 0 33764 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__B1
timestamp -25199
transform 1 0 33028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0528__B1
timestamp -25199
transform -1 0 33856 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__A2
timestamp -25199
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__X
timestamp -25199
transform -1 0 30636 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__B1
timestamp -25199
transform 1 0 6716 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__A2
timestamp -25199
transform 1 0 8556 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__B1
timestamp -25199
transform 1 0 8372 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0572__A2
timestamp -25199
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0572__B1
timestamp -25199
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__A2
timestamp -25199
transform 1 0 18860 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__B1
timestamp -25199
transform 1 0 17848 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__A2
timestamp -25199
transform 1 0 18216 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__B1
timestamp -25199
transform 1 0 18032 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__A2
timestamp -25199
transform -1 0 10856 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__B1
timestamp -25199
transform -1 0 10672 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__A2
timestamp -25199
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__B1
timestamp -25199
transform 1 0 9844 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__A2
timestamp -25199
transform -1 0 11040 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__C1
timestamp -25199
transform -1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__A2
timestamp -25199
transform -1 0 19044 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__C1
timestamp -25199
transform 1 0 18676 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__A2
timestamp -25199
transform -1 0 22540 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__B1
timestamp -25199
transform 1 0 4784 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__A2
timestamp -25199
transform 1 0 14168 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__B1
timestamp -25199
transform 1 0 13984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__A2
timestamp -25199
transform -1 0 21988 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__B1
timestamp -25199
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__A2
timestamp -25199
transform 1 0 5796 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__B1
timestamp -25199
transform 1 0 5612 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__A2
timestamp -25199
transform 1 0 13524 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__B1
timestamp -25199
transform 1 0 13340 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__A2
timestamp -25199
transform 1 0 14996 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__B1
timestamp -25199
transform 1 0 15180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__A2
timestamp -25199
transform 1 0 16008 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__C1
timestamp -25199
transform 1 0 15824 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A2
timestamp -25199
transform 1 0 23000 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__C1
timestamp -25199
transform 1 0 22356 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__B1
timestamp -25199
transform 1 0 4968 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__A2
timestamp -25199
transform 1 0 17480 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__B1
timestamp -25199
transform 1 0 17664 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__A2
timestamp -25199
transform 1 0 13248 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__B1
timestamp -25199
transform 1 0 13064 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__A2
timestamp -25199
transform 1 0 18768 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__B1
timestamp -25199
transform -1 0 19964 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__A2
timestamp -25199
transform 1 0 14720 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__B1
timestamp -25199
transform 1 0 14536 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__A2
timestamp -25199
transform 1 0 8004 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__B1
timestamp -25199
transform 1 0 7820 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0598__A2
timestamp -25199
transform 1 0 12604 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0598__B1
timestamp -25199
transform 1 0 12788 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__A2
timestamp -25199
transform 1 0 9292 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__C1
timestamp -25199
transform 1 0 9476 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__A2
timestamp -25199
transform 1 0 19964 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__C1
timestamp -25199
transform 1 0 19596 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__A2
timestamp -25199
transform -1 0 23000 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__B1
timestamp -25199
transform 1 0 20884 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__A2
timestamp -25199
transform 1 0 26404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__B1
timestamp -25199
transform 1 0 25668 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__A2
timestamp -25199
transform 1 0 24840 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__B1
timestamp -25199
transform 1 0 23920 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__A2
timestamp -25199
transform 1 0 27140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__B1
timestamp -25199
transform -1 0 26772 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__A2
timestamp -25199
transform -1 0 29348 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__B1
timestamp -25199
transform -1 0 28612 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__A2
timestamp -25199
transform -1 0 30268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__A2
timestamp -25199
transform -1 0 27508 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__B1
timestamp -25199
transform 1 0 27508 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__A2
timestamp -25199
transform 1 0 26128 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__D1
timestamp -25199
transform 1 0 27692 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__A2
timestamp -25199
transform 1 0 31464 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__B
timestamp -25199
transform 1 0 7636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__A2
timestamp -25199
transform 1 0 5888 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__B1
timestamp -25199
transform 1 0 5888 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__A2
timestamp -25199
transform 1 0 15364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__B1
timestamp -25199
transform 1 0 14352 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__A2
timestamp -25199
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__B1
timestamp -25199
transform 1 0 16284 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__A2
timestamp -25199
transform 1 0 11592 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__B1
timestamp -25199
transform 1 0 13156 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__B1
timestamp -25199
transform 1 0 8372 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__A2
timestamp -25199
transform 1 0 12512 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__B1
timestamp -25199
transform 1 0 11500 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__A2
timestamp -25199
transform 1 0 9752 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__B1
timestamp -25199
transform 1 0 9568 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__A
timestamp -25199
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__A2
timestamp -25199
transform 1 0 17480 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__C1
timestamp -25199
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__X
timestamp -25199
transform -1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0624__B1
timestamp -25199
transform 1 0 33764 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__A2
timestamp -25199
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__B1
timestamp -25199
transform 1 0 22816 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__A2
timestamp -25199
transform 1 0 19320 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__C1
timestamp -25199
transform 1 0 19504 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__A2
timestamp -25199
transform -1 0 21712 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__B1
timestamp -25199
transform 1 0 21712 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__A2
timestamp -25199
transform 1 0 23000 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__A2
timestamp -25199
transform 1 0 29716 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__B1
timestamp -25199
transform -1 0 29716 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__A2
timestamp -25199
transform 1 0 30084 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__A2
timestamp -25199
transform -1 0 27692 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__A2
timestamp -25199
transform 1 0 27784 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__B1
timestamp -25199
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__A2
timestamp -25199
transform 1 0 32108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__B1
timestamp -25199
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__A2
timestamp -25199
transform -1 0 15364 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__B1
timestamp -25199
transform 1 0 15272 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__A2
timestamp -25199
transform 1 0 17572 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__B1
timestamp -25199
transform 1 0 17388 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__A2
timestamp -25199
transform 1 0 10304 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__B1
timestamp -25199
transform 1 0 10488 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__A2
timestamp -25199
transform 1 0 9660 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__B1
timestamp -25199
transform 1 0 9476 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__B1
timestamp -25199
transform 1 0 5244 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__A2
timestamp -25199
transform 1 0 7176 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__B1
timestamp -25199
transform 1 0 7084 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__A2
timestamp -25199
transform 1 0 13708 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__B1
timestamp -25199
transform 1 0 13524 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__A2
timestamp -25199
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__C1
timestamp -25199
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__A2
timestamp -25199
transform 1 0 17940 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__C1
timestamp -25199
transform -1 0 17940 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__A2
timestamp -25199
transform 1 0 29256 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__A2
timestamp -25199
transform 1 0 20424 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__B1
timestamp -25199
transform -1 0 21344 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A2
timestamp -25199
transform 1 0 27416 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__A2
timestamp -25199
transform 1 0 23092 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__B1
timestamp -25199
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__A2
timestamp -25199
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__B1
timestamp -25199
transform 1 0 24564 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__A2
timestamp -25199
transform 1 0 24288 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__B1
timestamp -25199
transform 1 0 24104 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__A2
timestamp -25199
transform 1 0 20792 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__B1
timestamp -25199
transform 1 0 20424 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__A2
timestamp -25199
transform 1 0 21988 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__B1
timestamp -25199
transform 1 0 22172 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__A2
timestamp -25199
transform 1 0 30820 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__C1
timestamp -25199
transform -1 0 29440 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A2
timestamp -25199
transform -1 0 14536 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__B1
timestamp -25199
transform -1 0 14352 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__A2
timestamp -25199
transform -1 0 17112 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__B1
timestamp -25199
transform 1 0 17112 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__A2
timestamp -25199
transform 1 0 8004 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__B1
timestamp -25199
transform 1 0 7820 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__A2
timestamp -25199
transform -1 0 9016 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__B1
timestamp -25199
transform -1 0 8832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__A2
timestamp -25199
transform 1 0 5612 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__B1
timestamp -25199
transform 1 0 5428 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__A2
timestamp -25199
transform 1 0 5244 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__A2
timestamp -25199
transform 1 0 11868 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__B1
timestamp -25199
transform 1 0 11684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__A2
timestamp -25199
transform 1 0 10580 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__C1
timestamp -25199
transform 1 0 10764 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__A2
timestamp -25199
transform -1 0 17848 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__C1
timestamp -25199
transform 1 0 17480 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__B
timestamp -25199
transform 1 0 29992 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__A2
timestamp -25199
transform 1 0 29992 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__B1
timestamp -25199
transform -1 0 31280 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A2
timestamp -25199
transform 1 0 26680 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__B1
timestamp -25199
transform 1 0 25760 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__C1
timestamp -25199
transform -1 0 27968 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A2
timestamp -25199
transform 1 0 27968 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__B1
timestamp -25199
transform 1 0 28980 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A2
timestamp -25199
transform -1 0 24288 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__B1
timestamp -25199
transform -1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A2
timestamp -25199
transform 1 0 25484 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__B1
timestamp -25199
transform 1 0 26312 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A2
timestamp -25199
transform 1 0 23276 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__B1
timestamp -25199
transform 1 0 23092 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A2
timestamp -25199
transform 1 0 25392 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__B1
timestamp -25199
transform 1 0 25208 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A2
timestamp -25199
transform 1 0 31464 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__C1
timestamp -25199
transform 1 0 30452 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__A2
timestamp -25199
transform 1 0 16192 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__B1
timestamp -25199
transform -1 0 16284 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__B1
timestamp -25199
transform 1 0 7820 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__A2
timestamp -25199
transform 1 0 20148 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__B1
timestamp -25199
transform 1 0 20332 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A2
timestamp -25199
transform 1 0 18124 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__B1
timestamp -25199
transform 1 0 17940 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A2
timestamp -25199
transform 1 0 16008 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__B1
timestamp -25199
transform 1 0 15824 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__A2
timestamp -25199
transform 1 0 16928 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__B1
timestamp -25199
transform 1 0 18032 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__A2
timestamp -25199
transform 1 0 9568 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__C1
timestamp -25199
transform 1 0 9752 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__A2
timestamp -25199
transform 1 0 20976 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__C1
timestamp -25199
transform 1 0 20792 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A2
timestamp -25199
transform 1 0 28612 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__B1
timestamp -25199
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A2
timestamp -25199
transform 1 0 12328 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__B1
timestamp -25199
transform 1 0 12512 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A2
timestamp -25199
transform 1 0 12236 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__B1
timestamp -25199
transform 1 0 13156 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__C1
timestamp -25199
transform 1 0 13524 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__A2
timestamp -25199
transform 1 0 4876 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__B1
timestamp -25199
transform 1 0 5060 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__B1
timestamp -25199
transform 1 0 5980 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__B1
timestamp -25199
transform 1 0 9660 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A2
timestamp -25199
transform 1 0 10856 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__B1
timestamp -25199
transform 1 0 10672 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A2
timestamp -25199
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A2
timestamp -25199
transform -1 0 30544 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__B1
timestamp -25199
transform -1 0 30728 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__A2
timestamp -25199
transform 1 0 28244 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__B1
timestamp -25199
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A2
timestamp -25199
transform -1 0 26128 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__B1
timestamp -25199
transform 1 0 26128 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A2
timestamp -25199
transform -1 0 26680 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__B1
timestamp -25199
transform -1 0 26496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__B1
timestamp -25199
transform 1 0 27140 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A2
timestamp -25199
transform -1 0 24012 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__B1
timestamp -25199
transform -1 0 24196 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A2
timestamp -25199
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__C1
timestamp -25199
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A2
timestamp -25199
transform 1 0 31556 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__B
timestamp -25199
transform -1 0 15272 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A2
timestamp -25199
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__B1
timestamp -25199
transform 1 0 16192 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A2
timestamp -25199
transform 1 0 11132 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__B1
timestamp -25199
transform 1 0 10948 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A2
timestamp -25199
transform 1 0 12236 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__B1
timestamp -25199
transform 1 0 12604 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__C1
timestamp -25199
transform 1 0 12420 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A2
timestamp -25199
transform 1 0 10488 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__B1
timestamp -25199
transform 1 0 10304 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A2
timestamp -25199
transform -1 0 11592 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__B1
timestamp -25199
transform -1 0 11408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__B1
timestamp -25199
transform 1 0 4876 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__B1
timestamp -25199
transform -1 0 5704 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__A2
timestamp -25199
transform 1 0 17572 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__C1
timestamp -25199
transform 1 0 17480 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A2
timestamp -25199
transform -1 0 21436 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__B1
timestamp -25199
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A2
timestamp -25199
transform -1 0 28980 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__B1
timestamp -25199
transform 1 0 28612 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__B1
timestamp -25199
transform 1 0 28980 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A2
timestamp -25199
transform 1 0 21344 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__B1
timestamp -25199
transform 1 0 21160 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A2
timestamp -25199
transform 1 0 18676 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__B1
timestamp -25199
transform 1 0 18768 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A2
timestamp -25199
transform 1 0 19412 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__B1
timestamp -25199
transform 1 0 18492 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A2
timestamp -25199
transform -1 0 21528 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A2
timestamp -25199
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__C1
timestamp -25199
transform 1 0 21988 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A2
timestamp -25199
transform 1 0 30084 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A2
timestamp -25199
transform -1 0 15364 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__B1
timestamp -25199
transform -1 0 15180 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A2
timestamp -25199
transform -1 0 16100 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B1
timestamp -25199
transform -1 0 15916 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__B1
timestamp -25199
transform -1 0 8372 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A2
timestamp -25199
transform -1 0 8464 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__B1
timestamp -25199
transform -1 0 8280 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A2
timestamp -25199
transform -1 0 9200 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__B1
timestamp -25199
transform -1 0 9384 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B1
timestamp -25199
transform 1 0 9660 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A2
timestamp -25199
transform 1 0 14352 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__B1
timestamp -25199
transform 1 0 14260 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__A2
timestamp -25199
transform 1 0 13340 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__C1
timestamp -25199
transform -1 0 13708 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__A2
timestamp -25199
transform 1 0 18216 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__C1
timestamp -25199
transform -1 0 18216 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A1
timestamp -25199
transform 1 0 28980 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__S
timestamp -25199
transform -1 0 18860 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__S
timestamp -25199
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__S
timestamp -25199
transform 1 0 20056 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__S
timestamp -25199
transform -1 0 30636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__S
timestamp -25199
transform 1 0 17480 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__S
timestamp -25199
transform 1 0 30360 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__S
timestamp -25199
transform 1 0 17664 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__S
timestamp -25199
transform 1 0 30912 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__S
timestamp -25199
transform 1 0 17480 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__S
timestamp -25199
transform 1 0 31464 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__S
timestamp -25199
transform 1 0 20516 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A0
timestamp -25199
transform 1 0 29348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__S
timestamp -25199
transform 1 0 17480 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__S
timestamp -25199
transform -1 0 16744 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__S
timestamp -25199
transform 1 0 18584 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__S
timestamp -25199
transform -1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__S
timestamp -25199
transform 1 0 12420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__S
timestamp -25199
transform -1 0 28060 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__S
timestamp -25199
transform 1 0 12604 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__S
timestamp -25199
transform 1 0 20700 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__S
timestamp -25199
transform -1 0 13064 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__S
timestamp -25199
transform -1 0 24288 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__S
timestamp -25199
transform 1 0 12328 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__S
timestamp -25199
transform -1 0 26680 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__S
timestamp -25199
transform 1 0 17204 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__S
timestamp -25199
transform 1 0 12972 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__S
timestamp -25199
transform 1 0 27784 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__S
timestamp -25199
transform 1 0 12420 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__S
timestamp -25199
transform -1 0 21988 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__S
timestamp -25199
transform 1 0 13708 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__Y
timestamp -25199
transform -1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__S
timestamp -25199
transform 1 0 17480 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__S
timestamp -25199
transform -1 0 20332 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__S
timestamp -25199
transform 1 0 3772 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__S
timestamp -25199
transform 1 0 20148 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__S
timestamp -25199
transform 1 0 4968 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__S
timestamp -25199
transform 1 0 23736 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__S
timestamp -25199
transform 1 0 4600 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__S
timestamp -25199
transform -1 0 19136 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__S
timestamp -25199
transform 1 0 4600 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__S
timestamp -25199
transform 1 0 4876 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__S
timestamp -25199
transform -1 0 9936 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__S
timestamp -25199
transform 1 0 13616 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__S
timestamp -25199
transform 1 0 17664 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__S
timestamp -25199
transform 1 0 14996 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__S
timestamp -25199
transform 1 0 14904 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__S
timestamp -25199
transform 1 0 25760 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__S
timestamp -25199
transform 1 0 12972 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__S
timestamp -25199
transform 1 0 22448 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__S
timestamp -25199
transform 1 0 14904 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__S
timestamp -25199
transform 1 0 21620 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__S
timestamp -25199
transform 1 0 13616 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__S
timestamp -25199
transform 1 0 25668 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__S
timestamp -25199
transform 1 0 17756 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__S
timestamp -25199
transform 1 0 13340 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__S
timestamp -25199
transform -1 0 26312 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__S
timestamp -25199
transform 1 0 12512 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__S
timestamp -25199
transform -1 0 20240 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__S
timestamp -25199
transform -1 0 16560 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__S
timestamp -25199
transform -1 0 8372 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__S
timestamp -25199
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__S
timestamp -25199
transform 1 0 9752 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__S
timestamp -25199
transform 1 0 24656 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__S
timestamp -25199
transform 1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__S
timestamp -25199
transform 1 0 26588 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__S
timestamp -25199
transform -1 0 17664 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__S
timestamp -25199
transform -1 0 10028 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__S
timestamp -25199
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__S
timestamp -25199
transform 1 0 15916 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__S
timestamp -25199
transform 1 0 10948 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__S
timestamp -25199
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__S
timestamp -25199
transform -1 0 8372 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__S
timestamp -25199
transform 1 0 18216 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__S
timestamp -25199
transform 1 0 7176 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__S
timestamp -25199
transform 1 0 6900 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__S
timestamp -25199
transform 1 0 16284 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__S
timestamp -25199
transform 1 0 19412 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__S
timestamp -25199
transform 1 0 6624 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__S
timestamp -25199
transform -1 0 31464 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__S
timestamp -25199
transform 1 0 8004 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__S
timestamp -25199
transform 1 0 9660 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__S
timestamp -25199
transform -1 0 30360 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__S
timestamp -25199
transform 1 0 9660 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__S
timestamp -25199
transform 1 0 18584 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__S
timestamp -25199
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__S
timestamp -25199
transform -1 0 11408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A1
timestamp -25199
transform -1 0 4876 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__S
timestamp -25199
transform 1 0 5704 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__S
timestamp -25199
transform 1 0 10764 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__S
timestamp -25199
transform -1 0 28244 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__S
timestamp -25199
transform -1 0 17480 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__S
timestamp -25199
transform -1 0 31188 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__S
timestamp -25199
transform 1 0 11132 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__S
timestamp -25199
transform 1 0 25760 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__S
timestamp -25199
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__S
timestamp -25199
transform 1 0 29808 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__S
timestamp -25199
transform 1 0 19136 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A1
timestamp -25199
transform 1 0 26496 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__S
timestamp -25199
transform 1 0 28428 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__S
timestamp -25199
transform 1 0 22908 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__S
timestamp -25199
transform -1 0 11684 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__S
timestamp -25199
transform -1 0 21160 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__S
timestamp -25199
transform 1 0 6900 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__S
timestamp -25199
transform -1 0 9936 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__S
timestamp -25199
transform 1 0 21160 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__S
timestamp -25199
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__S
timestamp -25199
transform 1 0 21988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__S
timestamp -25199
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__S
timestamp -25199
transform 1 0 18860 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__S
timestamp -25199
transform -1 0 13432 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__S
timestamp -25199
transform 1 0 27600 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__S
timestamp -25199
transform -1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__S
timestamp -25199
transform -1 0 28704 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__S
timestamp -25199
transform 1 0 8832 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__S
timestamp -25199
transform 1 0 8464 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__S
timestamp -25199
transform -1 0 24564 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__S
timestamp -25199
transform -1 0 9108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__S
timestamp -25199
transform -1 0 27508 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__S
timestamp -25199
transform 1 0 10488 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__S
timestamp -25199
transform -1 0 9936 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__A1
timestamp -25199
transform -1 0 3680 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__S
timestamp -25199
transform 1 0 5888 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__S
timestamp -25199
transform 1 0 18860 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__S
timestamp -25199
transform 1 0 26864 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__S
timestamp -25199
transform 1 0 10764 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__S
timestamp -25199
transform 1 0 26036 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__S
timestamp -25199
transform 1 0 6256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A1
timestamp -25199
transform -1 0 26588 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__S
timestamp -25199
transform -1 0 26772 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__S
timestamp -25199
transform 1 0 15640 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__S
timestamp -25199
transform 1 0 26128 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__S
timestamp -25199
transform 1 0 16008 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__S
timestamp -25199
transform 1 0 4416 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__S
timestamp -25199
transform 1 0 22908 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__S
timestamp -25199
transform 1 0 5060 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__S
timestamp -25199
transform 1 0 22264 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__S
timestamp -25199
transform -1 0 15456 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__Y
timestamp -25199
transform -1 0 25852 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__S
timestamp -25199
transform 1 0 8096 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__S
timestamp -25199
transform 1 0 14996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__S
timestamp -25199
transform 1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__S
timestamp -25199
transform -1 0 28796 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__S
timestamp -25199
transform 1 0 15272 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__S
timestamp -25199
transform 1 0 22632 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__S
timestamp -25199
transform -1 0 9936 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__S
timestamp -25199
transform 1 0 21252 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__S
timestamp -25199
transform 1 0 8740 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__S
timestamp -25199
transform 1 0 24656 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A1
timestamp -25199
transform -1 0 26588 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__S
timestamp -25199
transform -1 0 15456 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__S
timestamp -25199
transform -1 0 8372 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__Y
timestamp -25199
transform -1 0 23552 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A1
timestamp -25199
transform 1 0 3128 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__S
timestamp -25199
transform 1 0 30728 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__S
timestamp -25199
transform 1 0 20884 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A1
timestamp -25199
transform -1 0 31556 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__S
timestamp -25199
transform 1 0 30728 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A1
timestamp -25199
transform 1 0 28888 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__S
timestamp -25199
transform 1 0 30360 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A1
timestamp -25199
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__S
timestamp -25199
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__S
timestamp -25199
transform 1 0 28980 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__S
timestamp -25199
transform 1 0 7820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__S
timestamp -25199
transform -1 0 14076 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__S
timestamp -25199
transform 1 0 11776 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__S
timestamp -25199
transform 1 0 23000 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__S
timestamp -25199
transform 1 0 10764 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__S
timestamp -25199
transform 1 0 17756 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__S
timestamp -25199
transform 1 0 7544 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__S
timestamp -25199
transform 1 0 22080 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__S
timestamp -25199
transform -1 0 8648 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__S
timestamp -25199
transform -1 0 22540 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__S
timestamp -25199
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__S
timestamp -25199
transform 1 0 12696 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__S
timestamp -25199
transform -1 0 24288 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__S
timestamp -25199
transform -1 0 12512 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__S
timestamp -25199
transform -1 0 19872 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__S
timestamp -25199
transform 1 0 14904 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__S
timestamp -25199
transform -1 0 11040 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A1
timestamp -25199
transform 1 0 11316 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__S
timestamp -25199
transform -1 0 12512 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__S
timestamp -25199
transform 1 0 17480 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__S
timestamp -25199
transform 1 0 27508 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__S
timestamp -25199
transform 1 0 15456 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__S
timestamp -25199
transform 1 0 27784 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__S
timestamp -25199
transform 1 0 11132 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__S
timestamp -25199
transform 1 0 23184 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__S
timestamp -25199
transform 1 0 15824 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A1
timestamp -25199
transform 1 0 26956 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__S
timestamp -25199
transform 1 0 17848 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A1
timestamp -25199
transform 1 0 25392 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__S
timestamp -25199
transform 1 0 15824 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__S
timestamp -25199
transform -1 0 19596 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__S
timestamp -25199
transform 1 0 13616 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__S
timestamp -25199
transform -1 0 4508 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A1
timestamp -25199
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__S
timestamp -25199
transform 1 0 4600 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__S
timestamp -25199
transform -1 0 18308 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__S
timestamp -25199
transform -1 0 24564 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__S
timestamp -25199
transform 1 0 3680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__S
timestamp -25199
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__S
timestamp -25199
transform 1 0 9752 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__S
timestamp -25199
transform -1 0 26128 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__S
timestamp -25199
transform 1 0 11224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__S
timestamp -25199
transform 1 0 24012 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__S
timestamp -25199
transform -1 0 18308 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__S
timestamp -25199
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__S
timestamp -25199
transform -1 0 24656 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__S
timestamp -25199
transform -1 0 4048 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__S
timestamp -25199
transform -1 0 18400 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__S
timestamp -25199
transform 1 0 6440 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__S
timestamp -25199
transform -1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__S
timestamp -25199
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__S
timestamp -25199
transform 1 0 7176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__S
timestamp -25199
transform 1 0 28244 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__S
timestamp -25199
transform -1 0 15732 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__S
timestamp -25199
transform 1 0 28612 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__S
timestamp -25199
transform 1 0 14444 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__S
timestamp -25199
transform 1 0 22080 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__S
timestamp -25199
transform 1 0 4968 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__S
timestamp -25199
transform 1 0 22632 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__S
timestamp -25199
transform 1 0 14904 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__S
timestamp -25199
transform 1 0 24932 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__S
timestamp -25199
transform 1 0 28244 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__S
timestamp -25199
transform 1 0 10212 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__S
timestamp -25199
transform 1 0 12880 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__S
timestamp -25199
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__S
timestamp -25199
transform -1 0 23828 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__S
timestamp -25199
transform 1 0 7176 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__S
timestamp -25199
transform 1 0 26036 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__S
timestamp -25199
transform 1 0 9200 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__S
timestamp -25199
transform 1 0 19044 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__S
timestamp -25199
transform 1 0 6900 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__S
timestamp -25199
transform 1 0 23828 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__S
timestamp -25199
transform 1 0 20148 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A1
timestamp -25199
transform 1 0 9936 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__S
timestamp -25199
transform 1 0 10948 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__S
timestamp -25199
transform 1 0 23644 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__S
timestamp -25199
transform 1 0 10948 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__S
timestamp -25199
transform 1 0 20056 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__S
timestamp -25199
transform 1 0 7084 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__RESET_B
timestamp -25199
transform 1 0 28152 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp -25199
transform 1 0 17940 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp -25199
transform 1 0 19964 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_clk_A
timestamp -25199
transform 1 0 13616 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_clk_X
timestamp -25199
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_clk_A
timestamp -25199
transform 1 0 13708 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_clk_X
timestamp -25199
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_clk_A
timestamp -25199
transform -1 0 24932 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_clk_X
timestamp -25199
transform 1 0 27140 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_clk_A
timestamp -25199
transform 1 0 24564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_clk_X
timestamp -25199
transform 1 0 26496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_clk_A
timestamp -25199
transform 1 0 4968 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_clk_A
timestamp -25199
transform 1 0 11408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_clk_A
timestamp -25199
transform 1 0 14260 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_clk_A
timestamp -25199
transform 1 0 9936 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_clk_A
timestamp -25199
transform 1 0 5152 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_clk_A
timestamp -25199
transform 1 0 6256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_clk_A
timestamp -25199
transform -1 0 7912 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_clk_A
timestamp -25199
transform 1 0 11132 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_clk_A
timestamp -25199
transform 1 0 15640 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_clk_A
timestamp -25199
transform 1 0 14168 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_clk_A
timestamp -25199
transform 1 0 17940 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_clk_A
timestamp -25199
transform 1 0 23000 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_12_clk_A
timestamp -25199
transform 1 0 23092 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_13_clk_A
timestamp -25199
transform 1 0 28612 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_14_clk_A
timestamp -25199
transform 1 0 30820 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_15_clk_A
timestamp -25199
transform -1 0 29532 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_16_clk_A
timestamp -25199
transform 1 0 26312 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_17_clk_A
timestamp -25199
transform 1 0 23920 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_18_clk_A
timestamp -25199
transform 1 0 29164 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_19_clk_A
timestamp -25199
transform 1 0 31924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_20_clk_A
timestamp -25199
transform 1 0 31004 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_21_clk_A
timestamp -25199
transform -1 0 29164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_22_clk_A
timestamp -25199
transform 1 0 22816 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_23_clk_A
timestamp -25199
transform 1 0 22908 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_24_clk_A
timestamp -25199
transform 1 0 15456 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_25_clk_A
timestamp -25199
transform 1 0 14536 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_26_clk_A
timestamp -25199
transform -1 0 14076 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_27_clk_A
timestamp -25199
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_28_clk_A
timestamp -25199
transform 1 0 7360 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload0_A
timestamp -25199
transform -1 0 12512 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload1_A
timestamp -25199
transform 1 0 23920 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload2_A
timestamp -25199
transform 1 0 25024 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout38_A
timestamp -25199
transform -1 0 26036 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout38_X
timestamp -25199
transform -1 0 26404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout39_A
timestamp -25199
transform 1 0 24012 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout39_X
timestamp -25199
transform -1 0 24564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout40_X
timestamp -25199
transform 1 0 23736 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout41_A
timestamp -25199
transform 1 0 15088 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout41_X
timestamp -25199
transform 1 0 14904 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout42_A
timestamp -25199
transform 1 0 5796 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout43_A
timestamp -25199
transform -1 0 22356 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout43_X
timestamp -25199
transform 1 0 22540 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout44_X
timestamp -25199
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout45_A
timestamp -25199
transform -1 0 4140 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout45_X
timestamp -25199
transform -1 0 4692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout46_A
timestamp -25199
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout46_X
timestamp -25199
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout47_X
timestamp -25199
transform -1 0 24840 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout48_A
timestamp -25199
transform -1 0 28060 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout48_X
timestamp -25199
transform -1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout49_A
timestamp -25199
transform 1 0 15732 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout49_X
timestamp -25199
transform 1 0 15548 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout50_A
timestamp -25199
transform -1 0 29256 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout51_X
timestamp -25199
transform -1 0 28244 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout52_A
timestamp -25199
transform -1 0 14536 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout52_X
timestamp -25199
transform 1 0 13708 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout53_A
timestamp -25199
transform 1 0 22448 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout53_X
timestamp -25199
transform 1 0 22264 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout54_X
timestamp -25199
transform 1 0 22172 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout55_A
timestamp -25199
transform -1 0 6900 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout56_A
timestamp -25199
transform 1 0 7452 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout57_A
timestamp -25199
transform -1 0 30452 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout57_X
timestamp -25199
transform 1 0 30452 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout58_A
timestamp -25199
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout58_X
timestamp -25199
transform 1 0 21804 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout59_A
timestamp -25199
transform 1 0 26312 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout60_A
timestamp -25199
transform -1 0 26864 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout60_X
timestamp -25199
transform 1 0 28244 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout61_A
timestamp -25199
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout61_X
timestamp -25199
transform 1 0 19412 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout62_A
timestamp -25199
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout62_X
timestamp -25199
transform -1 0 16652 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout63_X
timestamp -25199
transform -1 0 27140 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout64_A
timestamp -25199
transform -1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout64_X
timestamp -25199
transform -1 0 20608 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout65_A
timestamp -25199
transform 1 0 13708 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout65_X
timestamp -25199
transform 1 0 13524 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout66_X
timestamp -25199
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout67_A
timestamp -25199
transform 1 0 11500 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout67_X
timestamp -25199
transform 1 0 11316 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout68_A
timestamp -25199
transform 1 0 28428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout68_X
timestamp -25199
transform 1 0 28244 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout69_X
timestamp -25199
transform -1 0 28980 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout70_A
timestamp -25199
transform -1 0 18216 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout70_X
timestamp -25199
transform 1 0 17848 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout71_A
timestamp -25199
transform 1 0 30636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout72_A
timestamp -25199
transform 1 0 29532 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout72_X
timestamp -25199
transform 1 0 29348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout73_X
timestamp -25199
transform 1 0 29808 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout74_A
timestamp -25199
transform -1 0 25944 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout74_X
timestamp -25199
transform -1 0 25024 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout75_A
timestamp -25199
transform -1 0 23092 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout75_X
timestamp -25199
transform -1 0 22908 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout76_A
timestamp -25199
transform 1 0 27784 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout77_X
timestamp -25199
transform 1 0 25024 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout78_A
timestamp -25199
transform 1 0 25852 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout78_X
timestamp -25199
transform -1 0 26036 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout79_A
timestamp -25199
transform 1 0 26312 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout79_X
timestamp -25199
transform -1 0 28336 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout80_X
timestamp -25199
transform -1 0 26772 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout81_A
timestamp -25199
transform -1 0 18308 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout81_X
timestamp -25199
transform -1 0 19136 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout82_A
timestamp -25199
transform 1 0 22264 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout83_A
timestamp -25199
transform 1 0 20240 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout83_X
timestamp -25199
transform 1 0 20608 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout84_A
timestamp -25199
transform 1 0 18676 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout84_X
timestamp -25199
transform 1 0 18492 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout85_A
timestamp -25199
transform 1 0 27048 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout85_X
timestamp -25199
transform -1 0 28612 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout86_X
timestamp -25199
transform -1 0 29716 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout87_A
timestamp -25199
transform -1 0 22172 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout87_X
timestamp -25199
transform 1 0 22356 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout88_A
timestamp -25199
transform -1 0 31648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout88_X
timestamp -25199
transform -1 0 31832 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout89_A
timestamp -25199
transform -1 0 28704 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout90_X
timestamp -25199
transform 1 0 21988 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout91_X
timestamp -25199
transform -1 0 22816 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout92_X
timestamp -25199
transform 1 0 20516 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout95_A
timestamp -25199
transform 1 0 25300 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout95_X
timestamp -25199
transform -1 0 25300 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout96_A
timestamp -25199
transform 1 0 29348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout97_A
timestamp -25199
transform -1 0 27048 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout97_X
timestamp -25199
transform -1 0 26864 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout98_X
timestamp -25199
transform 1 0 28796 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout99_A
timestamp -25199
transform 1 0 20884 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout99_X
timestamp -25199
transform 1 0 20700 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout100_A
timestamp -25199
transform -1 0 31372 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout101_A
timestamp -25199
transform 1 0 29716 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout101_X
timestamp -25199
transform -1 0 30452 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout102_X
timestamp -25199
transform -1 0 31556 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout103_A
timestamp -25199
transform -1 0 28980 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout103_X
timestamp -25199
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout104_A
timestamp -25199
transform -1 0 27140 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout104_X
timestamp -25199
transform -1 0 27508 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout105_X
timestamp -25199
transform 1 0 24012 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout106_A
timestamp -25199
transform 1 0 16284 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout106_X
timestamp -25199
transform 1 0 15916 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout107_A
timestamp -25199
transform 1 0 16744 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout107_X
timestamp -25199
transform 1 0 16560 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout108_A
timestamp -25199
transform -1 0 26864 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout108_X
timestamp -25199
transform 1 0 26496 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout109_X
timestamp -25199
transform -1 0 27876 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout110_A
timestamp -25199
transform 1 0 25668 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout110_X
timestamp -25199
transform -1 0 25668 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout111_A
timestamp -25199
transform 1 0 24012 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout111_X
timestamp -25199
transform -1 0 24012 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout112_A
timestamp -25199
transform -1 0 29348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout113_X
timestamp -25199
transform 1 0 27968 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout114_A
timestamp -25199
transform 1 0 17112 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout114_X
timestamp -25199
transform -1 0 17112 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout115_A
timestamp -25199
transform 1 0 30544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout115_X
timestamp -25199
transform 1 0 30360 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout116_X
timestamp -25199
transform -1 0 31188 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout117_A
timestamp -25199
transform 1 0 23092 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout117_X
timestamp -25199
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout118_A
timestamp -25199
transform 1 0 28888 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout118_X
timestamp -25199
transform -1 0 28888 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout119_X
timestamp -25199
transform -1 0 29440 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout121_A
timestamp -25199
transform -1 0 33580 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout122_A
timestamp -25199
transform 1 0 32844 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout123_A
timestamp -25199
transform 1 0 34500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout124_A
timestamp -25199
transform -1 0 33028 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout125_X
timestamp -25199
transform 1 0 33212 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout126_A
timestamp -25199
transform -1 0 33856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout127_A
timestamp -25199
transform -1 0 32016 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout127_X
timestamp -25199
transform 1 0 32844 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout128_A
timestamp -25199
transform 1 0 29624 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout128_X
timestamp -25199
transform -1 0 29624 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout129_A
timestamp -25199
transform -1 0 29164 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout130_X
timestamp -25199
transform -1 0 32844 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout131_A
timestamp -25199
transform -1 0 10948 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout131_X
timestamp -25199
transform -1 0 10764 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout132_A
timestamp -25199
transform -1 0 26312 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout132_X
timestamp -25199
transform 1 0 26312 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout133_X
timestamp -25199
transform 1 0 23736 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout134_A
timestamp -25199
transform 1 0 26220 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout134_X
timestamp -25199
transform -1 0 26772 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout135_A
timestamp -25199
transform 1 0 25852 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout135_X
timestamp -25199
transform -1 0 25760 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout136_X
timestamp -25199
transform 1 0 26404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout137_A
timestamp -25199
transform 1 0 8188 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout138_A
timestamp -25199
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout139_A
timestamp -25199
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout139_X
timestamp -25199
transform 1 0 29072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout140_A
timestamp -25199
transform 1 0 19780 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout140_X
timestamp -25199
transform -1 0 19780 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout141_A
timestamp -25199
transform 1 0 16192 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout141_X
timestamp -25199
transform 1 0 16008 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout142_X
timestamp -25199
transform 1 0 23092 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout143_A
timestamp -25199
transform -1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout143_X
timestamp -25199
transform 1 0 26312 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout144_A
timestamp -25199
transform 1 0 20608 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout144_X
timestamp -25199
transform 1 0 20240 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout145_A
timestamp -25199
transform -1 0 28152 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout146_X
timestamp -25199
transform 1 0 22816 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout147_A
timestamp -25199
transform 1 0 15272 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout147_X
timestamp -25199
transform 1 0 15456 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout148_A
timestamp -25199
transform 1 0 5612 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout149_A
timestamp -25199
transform 1 0 27968 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout149_X
timestamp -25199
transform -1 0 31004 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout150_X
timestamp -25199
transform -1 0 29440 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout151_A
timestamp -25199
transform 1 0 31188 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout151_X
timestamp -25199
transform -1 0 31188 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout152_A
timestamp -25199
transform -1 0 32108 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout152_X
timestamp -25199
transform -1 0 31924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout153_X
timestamp -25199
transform -1 0 32936 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout154_A
timestamp -25199
transform -1 0 27876 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout154_X
timestamp -25199
transform -1 0 29348 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout155_A
timestamp -25199
transform 1 0 28336 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout155_X
timestamp -25199
transform 1 0 26128 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout156_X
timestamp -25199
transform -1 0 29348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout157_A
timestamp -25199
transform -1 0 28612 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout157_X
timestamp -25199
transform 1 0 28980 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout158_A
timestamp -25199
transform 1 0 28060 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout158_X
timestamp -25199
transform -1 0 28612 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout159_X
timestamp -25199
transform 1 0 24748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout192_A
timestamp -25199
transform 1 0 22816 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout194_A
timestamp -25199
transform -1 0 2944 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout195_X
timestamp -25199
transform -1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout206_A
timestamp -25199
transform 1 0 24932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout207_A
timestamp -25199
transform 1 0 32844 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout208_A
timestamp -25199
transform 1 0 24012 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout208_X
timestamp -25199
transform -1 0 24196 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout209_A
timestamp -25199
transform 1 0 31740 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout210_A
timestamp -25199
transform 1 0 33396 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout211_A
timestamp -25199
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout211_X
timestamp -25199
transform 1 0 22632 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout214_A
timestamp -25199
transform -1 0 23000 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout221_A
timestamp -25199
transform 1 0 19044 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout229_A
timestamp -25199
transform 1 0 18308 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout237_A
timestamp -25199
transform -1 0 21436 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout242_A
timestamp -25199
transform -1 0 19780 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout243_X
timestamp -25199
transform -1 0 3036 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp -25199
transform -1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_X
timestamp -25199
transform 1 0 1748 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp -25199
transform -1 0 2024 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_X
timestamp -25199
transform 1 0 1656 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp -25199
transform -1 0 1840 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp -25199
transform -1 0 1840 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp -25199
transform -1 0 1840 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp -25199
transform -1 0 1564 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_X
timestamp -25199
transform -1 0 2484 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp -25199
transform -1 0 1840 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp -25199
transform -1 0 1564 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp -25199
transform -1 0 2116 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp -25199
transform -1 0 1840 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp -25199
transform -1 0 1840 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp -25199
transform -1 0 2024 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_X
timestamp -25199
transform 1 0 1656 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp -25199
transform -1 0 1840 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp -25199
transform -1 0 2024 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_X
timestamp -25199
transform -1 0 1840 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp -25199
transform -1 0 1840 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp -25199
transform -1 0 2116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_X
timestamp -25199
transform 1 0 1748 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp -25199
transform -1 0 1840 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp -25199
transform -1 0 2116 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_X
timestamp -25199
transform 1 0 1748 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp -25199
transform -1 0 2116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_X
timestamp -25199
transform -1 0 1932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -25199
transform 1 0 18124 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp -25199
transform -1 0 13616 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp -25199
transform -1 0 13708 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp -25199
transform 1 0 24932 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp -25199
transform 1 0 24656 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_0_clk
timestamp -25199
transform -1 0 4968 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_1_clk
timestamp -25199
transform 1 0 10396 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_2_clk
timestamp -25199
transform -1 0 15456 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_3_clk
timestamp -25199
transform 1 0 8924 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_4_clk
timestamp -25199
transform -1 0 5152 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_5_clk
timestamp -25199
transform 1 0 5244 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_6_clk
timestamp -25199
transform 1 0 6348 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_7_clk
timestamp -25199
transform 1 0 10120 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_8_clk
timestamp -25199
transform 1 0 16192 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_9_clk
timestamp -25199
transform 1 0 14352 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_10_clk
timestamp -25199
transform 1 0 18124 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_11_clk
timestamp -25199
transform -1 0 22816 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_12_clk
timestamp -25199
transform -1 0 23092 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_13_clk
timestamp -25199
transform 1 0 28796 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_14_clk
timestamp -25199
transform 1 0 31004 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_15_clk
timestamp -25199
transform 1 0 29532 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_16_clk
timestamp -25199
transform 1 0 24472 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_17_clk
timestamp -25199
transform -1 0 23460 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_18_clk
timestamp -25199
transform 1 0 29256 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_19_clk
timestamp -25199
transform 1 0 32292 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_20_clk
timestamp -25199
transform 1 0 31188 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_21_clk
timestamp -25199
transform 1 0 29164 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_22_clk
timestamp -25199
transform -1 0 22816 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_23_clk
timestamp -25199
transform 1 0 21896 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_24_clk
timestamp -25199
transform 1 0 16468 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_25_clk
timestamp -25199
transform 1 0 14720 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_26_clk
timestamp -25199
transform 1 0 14076 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_27_clk
timestamp -25199
transform 1 0 6440 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_28_clk
timestamp -25199
transform 1 0 5980 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinvlp_4  clkload0
timestamp -25199
transform 1 0 11776 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkinvlp_4  clkload1
timestamp -25199
transform 1 0 24840 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_6  clkload2
timestamp -25199
transform 1 0 24012 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload3
timestamp -25199
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_6  clkload4
timestamp -25199
transform 1 0 16836 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload5
timestamp -25199
transform 1 0 15272 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_6  clkload6
timestamp -25199
transform 1 0 13248 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload7
timestamp -25199
transform 1 0 6440 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_2  clkload8
timestamp -25199
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  clkload9
timestamp -25199
transform 1 0 15456 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_2  clkload10
timestamp -25199
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  clkload11
timestamp -25199
transform 1 0 4140 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload12
timestamp -25199
transform 1 0 5428 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_6  clkload13
timestamp -25199
transform 1 0 6256 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  clkload14
timestamp -25199
transform 1 0 15824 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  clkload15
timestamp -25199
transform 1 0 14812 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__bufinv_16  clkload16
timestamp -25199
transform 1 0 19228 0 1 22848
box -38 -48 2246 592
use sky130_fd_sc_hd__bufinv_16  clkload17
timestamp -25199
transform 1 0 22080 0 1 17408
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinvlp_4  clkload18
timestamp -25199
transform 1 0 29532 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_4  clkload19
timestamp -25199
transform 1 0 33304 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_4  clkload20
timestamp -25199
transform 1 0 30728 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_6  clkload21
timestamp -25199
transform 1 0 29532 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload22
timestamp -25199
transform 1 0 21804 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload23
timestamp -25199
transform 1 0 22540 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  clkload24
timestamp -25199
transform 1 0 29808 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_6  clkload25
timestamp -25199
transform 1 0 31096 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload26
timestamp -25199
transform 1 0 30912 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload27
timestamp -25199
transform 1 0 24104 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout38
timestamp -25199
transform 1 0 25116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp -25199
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp -25199
transform 1 0 23368 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp -25199
transform 1 0 14536 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout42
timestamp -25199
transform -1 0 5796 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout43
timestamp -25199
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp -25199
transform -1 0 21436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp -25199
transform 1 0 4140 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout46
timestamp -25199
transform 1 0 23736 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout47
timestamp -25199
transform 1 0 24104 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout48
timestamp -25199
transform 1 0 27876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout49
timestamp -25199
transform -1 0 15548 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout50
timestamp -25199
transform -1 0 28980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout51
timestamp -25199
transform 1 0 27508 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout52
timestamp -25199
transform -1 0 14260 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout53
timestamp -25199
transform 1 0 21896 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp -25199
transform -1 0 22172 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout55
timestamp -25199
transform -1 0 6716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout56
timestamp -25199
transform 1 0 6532 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout57
timestamp -25199
transform 1 0 29532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout58
timestamp -25199
transform -1 0 21252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout59
timestamp -25199
transform -1 0 26864 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout60
timestamp -25199
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout61
timestamp -25199
transform -1 0 19044 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout62
timestamp -25199
transform -1 0 16284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout63
timestamp -25199
transform 1 0 25852 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout64
timestamp -25199
transform 1 0 19872 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout65
timestamp -25199
transform -1 0 13524 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout66
timestamp -25199
transform -1 0 20608 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout67
timestamp -25199
transform -1 0 11316 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout68
timestamp -25199
transform 1 0 27324 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout69
timestamp -25199
transform 1 0 27692 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout70
timestamp -25199
transform -1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout71
timestamp -25199
transform 1 0 29532 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout72
timestamp -25199
transform -1 0 29348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout73
timestamp -25199
transform 1 0 29440 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout74
timestamp -25199
transform 1 0 24288 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout75
timestamp -25199
transform -1 0 21988 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout76
timestamp -25199
transform 1 0 27968 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout77
timestamp -25199
transform -1 0 24840 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout78
timestamp -25199
transform 1 0 25024 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout79
timestamp -25199
transform 1 0 26496 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout80
timestamp -25199
transform 1 0 25392 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout81
timestamp -25199
transform 1 0 18584 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout82
timestamp -25199
transform -1 0 22172 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout83
timestamp -25199
transform -1 0 20240 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout84
timestamp -25199
transform -1 0 18492 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout85
timestamp -25199
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout86
timestamp -25199
transform 1 0 28612 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout87
timestamp -25199
transform 1 0 21988 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout88
timestamp -25199
transform -1 0 31464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout89
timestamp -25199
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout90
timestamp -25199
transform 1 0 21620 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout91
timestamp -25199
transform -1 0 21712 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout92
timestamp -25199
transform 1 0 20148 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout93
timestamp -25199
transform -1 0 20148 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout94
timestamp -25199
transform 1 0 24380 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout95
timestamp -25199
transform -1 0 24748 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout96
timestamp -25199
transform -1 0 29808 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout97
timestamp -25199
transform 1 0 25944 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout98
timestamp -25199
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout99
timestamp -25199
transform -1 0 20700 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout100
timestamp -25199
transform -1 0 31004 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout101
timestamp -25199
transform 1 0 29900 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout102
timestamp -25199
transform 1 0 30360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout103
timestamp -25199
transform 1 0 28428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout104
timestamp -25199
transform 1 0 26588 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout105
timestamp -25199
transform -1 0 24012 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout106
timestamp -25199
transform -1 0 15916 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout107
timestamp -25199
transform -1 0 16560 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout108
timestamp -25199
transform 1 0 26128 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout109
timestamp -25199
transform 1 0 26864 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout110
timestamp -25199
transform -1 0 25116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout111
timestamp -25199
transform -1 0 23000 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout112
timestamp -25199
transform -1 0 29440 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout113
timestamp -25199
transform 1 0 26864 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout114
timestamp -25199
transform 1 0 16560 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout115
timestamp -25199
transform 1 0 29992 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout116
timestamp -25199
transform 1 0 29808 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout117
timestamp -25199
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout118
timestamp -25199
transform 1 0 27968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout119
timestamp -25199
transform 1 0 28336 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout120
timestamp -25199
transform -1 0 33028 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout121
timestamp -25199
transform 1 0 33304 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout122
timestamp -25199
transform -1 0 32844 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout123
timestamp -25199
transform -1 0 35052 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout124
timestamp -25199
transform -1 0 33304 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout125
timestamp -25199
transform -1 0 33212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout126
timestamp -25199
transform -1 0 33304 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout127
timestamp -25199
transform 1 0 32476 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout128
timestamp -25199
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout129
timestamp -25199
transform -1 0 28980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout130
timestamp -25199
transform 1 0 32108 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout131
timestamp -25199
transform 1 0 10212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout132
timestamp -25199
transform 1 0 25576 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout133
timestamp -25199
transform -1 0 24288 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout134
timestamp -25199
transform -1 0 25668 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout135
timestamp -25199
transform 1 0 24656 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout136
timestamp -25199
transform 1 0 25484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout137
timestamp -25199
transform -1 0 8188 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout138
timestamp -25199
transform 1 0 8556 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout139
timestamp -25199
transform 1 0 28888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout140
timestamp -25199
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout141
timestamp -25199
transform -1 0 16008 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout142
timestamp -25199
transform -1 0 22356 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout143
timestamp -25199
transform 1 0 27508 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout144
timestamp -25199
transform -1 0 20240 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout145
timestamp -25199
transform -1 0 27968 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout146
timestamp -25199
transform -1 0 22816 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout147
timestamp -25199
transform 1 0 14720 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout148
timestamp -25199
transform 1 0 5336 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout149
timestamp -25199
transform 1 0 28980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout150
timestamp -25199
transform 1 0 28612 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout151
timestamp -25199
transform -1 0 30820 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout152
timestamp -25199
transform 1 0 31188 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout153
timestamp -25199
transform 1 0 31556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout154
timestamp -25199
transform 1 0 27140 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout155
timestamp -25199
transform 1 0 26036 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout156
timestamp -25199
transform 1 0 27600 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout157
timestamp -25199
transform -1 0 28244 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout158
timestamp -25199
transform 1 0 27692 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout159
timestamp -25199
transform -1 0 24748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout160
timestamp -25199
transform -1 0 29716 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout161
timestamp -25199
transform 1 0 23736 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout162
timestamp -25199
transform -1 0 23552 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout163
timestamp -25199
transform -1 0 23644 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout164
timestamp -25199
transform -1 0 24104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout165
timestamp -25199
transform -1 0 27692 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout166
timestamp -25199
transform 1 0 30084 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout167
timestamp -25199
transform -1 0 25668 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout168
timestamp -25199
transform -1 0 27600 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout169
timestamp -25199
transform 1 0 30452 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout170
timestamp -25199
transform -1 0 30820 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout171
timestamp -25199
transform 1 0 26036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout172
timestamp -25199
transform -1 0 28060 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout173
timestamp -25199
transform -1 0 32016 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout174
timestamp -25199
transform -1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout175
timestamp -25199
transform -1 0 26680 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout176
timestamp -25199
transform -1 0 28428 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout177
timestamp -25199
transform 1 0 32384 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  fanout178
timestamp -25199
transform -1 0 32384 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout179
timestamp -25199
transform 1 0 6348 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout180
timestamp -25199
transform -1 0 13892 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout181
timestamp -25199
transform 1 0 5336 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout182
timestamp -25199
transform 1 0 18768 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout183
timestamp -25199
transform 1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout184
timestamp -25199
transform 1 0 18492 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout185
timestamp -25199
transform 1 0 18768 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout186
timestamp -25199
transform -1 0 4692 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout187
timestamp -25199
transform 1 0 10396 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout188
timestamp -25199
transform 1 0 15548 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout189
timestamp -25199
transform 1 0 4048 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout190
timestamp -25199
transform -1 0 23276 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout191
timestamp -25199
transform 1 0 23552 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout192
timestamp -25199
transform 1 0 23276 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout193
timestamp -25199
transform -1 0 3588 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout194
timestamp -25199
transform -1 0 4232 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout195
timestamp -25199
transform 1 0 2944 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout196
timestamp -25199
transform 1 0 17480 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout197
timestamp -25199
transform -1 0 17480 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout198
timestamp -25199
transform 1 0 14352 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout199
timestamp -25199
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout200
timestamp -25199
transform 1 0 5336 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout201
timestamp -25199
transform 1 0 9292 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout202
timestamp -25199
transform 1 0 4968 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout203
timestamp -25199
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout204
timestamp -25199
transform 1 0 23460 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout205
timestamp -25199
transform -1 0 31280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout206
timestamp -25199
transform -1 0 23460 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout207
timestamp -25199
transform 1 0 33028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout208
timestamp -25199
transform -1 0 23736 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout209
timestamp -25199
transform 1 0 31924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout210
timestamp -25199
transform 1 0 34132 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout211
timestamp -25199
transform 1 0 22264 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout212
timestamp -25199
transform -1 0 21712 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout213
timestamp -25199
transform -1 0 26036 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout214
timestamp -25199
transform 1 0 22356 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout215
timestamp -25199
transform 1 0 3772 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout216
timestamp -25199
transform -1 0 8372 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout217
timestamp -25199
transform -1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout218
timestamp -25199
transform 1 0 4692 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout219
timestamp -25199
transform 1 0 18308 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout220
timestamp -25199
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout221
timestamp -25199
transform 1 0 19228 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout222
timestamp -25199
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout223
timestamp -25199
transform -1 0 12420 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout224
timestamp -25199
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout225
timestamp -25199
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout226
timestamp -25199
transform 1 0 18952 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout227
timestamp -25199
transform 1 0 22172 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout228
timestamp -25199
transform 1 0 27232 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout229
timestamp -25199
transform 1 0 18492 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout230
timestamp -25199
transform 1 0 3680 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout231
timestamp -25199
transform -1 0 11224 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout232
timestamp -25199
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout233
timestamp -25199
transform 1 0 3404 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout234
timestamp -25199
transform 1 0 21896 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout235
timestamp -25199
transform 1 0 27048 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout236
timestamp -25199
transform -1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout237
timestamp -25199
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout238
timestamp -25199
transform -1 0 12420 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout239
timestamp -25199
transform 1 0 16560 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout240
timestamp -25199
transform 1 0 3404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout241
timestamp -25199
transform 1 0 12604 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout242
timestamp -25199
transform 1 0 19780 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout243
timestamp -25199
transform 1 0 3036 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636943256
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636943256
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -25199
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636943256
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636943256
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -25199
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636943256
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636943256
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -25199
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636943256
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636943256
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -25199
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636943256
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636943256
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -25199
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636943256
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636943256
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -25199
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636943256
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636943256
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -25199
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636943256
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636943256
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -25199
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636943256
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636943256
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -25199
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636943256
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636943256
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -25199
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636943256
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636943256
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -25199
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636943256
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1636943256
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp -25199
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1636943256
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1636943256
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp -25199
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_365
timestamp -25199
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636943256
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636943256
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636943256
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636943256
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp -25199
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -25199
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636943256
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636943256
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636943256
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636943256
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp -25199
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -25199
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636943256
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636943256
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636943256
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636943256
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp -25199
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -25199
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636943256
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636943256
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636943256
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636943256
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp -25199
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp -25199
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636943256
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636943256
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636943256
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636943256
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp -25199
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp -25199
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636943256
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636943256
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636943256
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636943256
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp -25199
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp -25199
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636943256
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636943256
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_361
timestamp -25199
transform 1 0 34316 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_10
timestamp 1636943256
transform 1 0 2024 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_22
timestamp -25199
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636943256
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636943256
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636943256
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636943256
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp -25199
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -25199
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636943256
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636943256
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636943256
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636943256
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp -25199
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -25199
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636943256
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636943256
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636943256
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636943256
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp -25199
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp -25199
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636943256
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636943256
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636943256
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636943256
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp -25199
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp -25199
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636943256
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636943256
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636943256
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636943256
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp -25199
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp -25199
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_309
timestamp -25199
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636943256
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636943256
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636943256
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_357
timestamp -25199
transform 1 0 33948 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_365
timestamp -25199
transform 1 0 34684 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636943256
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636943256
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636943256
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636943256
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp -25199
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -25199
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636943256
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636943256
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636943256
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636943256
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp -25199
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -25199
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636943256
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636943256
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636943256
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636943256
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp -25199
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -25199
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636943256
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636943256
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636943256
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636943256
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp -25199
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp -25199
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_225
timestamp -25199
transform 1 0 21804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_231
timestamp -25199
transform 1 0 22356 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_239
timestamp 1636943256
transform 1 0 23092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_251
timestamp 1636943256
transform 1 0 24196 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_263
timestamp 1636943256
transform 1 0 25300 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_275
timestamp -25199
transform 1 0 26404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp -25199
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636943256
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_293
timestamp -25199
transform 1 0 28060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_328
timestamp -25199
transform 1 0 31280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_337
timestamp -25199
transform 1 0 32108 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_350
timestamp 1636943256
transform 1 0 33304 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_362
timestamp -25199
transform 1 0 34408 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_368
timestamp -25199
transform 1 0 34960 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636943256
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636943256
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -25199
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636943256
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636943256
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636943256
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636943256
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp -25199
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -25199
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636943256
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636943256
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636943256
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636943256
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp -25199
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp -25199
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636943256
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636943256
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636943256
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636943256
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp -25199
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp -25199
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636943256
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636943256
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_221
timestamp -25199
transform 1 0 21436 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_229
timestamp -25199
transform 1 0 22172 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636943256
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636943256
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636943256
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1636943256
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp -25199
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp -25199
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_309
timestamp -25199
transform 1 0 29532 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_324
timestamp -25199
transform 1 0 30912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_341
timestamp -25199
transform 1 0 32476 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_365
timestamp -25199
transform 1 0 34684 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_11
timestamp 1636943256
transform 1 0 2116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_23
timestamp 1636943256
transform 1 0 3220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_35
timestamp 1636943256
transform 1 0 4324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp -25199
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp -25199
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636943256
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636943256
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636943256
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636943256
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp -25199
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -25199
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636943256
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636943256
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636943256
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636943256
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp -25199
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -25199
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636943256
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636943256
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636943256
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636943256
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp -25199
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp -25199
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_225
timestamp -25199
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_233
timestamp -25199
transform 1 0 22540 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_245
timestamp -25199
transform 1 0 23644 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_275
timestamp -25199
transform 1 0 26404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp -25199
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636943256
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636943256
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636943256
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_317
timestamp -25199
transform 1 0 30268 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_325
timestamp -25199
transform 1 0 31004 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_333
timestamp -25199
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636943256
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_349
timestamp -25199
transform 1 0 33212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_353
timestamp -25199
transform 1 0 33580 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_356
timestamp -25199
transform 1 0 33856 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636943256
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636943256
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -25199
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636943256
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636943256
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636943256
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636943256
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp -25199
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp -25199
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636943256
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636943256
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636943256
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636943256
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp -25199
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp -25199
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636943256
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636943256
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636943256
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636943256
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp -25199
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp -25199
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636943256
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_209
timestamp -25199
transform 1 0 20332 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_217
timestamp -25199
transform 1 0 21068 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_238
timestamp -25199
transform 1 0 23000 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp -25199
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636943256
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636943256
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_277
timestamp -25199
transform 1 0 26588 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_281
timestamp -25199
transform 1 0 26956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_302
timestamp -25199
transform 1 0 28888 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_305
timestamp -25199
transform 1 0 29164 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_331
timestamp 1636943256
transform 1 0 31556 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_343
timestamp -25199
transform 1 0 32660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp -25199
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_365
timestamp -25199
transform 1 0 34684 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636943256
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636943256
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636943256
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636943256
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp -25199
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -25199
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636943256
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636943256
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636943256
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636943256
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp -25199
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp -25199
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636943256
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636943256
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_137
timestamp -25199
transform 1 0 13708 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_141
timestamp -25199
transform 1 0 14076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_153
timestamp 1636943256
transform 1 0 15180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp -25199
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636943256
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636943256
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636943256
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1636943256
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_232
timestamp -25199
transform 1 0 22448 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_261
timestamp -25199
transform 1 0 25116 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp -25199
transform 1 0 25852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp -25199
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636943256
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_293
timestamp -25199
transform 1 0 28060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_323
timestamp -25199
transform 1 0 30820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_333
timestamp -25199
transform 1 0 31740 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_355
timestamp 1636943256
transform 1 0 33764 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_367
timestamp -25199
transform 1 0 34868 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636943256
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636943256
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -25199
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636943256
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636943256
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636943256
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636943256
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp -25199
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp -25199
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636943256
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_108
timestamp -25199
transform 1 0 11040 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_124
timestamp 1636943256
transform 1 0 12512 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp -25199
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_157
timestamp -25199
transform 1 0 15548 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_177
timestamp -25199
transform 1 0 17388 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_181
timestamp -25199
transform 1 0 17756 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp -25199
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp -25199
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_205
timestamp -25199
transform 1 0 19964 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp -25199
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_268
timestamp -25199
transform 1 0 25760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_291
timestamp -25199
transform 1 0 27876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp -25199
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_316
timestamp -25199
transform 1 0 30176 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_322
timestamp -25199
transform 1 0 30728 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_329
timestamp -25199
transform 1 0 31372 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp -25199
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_365
timestamp -25199
transform 1 0 34684 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_11
timestamp 1636943256
transform 1 0 2116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_23
timestamp 1636943256
transform 1 0 3220 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_35
timestamp 1636943256
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp -25199
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -25199
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp -25199
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp -25199
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_129
timestamp -25199
transform 1 0 12972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_133
timestamp -25199
transform 1 0 13340 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_141
timestamp -25199
transform 1 0 14076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_153
timestamp 1636943256
transform 1 0 15180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp -25199
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_169
timestamp -25199
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_218
timestamp -25199
transform 1 0 21160 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_229
timestamp -25199
transform 1 0 22172 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_245
timestamp -25199
transform 1 0 23644 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp -25199
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636943256
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp -25199
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_299
timestamp -25199
transform 1 0 28612 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_303
timestamp -25199
transform 1 0 28980 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_309
timestamp 1636943256
transform 1 0 29532 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_321
timestamp -25199
transform 1 0 30636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_332
timestamp -25199
transform 1 0 31648 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636943256
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636943256
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -25199
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636943256
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636943256
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_53
timestamp -25199
transform 1 0 5980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_57
timestamp -25199
transform 1 0 6348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_78
timestamp -25199
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_96
timestamp 1636943256
transform 1 0 9936 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_108
timestamp 1636943256
transform 1 0 11040 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_120
timestamp -25199
transform 1 0 12144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_131
timestamp -25199
transform 1 0 13156 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp -25199
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_152
timestamp 1636943256
transform 1 0 15088 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_164
timestamp -25199
transform 1 0 16192 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_188
timestamp -25199
transform 1 0 18400 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_197
timestamp -25199
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_203
timestamp -25199
transform 1 0 19780 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_231
timestamp -25199
transform 1 0 22356 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp -25199
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1636943256
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1636943256
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_277
timestamp -25199
transform 1 0 26588 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_281
timestamp -25199
transform 1 0 26956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_293
timestamp 1636943256
transform 1 0 28060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_305
timestamp -25199
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_329
timestamp -25199
transform 1 0 31372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_333
timestamp -25199
transform 1 0 31740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_347
timestamp -25199
transform 1 0 33028 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_351
timestamp -25199
transform 1 0 33396 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_357
timestamp -25199
transform 1 0 33948 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_365
timestamp -25199
transform 1 0 34684 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636943256
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636943256
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_27
timestamp -25199
transform 1 0 3588 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1636943256
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp -25199
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp -25199
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp -25199
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_71
timestamp 1636943256
transform 1 0 7636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_83
timestamp 1636943256
transform 1 0 8740 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_106
timestamp -25199
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp -25199
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_132
timestamp -25199
transform 1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_195
timestamp -25199
transform 1 0 19044 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_203
timestamp -25199
transform 1 0 19780 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_229
timestamp -25199
transform 1 0 22172 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_233
timestamp -25199
transform 1 0 22540 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_244
timestamp 1636943256
transform 1 0 23552 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_256
timestamp 1636943256
transform 1 0 24656 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_268
timestamp 1636943256
transform 1 0 25760 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_301
timestamp 1636943256
transform 1 0 28796 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_313
timestamp -25199
transform 1 0 29900 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_324
timestamp 1636943256
transform 1 0 30912 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_357
timestamp -25199
transform 1 0 33948 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_8
timestamp 1636943256
transform 1 0 1840 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp -25199
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_63
timestamp -25199
transform 1 0 6900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_67
timestamp -25199
transform 1 0 7268 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp -25199
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp -25199
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_112
timestamp 1636943256
transform 1 0 11408 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_124
timestamp -25199
transform 1 0 12512 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp -25199
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp -25199
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_155
timestamp 1636943256
transform 1 0 15364 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_167
timestamp 1636943256
transform 1 0 16468 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_179
timestamp -25199
transform 1 0 17572 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp -25199
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_240
timestamp 1636943256
transform 1 0 23184 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_263
timestamp -25199
transform 1 0 25300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp -25199
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_311
timestamp 1636943256
transform 1 0 29716 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_323
timestamp 1636943256
transform 1 0 30820 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_335
timestamp -25199
transform 1 0 31924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_343
timestamp -25199
transform 1 0 32660 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_365
timestamp -25199
transform 1 0 34684 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636943256
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_46
timestamp -25199
transform 1 0 5336 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_61
timestamp -25199
transform 1 0 6716 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_78
timestamp -25199
transform 1 0 8280 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_95
timestamp -25199
transform 1 0 9844 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp -25199
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_130
timestamp -25199
transform 1 0 13064 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_138
timestamp -25199
transform 1 0 13800 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_141
timestamp -25199
transform 1 0 14076 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_154
timestamp 1636943256
transform 1 0 15272 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp -25199
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_171
timestamp -25199
transform 1 0 16836 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1636943256
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_205
timestamp -25199
transform 1 0 19964 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp -25199
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_227
timestamp -25199
transform 1 0 21988 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_235
timestamp -25199
transform 1 0 22724 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_244
timestamp -25199
transform 1 0 23552 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_269
timestamp -25199
transform 1 0 25852 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_273
timestamp -25199
transform 1 0 26220 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_324
timestamp -25199
transform 1 0 30912 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_327
timestamp -25199
transform 1 0 31188 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp -25199
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1636943256
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_349
timestamp -25199
transform 1 0 33212 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_355
timestamp -25199
transform 1 0 33764 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_362
timestamp -25199
transform 1 0 34408 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_368
timestamp -25199
transform 1 0 34960 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636943256
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_15
timestamp -25199
transform 1 0 2484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_21
timestamp -25199
transform 1 0 3036 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_24
timestamp -25199
transform 1 0 3312 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_49
timestamp -25199
transform 1 0 5612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_53
timestamp -25199
transform 1 0 5980 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_63
timestamp -25199
transform 1 0 6900 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp -25199
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp -25199
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_92
timestamp -25199
transform 1 0 9568 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_150
timestamp -25199
transform 1 0 14904 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_158
timestamp -25199
transform 1 0 15640 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_184
timestamp -25199
transform 1 0 18032 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp -25199
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1636943256
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_225
timestamp -25199
transform 1 0 21804 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_233
timestamp -25199
transform 1 0 22540 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_247
timestamp -25199
transform 1 0 23828 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp -25199
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_256
timestamp 1636943256
transform 1 0 24656 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_268
timestamp -25199
transform 1 0 25760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_276
timestamp -25199
transform 1 0 26496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp -25199
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_321
timestamp -25199
transform 1 0 30636 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_338
timestamp 1636943256
transform 1 0 32200 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_350
timestamp 1636943256
transform 1 0 33304 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp -25199
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_365
timestamp -25199
transform 1 0 34684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp -25199
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp -25199
transform 1 0 1748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_40
timestamp -25199
transform 1 0 4784 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp -25199
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636943256
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1636943256
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1636943256
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_93
timestamp -25199
transform 1 0 9660 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_101
timestamp -25199
transform 1 0 10396 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_105
timestamp -25199
transform 1 0 10764 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1636943256
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_130
timestamp -25199
transform 1 0 13064 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_136
timestamp -25199
transform 1 0 13616 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_143
timestamp -25199
transform 1 0 14260 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_188
timestamp -25199
transform 1 0 18400 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_235
timestamp 1636943256
transform 1 0 22724 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_247
timestamp 1636943256
transform 1 0 23828 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_270
timestamp -25199
transform 1 0 25944 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp -25199
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_322
timestamp 1636943256
transform 1 0 30728 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp -25199
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1636943256
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_8
timestamp -25199
transform 1 0 1840 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_16
timestamp -25199
transform 1 0 2576 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_25
timestamp -25199
transform 1 0 3404 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_38
timestamp -25199
transform 1 0 4600 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_70
timestamp -25199
transform 1 0 7544 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp -25199
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp -25199
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_89
timestamp -25199
transform 1 0 9292 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_106
timestamp -25199
transform 1 0 10856 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_118
timestamp -25199
transform 1 0 11960 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp -25199
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_144
timestamp -25199
transform 1 0 14352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_177
timestamp -25199
transform 1 0 17388 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_180
timestamp -25199
transform 1 0 17664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp -25199
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp -25199
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_206
timestamp -25199
transform 1 0 20056 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_214
timestamp -25199
transform 1 0 20792 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_223
timestamp -25199
transform 1 0 21620 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_238
timestamp 1636943256
transform 1 0 23000 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp -25199
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_271
timestamp -25199
transform 1 0 26036 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_295
timestamp -25199
transform 1 0 28244 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp -25199
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_323
timestamp 1636943256
transform 1 0 30820 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_335
timestamp 1636943256
transform 1 0 31924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_347
timestamp -25199
transform 1 0 33028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_355
timestamp -25199
transform 1 0 33764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp -25199
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_365
timestamp -25199
transform 1 0 34684 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636943256
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp -25199
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp -25199
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp -25199
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_61
timestamp -25199
transform 1 0 6716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_113
timestamp -25199
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_132
timestamp -25199
transform 1 0 13248 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_142
timestamp -25199
transform 1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_146
timestamp -25199
transform 1 0 14536 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp -25199
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_178
timestamp -25199
transform 1 0 17480 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_195
timestamp 1636943256
transform 1 0 19044 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_218
timestamp -25199
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_241
timestamp -25199
transform 1 0 23276 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp -25199
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_281
timestamp -25199
transform 1 0 26956 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_291
timestamp -25199
transform 1 0 27876 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_314
timestamp -25199
transform 1 0 29992 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp -25199
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1636943256
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1636943256
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_361
timestamp -25199
transform 1 0 34316 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636943256
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636943256
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp -25199
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636943256
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636943256
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_87
timestamp 1636943256
transform 1 0 9108 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_99
timestamp 1636943256
transform 1 0 10212 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_111
timestamp 1636943256
transform 1 0 11316 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_134
timestamp -25199
transform 1 0 13432 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1636943256
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1636943256
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1636943256
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1636943256
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp -25199
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_201
timestamp -25199
transform 1 0 19596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp -25199
transform 1 0 21252 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_224
timestamp -25199
transform 1 0 21712 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_271
timestamp -25199
transform 1 0 26036 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_282
timestamp -25199
transform 1 0 27048 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_297
timestamp -25199
transform 1 0 28428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_305
timestamp -25199
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_309
timestamp -25199
transform 1 0 29532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_328
timestamp -25199
transform 1 0 31280 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_339
timestamp -25199
transform 1 0 32292 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_351
timestamp 1636943256
transform 1 0 33396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp -25199
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_365
timestamp -25199
transform 1 0 34684 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_8
timestamp 1636943256
transform 1 0 1840 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_40
timestamp 1636943256
transform 1 0 4784 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp -25199
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_70
timestamp 1636943256
transform 1 0 7544 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1636943256
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp -25199
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp -25199
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1636943256
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1636943256
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp -25199
transform 1 0 15180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_157
timestamp -25199
transform 1 0 15548 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp -25199
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_182
timestamp -25199
transform 1 0 17848 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_207
timestamp -25199
transform 1 0 20148 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_225
timestamp -25199
transform 1 0 21804 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_262
timestamp -25199
transform 1 0 25208 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp -25199
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_303
timestamp 1636943256
transform 1 0 28980 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_315
timestamp 1636943256
transform 1 0 30084 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_327
timestamp -25199
transform 1 0 31188 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp -25199
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_357
timestamp -25199
transform 1 0 33948 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp -25199
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_11
timestamp -25199
transform 1 0 2116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_45
timestamp -25199
transform 1 0 5244 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_64
timestamp -25199
transform 1 0 6992 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_96
timestamp -25199
transform 1 0 9936 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_118
timestamp -25199
transform 1 0 11960 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_126
timestamp -25199
transform 1 0 12696 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp -25199
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_171
timestamp -25199
transform 1 0 16836 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_175
timestamp -25199
transform 1 0 17204 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp -25199
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_191
timestamp -25199
transform 1 0 18676 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp -25199
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_208
timestamp -25199
transform 1 0 20240 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_239
timestamp -25199
transform 1 0 23092 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_247
timestamp -25199
transform 1 0 23828 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp -25199
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_255
timestamp -25199
transform 1 0 24564 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1636943256
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1636943256
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1636943256
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1636943256
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp -25199
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp -25199
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_365
timestamp -25199
transform 1 0 34684 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636943256
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_15
timestamp -25199
transform 1 0 2484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_23
timestamp -25199
transform 1 0 3220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_28
timestamp -25199
transform 1 0 3680 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_34
timestamp -25199
transform 1 0 4232 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_44
timestamp 1636943256
transform 1 0 5152 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_77
timestamp 1636943256
transform 1 0 8188 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp -25199
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp -25199
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_150
timestamp 1636943256
transform 1 0 14904 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_162
timestamp -25199
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_169
timestamp -25199
transform 1 0 16652 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_186
timestamp -25199
transform 1 0 18216 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_203
timestamp 1636943256
transform 1 0 19780 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_215
timestamp -25199
transform 1 0 20884 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp -25199
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_283
timestamp -25199
transform 1 0 27140 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_291
timestamp -25199
transform 1 0 27876 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_310
timestamp -25199
transform 1 0 29624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_327
timestamp -25199
transform 1 0 31188 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp -25199
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1636943256
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1636943256
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_361
timestamp -25199
transform 1 0 34316 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636943256
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636943256
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp -25199
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636943256
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_41
timestamp -25199
transform 1 0 4876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_45
timestamp -25199
transform 1 0 5244 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_62
timestamp 1636943256
transform 1 0 6808 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_74
timestamp -25199
transform 1 0 7912 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp -25199
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp -25199
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp -25199
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_104
timestamp -25199
transform 1 0 10672 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_129
timestamp -25199
transform 1 0 12972 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp -25199
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_141
timestamp -25199
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_174
timestamp 1636943256
transform 1 0 17112 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_186
timestamp -25199
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp -25199
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp -25199
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_215
timestamp -25199
transform 1 0 20884 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_221
timestamp -25199
transform 1 0 21436 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_226
timestamp -25199
transform 1 0 21896 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_234
timestamp -25199
transform 1 0 22632 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_275
timestamp -25199
transform 1 0 26404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp -25199
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_313
timestamp -25199
transform 1 0 29900 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_327
timestamp 1636943256
transform 1 0 31188 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_339
timestamp 1636943256
transform 1 0 32292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_351
timestamp -25199
transform 1 0 33396 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp -25199
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_365
timestamp -25199
transform 1 0 34684 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_10
timestamp -25199
transform 1 0 2024 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_18
timestamp -25199
transform 1 0 2760 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_30
timestamp -25199
transform 1 0 3864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_44
timestamp -25199
transform 1 0 5152 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp -25199
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_57
timestamp -25199
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_65
timestamp -25199
transform 1 0 7084 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_84
timestamp 1636943256
transform 1 0 8832 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_107
timestamp -25199
transform 1 0 10948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_119
timestamp -25199
transform 1 0 12052 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_131
timestamp -25199
transform 1 0 13156 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_139
timestamp -25199
transform 1 0 13892 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_157
timestamp -25199
transform 1 0 15548 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_163
timestamp -25199
transform 1 0 16100 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_180
timestamp -25199
transform 1 0 17664 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_192
timestamp 1636943256
transform 1 0 18768 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_204
timestamp -25199
transform 1 0 19872 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_236
timestamp -25199
transform 1 0 22816 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_303
timestamp -25199
transform 1 0 28980 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp -25199
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_346
timestamp -25199
transform 1 0 32936 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp -25199
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_11
timestamp -25199
transform 1 0 2116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_65
timestamp -25199
transform 1 0 7084 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_73
timestamp -25199
transform 1 0 7820 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp -25199
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_89
timestamp -25199
transform 1 0 9292 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_114
timestamp -25199
transform 1 0 11592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp -25199
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp -25199
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1636943256
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_153
timestamp -25199
transform 1 0 15180 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp -25199
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_205
timestamp -25199
transform 1 0 19964 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_217
timestamp -25199
transform 1 0 21068 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_235
timestamp -25199
transform 1 0 22724 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_238
timestamp -25199
transform 1 0 23000 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_255
timestamp -25199
transform 1 0 24564 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_294
timestamp -25199
transform 1 0 28152 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_317
timestamp -25199
transform 1 0 30268 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_334
timestamp -25199
transform 1 0 31832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_357
timestamp -25199
transform 1 0 33948 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_365
timestamp -25199
transform 1 0 34684 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1636943256
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_15
timestamp -25199
transform 1 0 2484 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_23
timestamp -25199
transform 1 0 3220 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_31
timestamp -25199
transform 1 0 3956 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_41
timestamp 1636943256
transform 1 0 4876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp -25199
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_73
timestamp -25199
transform 1 0 7820 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_96
timestamp -25199
transform 1 0 9936 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp -25199
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp -25199
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_127
timestamp -25199
transform 1 0 12788 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp -25199
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_180
timestamp -25199
transform 1 0 17664 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_188
timestamp -25199
transform 1 0 18400 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_216
timestamp -25199
transform 1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_240
timestamp -25199
transform 1 0 23184 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp -25199
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_289
timestamp -25199
transform 1 0 27692 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_317
timestamp -25199
transform 1 0 30268 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp -25199
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_339
timestamp -25199
transform 1 0 32292 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_360
timestamp -25199
transform 1 0 34224 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_368
timestamp -25199
transform 1 0 34960 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_8
timestamp 1636943256
transform 1 0 1840 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_20
timestamp -25199
transform 1 0 2944 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp -25199
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_44
timestamp -25199
transform 1 0 5152 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_62
timestamp -25199
transform 1 0 6808 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1636943256
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_97
timestamp -25199
transform 1 0 10028 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_114
timestamp -25199
transform 1 0 11592 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_153
timestamp -25199
transform 1 0 15180 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_158
timestamp -25199
transform 1 0 15640 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_178
timestamp -25199
transform 1 0 17480 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp -25199
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_197
timestamp -25199
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_202
timestamp 1636943256
transform 1 0 19688 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp -25199
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_270
timestamp -25199
transform 1 0 25944 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_291
timestamp -25199
transform 1 0 27876 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp -25199
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_347
timestamp -25199
transform 1 0 33028 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_355
timestamp -25199
transform 1 0 33764 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_365
timestamp -25199
transform 1 0 34684 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636943256
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_15
timestamp -25199
transform 1 0 2484 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_23
timestamp -25199
transform 1 0 3220 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_42
timestamp 1636943256
transform 1 0 4968 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp -25199
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_81
timestamp -25199
transform 1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp -25199
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp -25199
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_129
timestamp -25199
transform 1 0 12972 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_137
timestamp -25199
transform 1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp -25199
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_177
timestamp -25199
transform 1 0 17388 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_197
timestamp -25199
transform 1 0 19228 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_203
timestamp -25199
transform 1 0 19780 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_215
timestamp -25199
transform 1 0 20884 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_221
timestamp -25199
transform 1 0 21436 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp -25199
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_285
timestamp -25199
transform 1 0 27324 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_293
timestamp -25199
transform 1 0 28060 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_316
timestamp 1636943256
transform 1 0 30176 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_328
timestamp -25199
transform 1 0 31280 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1636943256
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1636943256
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_361
timestamp -25199
transform 1 0 34316 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636943256
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636943256
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp -25199
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636943256
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636943256
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1636943256
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1636943256
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp -25199
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp -25199
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp -25199
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp -25199
transform 1 0 9660 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_104
timestamp -25199
transform 1 0 10672 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_115
timestamp -25199
transform 1 0 11684 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_126
timestamp 1636943256
transform 1 0 12696 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp -25199
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_159
timestamp 1636943256
transform 1 0 15732 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_182
timestamp -25199
transform 1 0 17848 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_186
timestamp -25199
transform 1 0 18216 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp -25199
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_197
timestamp -25199
transform 1 0 19228 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_214
timestamp 1636943256
transform 1 0 20792 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_226
timestamp -25199
transform 1 0 21896 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_253
timestamp -25199
transform 1 0 24380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_257
timestamp -25199
transform 1 0 24748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_274
timestamp -25199
transform 1 0 26312 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_293
timestamp -25199
transform 1 0 28060 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp -25199
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_312
timestamp -25199
transform 1 0 29808 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_319
timestamp -25199
transform 1 0 30452 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_332
timestamp 1636943256
transform 1 0 31648 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_365
timestamp -25199
transform 1 0 34684 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636943256
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1636943256
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_27
timestamp -25199
transform 1 0 3588 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_38
timestamp 1636943256
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp -25199
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636943256
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_69
timestamp -25199
transform 1 0 7452 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_90
timestamp -25199
transform 1 0 9384 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_96
timestamp -25199
transform 1 0 9936 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp -25199
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1636943256
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp -25199
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_129
timestamp -25199
transform 1 0 12972 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_154
timestamp 1636943256
transform 1 0 15272 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp -25199
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_185
timestamp -25199
transform 1 0 18124 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_193
timestamp -25199
transform 1 0 18860 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_197
timestamp -25199
transform 1 0 19228 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_207
timestamp 1636943256
transform 1 0 20148 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_219
timestamp -25199
transform 1 0 21252 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_229
timestamp -25199
transform 1 0 22172 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_252
timestamp -25199
transform 1 0 24288 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp -25199
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_281
timestamp -25199
transform 1 0 26956 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_285
timestamp -25199
transform 1 0 27324 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_289
timestamp -25199
transform 1 0 27692 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_297
timestamp -25199
transform 1 0 28428 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_309
timestamp -25199
transform 1 0 29532 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_337
timestamp -25199
transform 1 0 32108 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_358
timestamp -25199
transform 1 0 34040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_362
timestamp -25199
transform 1 0 34408 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_10
timestamp 1636943256
transform 1 0 2024 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_22
timestamp -25199
transform 1 0 3128 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_47
timestamp -25199
transform 1 0 5428 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp -25199
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_110
timestamp -25199
transform 1 0 11224 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_129
timestamp -25199
transform 1 0 12972 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp -25199
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_144
timestamp -25199
transform 1 0 14352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_147
timestamp -25199
transform 1 0 14628 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_166
timestamp -25199
transform 1 0 16376 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_185
timestamp -25199
transform 1 0 18124 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp -25199
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_227
timestamp -25199
transform 1 0 21988 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp -25199
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_253
timestamp -25199
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_261
timestamp -25199
transform 1 0 25116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_267
timestamp -25199
transform 1 0 25668 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_276
timestamp -25199
transform 1 0 26496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp -25199
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_321
timestamp -25199
transform 1 0 30636 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_349
timestamp -25199
transform 1 0 33212 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp -25199
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_365
timestamp -25199
transform 1 0 34684 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp -25199
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp -25199
transform 1 0 2116 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_45
timestamp -25199
transform 1 0 5244 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp -25199
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_65
timestamp -25199
transform 1 0 7084 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_95
timestamp -25199
transform 1 0 9844 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_115
timestamp -25199
transform 1 0 11684 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_135
timestamp -25199
transform 1 0 13524 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_145
timestamp -25199
transform 1 0 14444 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_153
timestamp -25199
transform 1 0 15180 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp -25199
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp -25199
transform 1 0 17756 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp -25199
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_241
timestamp -25199
transform 1 0 23276 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_254
timestamp -25199
transform 1 0 24472 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp -25199
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_281
timestamp -25199
transform 1 0 26956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_288
timestamp -25199
transform 1 0 27600 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_297
timestamp -25199
transform 1 0 28428 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_311
timestamp -25199
transform 1 0 29716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp -25199
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp -25199
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_343
timestamp 1636943256
transform 1 0 32660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_355
timestamp -25199
transform 1 0 33764 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_365
timestamp -25199
transform 1 0 34684 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636943256
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_15
timestamp -25199
transform 1 0 2484 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp -25199
transform 1 0 3220 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_32
timestamp -25199
transform 1 0 4048 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_58
timestamp -25199
transform 1 0 6440 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_64
timestamp -25199
transform 1 0 6992 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_67
timestamp 1636943256
transform 1 0 7268 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_79
timestamp -25199
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp -25199
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1636943256
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_97
timestamp -25199
transform 1 0 10028 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_104
timestamp 1636943256
transform 1 0 10672 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_116
timestamp 1636943256
transform 1 0 11776 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_130
timestamp -25199
transform 1 0 13064 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp -25199
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_152
timestamp -25199
transform 1 0 15088 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_155
timestamp -25199
transform 1 0 15364 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_175
timestamp -25199
transform 1 0 17204 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_179
timestamp -25199
transform 1 0 17572 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_242
timestamp -25199
transform 1 0 23368 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp -25199
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_259
timestamp 1636943256
transform 1 0 24932 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_271
timestamp 1636943256
transform 1 0 26036 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_283
timestamp -25199
transform 1 0 27140 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_287
timestamp -25199
transform 1 0 27508 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_290
timestamp 1636943256
transform 1 0 27784 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_302
timestamp -25199
transform 1 0 28888 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_309
timestamp -25199
transform 1 0 29532 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_317
timestamp -25199
transform 1 0 30268 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_323
timestamp -25199
transform 1 0 30820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_331
timestamp -25199
transform 1 0 31556 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_339
timestamp 1636943256
transform 1 0 32292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_351
timestamp -25199
transform 1 0 33396 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp -25199
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_8
timestamp 1636943256
transform 1 0 1840 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_20
timestamp 1636943256
transform 1 0 2944 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_32
timestamp 1636943256
transform 1 0 4048 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_44
timestamp 1636943256
transform 1 0 5152 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1636943256
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_69
timestamp -25199
transform 1 0 7452 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_75
timestamp -25199
transform 1 0 8004 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_92
timestamp -25199
transform 1 0 9568 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp -25199
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_134
timestamp -25199
transform 1 0 13432 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_151
timestamp 1636943256
transform 1 0 14996 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp -25199
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp -25199
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_180
timestamp 1636943256
transform 1 0 17664 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_192
timestamp 1636943256
transform 1 0 18768 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp -25199
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp -25199
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_239
timestamp -25199
transform 1 0 23092 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_247
timestamp -25199
transform 1 0 23828 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_257
timestamp -25199
transform 1 0 24748 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_270
timestamp -25199
transform 1 0 25944 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_274
timestamp -25199
transform 1 0 26312 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp -25199
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_299
timestamp -25199
transform 1 0 28612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_305
timestamp -25199
transform 1 0 29164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp -25199
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp -25199
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1636943256
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636943256
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636943256
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp -25199
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_29
timestamp -25199
transform 1 0 3772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_44
timestamp -25199
transform 1 0 5152 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_50
timestamp -25199
transform 1 0 5704 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_62
timestamp -25199
transform 1 0 6808 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp -25199
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp -25199
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_110
timestamp -25199
transform 1 0 11224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_130
timestamp -25199
transform 1 0 13064 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp -25199
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp -25199
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_169
timestamp -25199
transform 1 0 16652 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_177
timestamp -25199
transform 1 0 17388 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_180
timestamp -25199
transform 1 0 17664 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_184
timestamp -25199
transform 1 0 18032 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp -25199
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_212
timestamp 1636943256
transform 1 0 20608 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_224
timestamp -25199
transform 1 0 21712 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_241
timestamp -25199
transform 1 0 23276 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_303
timestamp -25199
transform 1 0 28980 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_309
timestamp -25199
transform 1 0 29532 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_334
timestamp 1636943256
transform 1 0 31832 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_346
timestamp 1636943256
transform 1 0 32936 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_365
timestamp -25199
transform 1 0 34684 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp -25199
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_7
timestamp -25199
transform 1 0 1748 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_57
timestamp -25199
transform 1 0 6348 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_85
timestamp -25199
transform 1 0 8924 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_93
timestamp -25199
transform 1 0 9660 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_96
timestamp -25199
transform 1 0 9936 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_107
timestamp -25199
transform 1 0 10948 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp -25199
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1636943256
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_125
timestamp -25199
transform 1 0 12604 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_138
timestamp -25199
transform 1 0 13800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_142
timestamp -25199
transform 1 0 14168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_165
timestamp -25199
transform 1 0 16284 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_178
timestamp -25199
transform 1 0 17480 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp -25199
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp -25199
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp -25199
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_285
timestamp -25199
transform 1 0 27324 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_309
timestamp -25199
transform 1 0 29532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_312
timestamp -25199
transform 1 0 29808 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_326
timestamp -25199
transform 1 0 31096 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_334
timestamp -25199
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1636943256
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1636943256
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_361
timestamp -25199
transform 1 0 34316 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636943256
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636943256
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp -25199
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_47
timestamp 1636943256
transform 1 0 5428 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_59
timestamp 1636943256
transform 1 0 6532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_71
timestamp 1636943256
transform 1 0 7636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp -25199
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_85
timestamp -25199
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_93
timestamp -25199
transform 1 0 9660 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_97
timestamp -25199
transform 1 0 10028 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_112
timestamp -25199
transform 1 0 11408 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp -25199
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp -25199
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_162
timestamp -25199
transform 1 0 16008 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_179
timestamp -25199
transform 1 0 17572 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp -25199
transform 1 0 20700 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_241
timestamp -25199
transform 1 0 23276 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_245
timestamp -25199
transform 1 0 23644 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_253
timestamp -25199
transform 1 0 24380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_278
timestamp -25199
transform 1 0 26680 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_331
timestamp 1636943256
transform 1 0 31556 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_343
timestamp -25199
transform 1 0 32660 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_365
timestamp -25199
transform 1 0 34684 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_11
timestamp 1636943256
transform 1 0 2116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_23
timestamp -25199
transform 1 0 3220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp -25199
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp -25199
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1636943256
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_69
timestamp -25199
transform 1 0 7452 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_73
timestamp -25199
transform 1 0 7820 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp -25199
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1636943256
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_125
timestamp -25199
transform 1 0 12604 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_146
timestamp -25199
transform 1 0 14536 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_182
timestamp -25199
transform 1 0 17848 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_192
timestamp -25199
transform 1 0 18768 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_197
timestamp -25199
transform 1 0 19228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp -25199
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp -25199
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_230
timestamp 1636943256
transform 1 0 22264 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_242
timestamp -25199
transform 1 0 23368 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp -25199
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp -25199
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_281
timestamp -25199
transform 1 0 26956 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_284
timestamp -25199
transform 1 0 27232 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_331
timestamp -25199
transform 1 0 31556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp -25199
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1636943256
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_349
timestamp -25199
transform 1 0 33212 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636943256
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636943256
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp -25199
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp -25199
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_46
timestamp -25199
transform 1 0 5336 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_63
timestamp -25199
transform 1 0 6900 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp -25199
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_107
timestamp -25199
transform 1 0 10948 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_119
timestamp -25199
transform 1 0 12052 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp -25199
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp -25199
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_167
timestamp -25199
transform 1 0 16468 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_176
timestamp -25199
transform 1 0 17296 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_182
timestamp -25199
transform 1 0 17848 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_237
timestamp -25199
transform 1 0 22908 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp -25199
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_269
timestamp -25199
transform 1 0 25852 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_273
timestamp -25199
transform 1 0 26220 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_280
timestamp -25199
transform 1 0 26864 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_292
timestamp -25199
transform 1 0 27968 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_300
timestamp -25199
transform 1 0 28704 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_320
timestamp 1636943256
transform 1 0 30544 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_332
timestamp 1636943256
transform 1 0 31648 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_344
timestamp 1636943256
transform 1 0 32752 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_356
timestamp -25199
transform 1 0 33856 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_365
timestamp -25199
transform 1 0 34684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_3
timestamp -25199
transform 1 0 1380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_11
timestamp -25199
transform 1 0 2116 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp -25199
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_59
timestamp -25199
transform 1 0 6532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_79
timestamp -25199
transform 1 0 8372 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_124
timestamp -25199
transform 1 0 12512 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_130
timestamp -25199
transform 1 0 13064 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_139
timestamp 1636943256
transform 1 0 13892 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_151
timestamp -25199
transform 1 0 14996 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp -25199
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp -25199
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_169
timestamp -25199
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_193
timestamp -25199
transform 1 0 18860 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_210
timestamp -25199
transform 1 0 20424 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_214
timestamp -25199
transform 1 0 20792 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_227
timestamp -25199
transform 1 0 21988 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_315
timestamp -25199
transform 1 0 30084 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp -25199
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1636943256
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_349
timestamp -25199
transform 1 0 33212 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_8
timestamp 1636943256
transform 1 0 1840 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp -25199
transform 1 0 2944 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_32
timestamp -25199
transform 1 0 4048 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_42
timestamp 1636943256
transform 1 0 4968 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1636943256
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp -25199
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp -25199
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_89
timestamp -25199
transform 1 0 9292 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_95
timestamp -25199
transform 1 0 9844 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_98
timestamp 1636943256
transform 1 0 10120 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp -25199
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_115
timestamp -25199
transform 1 0 11684 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_119
timestamp -25199
transform 1 0 12052 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_131
timestamp -25199
transform 1 0 13156 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp -25199
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_143
timestamp 1636943256
transform 1 0 14260 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_155
timestamp -25199
transform 1 0 15364 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1636943256
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp -25199
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp -25199
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1636943256
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_221
timestamp -25199
transform 1 0 21436 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_227
timestamp -25199
transform 1 0 21988 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp -25199
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_257
timestamp -25199
transform 1 0 24748 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_267
timestamp -25199
transform 1 0 25668 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp -25199
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_316
timestamp -25199
transform 1 0 30176 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_334
timestamp -25199
transform 1 0 31832 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_342
timestamp -25199
transform 1 0 32568 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_365
timestamp -25199
transform 1 0 34684 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636943256
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_15
timestamp -25199
transform 1 0 2484 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_35
timestamp -25199
transform 1 0 4324 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_46
timestamp -25199
transform 1 0 5336 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp -25199
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_66
timestamp 1636943256
transform 1 0 7176 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_94
timestamp -25199
transform 1 0 9752 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_109
timestamp -25199
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_113
timestamp -25199
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp -25199
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_183
timestamp 1636943256
transform 1 0 17940 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_195
timestamp -25199
transform 1 0 19044 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_201
timestamp -25199
transform 1 0 19596 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_211
timestamp 1636943256
transform 1 0 20516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp -25199
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_238
timestamp -25199
transform 1 0 23000 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_270
timestamp -25199
transform 1 0 25944 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_308
timestamp -25199
transform 1 0 29440 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_332
timestamp -25199
transform 1 0 31648 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1636943256
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1636943256
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_361
timestamp -25199
transform 1 0 34316 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636943256
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1636943256
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp -25199
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_29
timestamp -25199
transform 1 0 3772 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_78
timestamp -25199
transform 1 0 8280 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp -25199
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_92
timestamp -25199
transform 1 0 9568 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_109
timestamp -25199
transform 1 0 11132 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_113
timestamp -25199
transform 1 0 11500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_130
timestamp -25199
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp -25199
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_141
timestamp -25199
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_163
timestamp -25199
transform 1 0 16100 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_177
timestamp -25199
transform 1 0 17388 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_197
timestamp -25199
transform 1 0 19228 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_214
timestamp -25199
transform 1 0 20792 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp -25199
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_253
timestamp -25199
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_271
timestamp -25199
transform 1 0 26036 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_290
timestamp -25199
transform 1 0 27784 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_330
timestamp 1636943256
transform 1 0 31464 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_342
timestamp 1636943256
transform 1 0 32568 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_354
timestamp -25199
transform 1 0 33672 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_362
timestamp -25199
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_365
timestamp -25199
transform 1 0 34684 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636943256
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636943256
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_38
timestamp -25199
transform 1 0 4600 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp -25199
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp -25199
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_69
timestamp -25199
transform 1 0 7452 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_95
timestamp -25199
transform 1 0 9844 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp -25199
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_113
timestamp -25199
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_121
timestamp -25199
transform 1 0 12236 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_135
timestamp -25199
transform 1 0 13524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp -25199
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_185
timestamp -25199
transform 1 0 18124 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_198
timestamp -25199
transform 1 0 19320 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_211
timestamp 1636943256
transform 1 0 20516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp -25199
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_225
timestamp -25199
transform 1 0 21804 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_234
timestamp 1636943256
transform 1 0 22632 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_246
timestamp -25199
transform 1 0 23736 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_271
timestamp -25199
transform 1 0 26036 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp -25199
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1636943256
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1636943256
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_305
timestamp -25199
transform 1 0 29164 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_311
timestamp -25199
transform 1 0 29716 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_316
timestamp -25199
transform 1 0 30176 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_326
timestamp -25199
transform 1 0 31096 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_334
timestamp -25199
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1636943256
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_11
timestamp 1636943256
transform 1 0 2116 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_23
timestamp -25199
transform 1 0 3220 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp -25199
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_31
timestamp 1636943256
transform 1 0 3956 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_43
timestamp -25199
transform 1 0 5060 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_51
timestamp 1636943256
transform 1 0 5796 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_63
timestamp -25199
transform 1 0 6900 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_71
timestamp 1636943256
transform 1 0 7636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp -25199
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_87
timestamp -25199
transform 1 0 9108 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_95
timestamp 1636943256
transform 1 0 9844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_107
timestamp -25199
transform 1 0 10948 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_116
timestamp -25199
transform 1 0 11776 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp -25199
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_141
timestamp -25199
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_149
timestamp -25199
transform 1 0 14812 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_163
timestamp -25199
transform 1 0 16100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_169
timestamp -25199
transform 1 0 16652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_187
timestamp -25199
transform 1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp -25199
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1636943256
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1636943256
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_232
timestamp -25199
transform 1 0 22448 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp -25199
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp -25199
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp -25199
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_276
timestamp -25199
transform 1 0 26496 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_286
timestamp 1636943256
transform 1 0 27416 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_298
timestamp -25199
transform 1 0 28520 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_311
timestamp -25199
transform 1 0 29716 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_331
timestamp 1636943256
transform 1 0 31556 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_343
timestamp 1636943256
transform 1 0 32660 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_361
timestamp -25199
transform 1 0 34316 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_365
timestamp -25199
transform 1 0 34684 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1636943256
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_15
timestamp -25199
transform 1 0 2484 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_43
timestamp 1636943256
transform 1 0 5060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp -25199
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_57
timestamp -25199
transform 1 0 6348 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_61
timestamp -25199
transform 1 0 6716 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_71
timestamp -25199
transform 1 0 7636 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_90
timestamp -25199
transform 1 0 9384 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp -25199
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_120
timestamp -25199
transform 1 0 12144 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp -25199
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_169
timestamp -25199
transform 1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_195
timestamp -25199
transform 1 0 19044 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_203
timestamp -25199
transform 1 0 19780 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_218
timestamp -25199
transform 1 0 21160 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_229
timestamp -25199
transform 1 0 22172 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_246
timestamp -25199
transform 1 0 23736 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_267
timestamp -25199
transform 1 0 25668 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_273
timestamp -25199
transform 1 0 26220 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_297
timestamp -25199
transform 1 0 28428 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_314
timestamp -25199
transform 1 0 29992 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_322
timestamp -25199
transform 1 0 30728 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1636943256
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_349
timestamp -25199
transform 1 0 33212 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_361
timestamp -25199
transform 1 0 34316 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_3
timestamp -25199
transform 1 0 1380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_11
timestamp -25199
transform 1 0 2116 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_29
timestamp -25199
transform 1 0 3772 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_71
timestamp -25199
transform 1 0 7636 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_108
timestamp -25199
transform 1 0 11040 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_121
timestamp -25199
transform 1 0 12236 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_128
timestamp -25199
transform 1 0 12880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_143
timestamp -25199
transform 1 0 14260 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_169
timestamp -25199
transform 1 0 16652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_179
timestamp -25199
transform 1 0 17572 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_213
timestamp -25199
transform 1 0 20700 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_253
timestamp -25199
transform 1 0 24380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_261
timestamp -25199
transform 1 0 25116 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_275
timestamp -25199
transform 1 0 26404 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_294
timestamp -25199
transform 1 0 28152 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_318
timestamp -25199
transform 1 0 30360 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_333
timestamp -25199
transform 1 0 31740 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_341
timestamp -25199
transform 1 0 32476 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_365
timestamp -25199
transform 1 0 34684 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_8
timestamp -25199
transform 1 0 1840 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_16
timestamp -25199
transform 1 0 2576 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_45
timestamp -25199
transform 1 0 5244 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_77
timestamp -25199
transform 1 0 8188 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_83
timestamp -25199
transform 1 0 8740 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_86
timestamp 1636943256
transform 1 0 9016 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_98
timestamp 1636943256
transform 1 0 10120 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp -25199
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_129
timestamp 1636943256
transform 1 0 12972 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_141
timestamp -25199
transform 1 0 14076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_155
timestamp -25199
transform 1 0 15364 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp -25199
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_187
timestamp 1636943256
transform 1 0 18308 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_199
timestamp -25199
transform 1 0 19412 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_213
timestamp -25199
transform 1 0 20700 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_240
timestamp 1636943256
transform 1 0 23184 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_252
timestamp -25199
transform 1 0 24288 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_301
timestamp -25199
transform 1 0 28796 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_309
timestamp 1636943256
transform 1 0 29532 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_321
timestamp 1636943256
transform 1 0 30636 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_333
timestamp -25199
transform 1 0 31740 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1636943256
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1636943256
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_361
timestamp -25199
transform 1 0 34316 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636943256
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_15
timestamp -25199
transform 1 0 2484 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_23
timestamp -25199
transform 1 0 3220 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_26
timestamp -25199
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1636943256
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_41
timestamp -25199
transform 1 0 4876 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_51
timestamp -25199
transform 1 0 5796 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_55
timestamp -25199
transform 1 0 6164 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_60
timestamp 1636943256
transform 1 0 6624 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_72
timestamp 1636943256
transform 1 0 7728 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1636943256
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1636943256
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1636943256
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1636943256
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp -25199
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp -25199
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_141
timestamp -25199
transform 1 0 14076 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_154
timestamp 1636943256
transform 1 0 15272 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_166
timestamp -25199
transform 1 0 16376 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_174
timestamp -25199
transform 1 0 17112 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_178
timestamp 1636943256
transform 1 0 17480 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_190
timestamp -25199
transform 1 0 18584 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_48_197
timestamp -25199
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_205
timestamp -25199
transform 1 0 19964 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_217
timestamp 1636943256
transform 1 0 21068 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_229
timestamp -25199
transform 1 0 22172 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp -25199
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1636943256
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1636943256
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_277
timestamp -25199
transform 1 0 26588 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_299
timestamp -25199
transform 1 0 28612 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_305
timestamp -25199
transform 1 0 29164 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_320
timestamp 1636943256
transform 1 0 30544 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_332
timestamp 1636943256
transform 1 0 31648 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_344
timestamp 1636943256
transform 1 0 32752 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_356
timestamp -25199
transform 1 0 33856 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_365
timestamp -25199
transform 1 0 34684 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1636943256
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_15
timestamp -25199
transform 1 0 2484 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_32
timestamp -25199
transform 1 0 4048 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_43
timestamp -25199
transform 1 0 5060 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_66
timestamp -25199
transform 1 0 7176 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_95
timestamp -25199
transform 1 0 9844 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_109
timestamp -25199
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1636943256
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_125
timestamp -25199
transform 1 0 12604 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_156
timestamp -25199
transform 1 0 15456 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_171
timestamp -25199
transform 1 0 16836 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_188
timestamp 1636943256
transform 1 0 18400 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_200
timestamp -25199
transform 1 0 19504 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_218
timestamp -25199
transform 1 0 21160 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_250
timestamp -25199
transform 1 0 24104 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_265
timestamp 1636943256
transform 1 0 25484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_277
timestamp -25199
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_292
timestamp -25199
transform 1 0 27968 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_307
timestamp -25199
transform 1 0 29348 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_324
timestamp 1636943256
transform 1 0 30912 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1636943256
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1636943256
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_361
timestamp -25199
transform 1 0 34316 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_3
timestamp -25199
transform 1 0 1380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_11
timestamp -25199
transform 1 0 2116 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_85
timestamp -25199
transform 1 0 8924 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_90
timestamp -25199
transform 1 0 9384 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_108
timestamp -25199
transform 1 0 11040 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp -25199
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp -25199
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_145
timestamp -25199
transform 1 0 14444 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_154
timestamp -25199
transform 1 0 15272 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_171
timestamp -25199
transform 1 0 16836 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_188
timestamp -25199
transform 1 0 18400 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_193
timestamp -25199
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_222
timestamp -25199
transform 1 0 21528 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_226
timestamp -25199
transform 1 0 21896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_236
timestamp -25199
transform 1 0 22816 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_246
timestamp -25199
transform 1 0 23736 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_269
timestamp -25199
transform 1 0 25852 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_287
timestamp -25199
transform 1 0 27508 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_291
timestamp -25199
transform 1 0 27876 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_322
timestamp 1636943256
transform 1 0 30728 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_334
timestamp -25199
transform 1 0 31832 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_342
timestamp -25199
transform 1 0 32568 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_365
timestamp -25199
transform 1 0 34684 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_8
timestamp 1636943256
transform 1 0 1840 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_20
timestamp 1636943256
transform 1 0 2944 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_32
timestamp -25199
transform 1 0 4048 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_45
timestamp -25199
transform 1 0 5244 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_53
timestamp -25199
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1636943256
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1636943256
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_81
timestamp -25199
transform 1 0 8556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_96
timestamp -25199
transform 1 0 9936 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp -25199
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1636943256
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_125
timestamp -25199
transform 1 0 12604 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_143
timestamp -25199
transform 1 0 14260 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_155
timestamp -25199
transform 1 0 15364 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1636943256
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_181
timestamp -25199
transform 1 0 17756 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_191
timestamp -25199
transform 1 0 18676 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_203
timestamp -25199
transform 1 0 19780 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_211
timestamp -25199
transform 1 0 20516 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp -25199
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_227
timestamp -25199
transform 1 0 21988 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_235
timestamp -25199
transform 1 0 22724 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_247
timestamp 1636943256
transform 1 0 23828 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1636943256
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_273
timestamp -25199
transform 1 0 26220 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_277
timestamp -25199
transform 1 0 26588 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_299
timestamp -25199
transform 1 0 28612 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_311
timestamp 1636943256
transform 1 0 29716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_323
timestamp 1636943256
transform 1 0 30820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp -25199
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1636943256
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_349
timestamp -25199
transform 1 0 33212 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1636943256
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1636943256
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp -25199
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp -25199
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_50
timestamp -25199
transform 1 0 5704 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_67
timestamp 1636943256
transform 1 0 7268 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_79
timestamp -25199
transform 1 0 8372 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp -25199
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1636943256
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1636943256
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1636943256
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp -25199
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_162
timestamp 1636943256
transform 1 0 16008 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_174
timestamp -25199
transform 1 0 17112 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_180
timestamp -25199
transform 1 0 17664 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_188
timestamp -25199
transform 1 0 18400 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp -25199
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_208
timestamp -25199
transform 1 0 20240 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_226
timestamp -25199
transform 1 0 21896 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_246
timestamp -25199
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_274
timestamp 1636943256
transform 1 0 26312 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_286
timestamp -25199
transform 1 0 27416 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_294
timestamp -25199
transform 1 0 28152 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp -25199
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_309
timestamp -25199
transform 1 0 29532 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_317
timestamp -25199
transform 1 0 30268 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_337
timestamp 1636943256
transform 1 0 32108 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_349
timestamp -25199
transform 1 0 33212 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_357
timestamp -25199
transform 1 0 33948 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_365
timestamp -25199
transform 1 0 34684 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_5
timestamp -25199
transform 1 0 1564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_13
timestamp -25199
transform 1 0 2300 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp -25199
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp -25199
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_73
timestamp -25199
transform 1 0 7820 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_101
timestamp -25199
transform 1 0 10396 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_105
timestamp -25199
transform 1 0 10764 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_127
timestamp 1636943256
transform 1 0 12788 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_139
timestamp 1636943256
transform 1 0 13892 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_151
timestamp 1636943256
transform 1 0 14996 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_163
timestamp -25199
transform 1 0 16100 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp -25199
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_178
timestamp -25199
transform 1 0 17480 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_206
timestamp -25199
transform 1 0 20056 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_210
timestamp -25199
transform 1 0 20424 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp -25199
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_225
timestamp -25199
transform 1 0 21804 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_233
timestamp -25199
transform 1 0 22540 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_251
timestamp -25199
transform 1 0 24196 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_283
timestamp -25199
transform 1 0 27140 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_291
timestamp -25199
transform 1 0 27876 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_309
timestamp -25199
transform 1 0 29532 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_313
timestamp -25199
transform 1 0 29900 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_330
timestamp -25199
transform 1 0 31464 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1636943256
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_349
timestamp -25199
transform 1 0 33212 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1636943256
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp -25199
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_39
timestamp -25199
transform 1 0 4692 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_79
timestamp -25199
transform 1 0 8372 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp -25199
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_95
timestamp -25199
transform 1 0 9844 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_125
timestamp -25199
transform 1 0 12604 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp -25199
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1636943256
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_153
timestamp -25199
transform 1 0 15180 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_170
timestamp -25199
transform 1 0 16744 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_174
timestamp -25199
transform 1 0 17112 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_191
timestamp -25199
transform 1 0 18676 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp -25199
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1636943256
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1636943256
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_232
timestamp -25199
transform 1 0 22448 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_236
timestamp -25199
transform 1 0 22816 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp -25199
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1636943256
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_265
timestamp -25199
transform 1 0 25484 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_274
timestamp -25199
transform 1 0 26312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_305
timestamp -25199
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_327
timestamp 1636943256
transform 1 0 31188 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_339
timestamp -25199
transform 1 0 32292 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_343
timestamp -25199
transform 1 0 32660 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_365
timestamp -25199
transform 1 0 34684 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1636943256
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_15
timestamp -25199
transform 1 0 2484 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_23
timestamp -25199
transform 1 0 3220 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_41
timestamp 1636943256
transform 1 0 4876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp -25199
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_60
timestamp 1636943256
transform 1 0 6624 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_97
timestamp -25199
transform 1 0 10028 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp -25199
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_113
timestamp -25199
transform 1 0 11500 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_121
timestamp -25199
transform 1 0 12236 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_138
timestamp -25199
transform 1 0 13800 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_144
timestamp -25199
transform 1 0 14352 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_156
timestamp 1636943256
transform 1 0 15456 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_180
timestamp 1636943256
transform 1 0 17664 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_192
timestamp -25199
transform 1 0 18768 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_198
timestamp -25199
transform 1 0 19320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_210
timestamp -25199
transform 1 0 20424 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp -25199
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_229
timestamp -25199
transform 1 0 22172 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_249
timestamp -25199
transform 1 0 24012 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_262
timestamp 1636943256
transform 1 0 25208 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_274
timestamp -25199
transform 1 0 26312 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_281
timestamp -25199
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_289
timestamp -25199
transform 1 0 27692 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_323
timestamp 1636943256
transform 1 0 30820 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp -25199
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1636943256
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1636943256
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_361
timestamp -25199
transform 1 0 34316 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636943256
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1636943256
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp -25199
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1636943256
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_41
timestamp -25199
transform 1 0 4876 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_56_65
timestamp -25199
transform 1 0 7084 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_80
timestamp -25199
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_85
timestamp -25199
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_95
timestamp -25199
transform 1 0 9844 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_104
timestamp -25199
transform 1 0 10672 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_112
timestamp -25199
transform 1 0 11408 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_137
timestamp -25199
transform 1 0 13708 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_157
timestamp -25199
transform 1 0 15548 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_188
timestamp -25199
transform 1 0 18400 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_213
timestamp -25199
transform 1 0 20700 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_239
timestamp -25199
transform 1 0 23092 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_243
timestamp -25199
transform 1 0 23460 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_247
timestamp -25199
transform 1 0 23828 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp -25199
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_287
timestamp 1636943256
transform 1 0 27508 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_303
timestamp -25199
transform 1 0 28980 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp -25199
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_325
timestamp 1636943256
transform 1 0 31004 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_337
timestamp -25199
transform 1 0 32108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_365
timestamp -25199
transform 1 0 34684 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1636943256
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1636943256
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1636943256
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_39
timestamp -25199
transform 1 0 4692 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_79
timestamp -25199
transform 1 0 8372 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_83
timestamp -25199
transform 1 0 8740 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_104
timestamp -25199
transform 1 0 10672 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_129
timestamp 1636943256
transform 1 0 12972 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_141
timestamp -25199
transform 1 0 14076 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_149
timestamp -25199
transform 1 0 14812 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_185
timestamp -25199
transform 1 0 18124 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_201
timestamp -25199
transform 1 0 19596 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_209
timestamp -25199
transform 1 0 20332 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp -25199
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_227
timestamp -25199
transform 1 0 21988 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_241
timestamp 1636943256
transform 1 0 23276 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_253
timestamp -25199
transform 1 0 24380 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_261
timestamp -25199
transform 1 0 25116 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_290
timestamp -25199
transform 1 0 27784 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_294
timestamp -25199
transform 1 0 28152 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_305
timestamp -25199
transform 1 0 29164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1636943256
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp -25199
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp -25199
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_363
timestamp -25199
transform 1 0 34500 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_8
timestamp 1636943256
transform 1 0 1840 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_20
timestamp -25199
transform 1 0 2944 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1636943256
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_41
timestamp -25199
transform 1 0 4876 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_45
timestamp -25199
transform 1 0 5244 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_74
timestamp -25199
transform 1 0 7912 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp -25199
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_101
timestamp -25199
transform 1 0 10396 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_114
timestamp 1636943256
transform 1 0 11592 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_126
timestamp -25199
transform 1 0 12696 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_130
timestamp -25199
transform 1 0 13064 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_143
timestamp -25199
transform 1 0 14260 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_155
timestamp -25199
transform 1 0 15364 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_163
timestamp -25199
transform 1 0 16100 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_167
timestamp -25199
transform 1 0 16468 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_170
timestamp -25199
transform 1 0 16744 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_176
timestamp -25199
transform 1 0 17296 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1636943256
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_209
timestamp -25199
transform 1 0 20332 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_217
timestamp -25199
transform 1 0 21068 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_221
timestamp -25199
transform 1 0 21436 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_227
timestamp -25199
transform 1 0 21988 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_239
timestamp -25199
transform 1 0 23092 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp -25199
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_253
timestamp -25199
transform 1 0 24380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_261
timestamp -25199
transform 1 0 25116 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_282
timestamp -25199
transform 1 0 27048 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp -25199
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp -25199
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1636943256
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1636943256
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1636943256
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_350
timestamp -25199
transform 1 0 33304 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_365
timestamp -25199
transform 1 0 34684 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1636943256
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1636943256
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1636943256
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1636943256
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp -25199
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp -25199
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1636943256
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_69
timestamp -25199
transform 1 0 7452 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_75
timestamp -25199
transform 1 0 8004 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_87
timestamp -25199
transform 1 0 9108 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_91
timestamp -25199
transform 1 0 9476 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp -25199
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_115
timestamp -25199
transform 1 0 11684 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_150
timestamp -25199
transform 1 0 14904 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_156
timestamp -25199
transform 1 0 15456 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1636943256
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_181
timestamp -25199
transform 1 0 17756 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_204
timestamp -25199
transform 1 0 19872 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_218
timestamp -25199
transform 1 0 21160 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_252
timestamp -25199
transform 1 0 24288 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_264
timestamp 1636943256
transform 1 0 25392 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp -25199
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_281
timestamp -25199
transform 1 0 26956 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_298
timestamp 1636943256
transform 1 0 28520 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_310
timestamp 1636943256
transform 1 0 29624 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_322
timestamp 1636943256
transform 1 0 30728 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp -25199
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1636943256
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1636943256
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_361
timestamp -25199
transform 1 0 34316 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_5
timestamp 1636943256
transform 1 0 1564 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_17
timestamp -25199
transform 1 0 2668 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_25
timestamp -25199
transform 1 0 3404 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1636943256
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1636943256
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1636943256
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_65
timestamp -25199
transform 1 0 7084 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_85
timestamp -25199
transform 1 0 8924 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_107
timestamp -25199
transform 1 0 10948 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_124
timestamp 1636943256
transform 1 0 12512 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp -25199
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_168
timestamp 1636943256
transform 1 0 16560 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_197
timestamp -25199
transform 1 0 19228 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_217
timestamp 1636943256
transform 1 0 21068 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp -25199
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp -25199
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp -25199
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp -25199
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1636943256
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1636943256
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1636943256
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1636943256
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp -25199
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp -25199
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_365
timestamp -25199
transform 1 0 34684 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_11
timestamp 1636943256
transform 1 0 2116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_23
timestamp -25199
transform 1 0 3220 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_27
timestamp -25199
transform 1 0 3588 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_29
timestamp 1636943256
transform 1 0 3772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_41
timestamp 1636943256
transform 1 0 4876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_53
timestamp -25199
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1636943256
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1636943256
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_81
timestamp -25199
transform 1 0 8556 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_85
timestamp 1636943256
transform 1 0 8924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_97
timestamp 1636943256
transform 1 0 10028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_109
timestamp -25199
transform 1 0 11132 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_124
timestamp 1636943256
transform 1 0 12512 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_136
timestamp -25199
transform 1 0 13616 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_141
timestamp 1636943256
transform 1 0 14076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_153
timestamp 1636943256
transform 1 0 15180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_165
timestamp -25199
transform 1 0 16284 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1636943256
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_181
timestamp -25199
transform 1 0 17756 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_208
timestamp 1636943256
transform 1 0 20240 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp -25199
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1636943256
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1636943256
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_249
timestamp -25199
transform 1 0 24012 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_253
timestamp -25199
transform 1 0 24380 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_261
timestamp -25199
transform 1 0 25116 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_274
timestamp -25199
transform 1 0 26312 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_281
timestamp -25199
transform 1 0 26956 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_296
timestamp 1636943256
transform 1 0 28336 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_309
timestamp 1636943256
transform 1 0 29532 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_321
timestamp 1636943256
transform 1 0 30636 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_333
timestamp -25199
transform 1 0 31740 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1636943256
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_349
timestamp -25199
transform 1 0 33212 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_357
timestamp -25199
transform 1 0 33948 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_365
timestamp -25199
transform 1 0 34684 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp -25199
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2
timestamp -25199
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp -25199
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp -25199
transform -1 0 1656 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp -25199
transform -1 0 1656 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp -25199
transform 1 0 1380 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp -25199
transform -1 0 1656 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp -25199
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp -25199
transform -1 0 1932 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp -25199
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp -25199
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp -25199
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp -25199
transform -1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp -25199
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp -25199
transform -1 0 1656 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp -25199
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp -25199
transform -1 0 1656 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp -25199
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp -25199
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output20
timestamp -25199
transform 1 0 34500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output21
timestamp -25199
transform 1 0 34040 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output22
timestamp -25199
transform -1 0 34592 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output23
timestamp -25199
transform 1 0 34500 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output24
timestamp -25199
transform 1 0 34500 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output25
timestamp -25199
transform 1 0 34040 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output26
timestamp -25199
transform 1 0 34500 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output27
timestamp -25199
transform 1 0 34040 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output28
timestamp -25199
transform -1 0 34592 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output29
timestamp -25199
transform 1 0 34500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output30
timestamp -25199
transform 1 0 34500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output31
timestamp -25199
transform 1 0 34500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output32
timestamp -25199
transform -1 0 34592 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output33
timestamp -25199
transform 1 0 34040 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output34
timestamp -25199
transform 1 0 34500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output35
timestamp -25199
transform -1 0 34592 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output36
timestamp -25199
transform 1 0 34500 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output37
timestamp -25199
transform 1 0 34500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_62
timestamp -25199
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -25199
transform -1 0 35328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_63
timestamp -25199
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -25199
transform -1 0 35328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_64
timestamp -25199
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -25199
transform -1 0 35328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_65
timestamp -25199
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -25199
transform -1 0 35328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_66
timestamp -25199
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -25199
transform -1 0 35328 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_67
timestamp -25199
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -25199
transform -1 0 35328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_68
timestamp -25199
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -25199
transform -1 0 35328 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_69
timestamp -25199
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -25199
transform -1 0 35328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_70
timestamp -25199
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -25199
transform -1 0 35328 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_71
timestamp -25199
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -25199
transform -1 0 35328 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_72
timestamp -25199
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -25199
transform -1 0 35328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_73
timestamp -25199
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -25199
transform -1 0 35328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_74
timestamp -25199
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -25199
transform -1 0 35328 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_75
timestamp -25199
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -25199
transform -1 0 35328 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_76
timestamp -25199
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -25199
transform -1 0 35328 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_77
timestamp -25199
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -25199
transform -1 0 35328 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_78
timestamp -25199
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -25199
transform -1 0 35328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_79
timestamp -25199
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -25199
transform -1 0 35328 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_80
timestamp -25199
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -25199
transform -1 0 35328 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_81
timestamp -25199
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -25199
transform -1 0 35328 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_82
timestamp -25199
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -25199
transform -1 0 35328 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_83
timestamp -25199
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -25199
transform -1 0 35328 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_84
timestamp -25199
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -25199
transform -1 0 35328 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_85
timestamp -25199
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -25199
transform -1 0 35328 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_86
timestamp -25199
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -25199
transform -1 0 35328 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_87
timestamp -25199
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp -25199
transform -1 0 35328 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_88
timestamp -25199
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp -25199
transform -1 0 35328 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_89
timestamp -25199
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp -25199
transform -1 0 35328 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_90
timestamp -25199
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp -25199
transform -1 0 35328 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_91
timestamp -25199
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp -25199
transform -1 0 35328 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_92
timestamp -25199
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp -25199
transform -1 0 35328 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_93
timestamp -25199
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp -25199
transform -1 0 35328 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_94
timestamp -25199
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp -25199
transform -1 0 35328 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_95
timestamp -25199
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp -25199
transform -1 0 35328 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_96
timestamp -25199
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp -25199
transform -1 0 35328 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_97
timestamp -25199
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp -25199
transform -1 0 35328 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_98
timestamp -25199
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp -25199
transform -1 0 35328 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_99
timestamp -25199
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp -25199
transform -1 0 35328 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_100
timestamp -25199
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp -25199
transform -1 0 35328 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_101
timestamp -25199
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp -25199
transform -1 0 35328 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_102
timestamp -25199
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp -25199
transform -1 0 35328 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_103
timestamp -25199
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp -25199
transform -1 0 35328 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_104
timestamp -25199
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp -25199
transform -1 0 35328 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_105
timestamp -25199
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp -25199
transform -1 0 35328 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_106
timestamp -25199
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp -25199
transform -1 0 35328 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_107
timestamp -25199
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp -25199
transform -1 0 35328 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_108
timestamp -25199
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp -25199
transform -1 0 35328 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_109
timestamp -25199
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp -25199
transform -1 0 35328 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_110
timestamp -25199
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp -25199
transform -1 0 35328 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_111
timestamp -25199
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp -25199
transform -1 0 35328 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_112
timestamp -25199
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp -25199
transform -1 0 35328 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_113
timestamp -25199
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp -25199
transform -1 0 35328 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_114
timestamp -25199
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp -25199
transform -1 0 35328 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_115
timestamp -25199
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp -25199
transform -1 0 35328 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_116
timestamp -25199
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp -25199
transform -1 0 35328 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_117
timestamp -25199
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp -25199
transform -1 0 35328 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_118
timestamp -25199
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp -25199
transform -1 0 35328 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_119
timestamp -25199
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp -25199
transform -1 0 35328 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_120
timestamp -25199
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp -25199
transform -1 0 35328 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_121
timestamp -25199
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp -25199
transform -1 0 35328 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_122
timestamp -25199
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp -25199
transform -1 0 35328 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_123
timestamp -25199
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp -25199
transform -1 0 35328 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_124
timestamp -25199
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_125
timestamp -25199
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_126
timestamp -25199
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_127
timestamp -25199
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_128
timestamp -25199
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_129
timestamp -25199
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_130
timestamp -25199
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_131
timestamp -25199
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_132
timestamp -25199
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_133
timestamp -25199
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_134
timestamp -25199
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_135
timestamp -25199
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_136
timestamp -25199
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_137
timestamp -25199
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_138
timestamp -25199
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_139
timestamp -25199
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_140
timestamp -25199
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_141
timestamp -25199
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_142
timestamp -25199
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_143
timestamp -25199
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_144
timestamp -25199
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_145
timestamp -25199
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_146
timestamp -25199
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_147
timestamp -25199
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_148
timestamp -25199
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_149
timestamp -25199
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_150
timestamp -25199
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_151
timestamp -25199
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_152
timestamp -25199
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_153
timestamp -25199
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_154
timestamp -25199
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_155
timestamp -25199
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_156
timestamp -25199
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_157
timestamp -25199
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_158
timestamp -25199
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_159
timestamp -25199
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_160
timestamp -25199
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_161
timestamp -25199
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_162
timestamp -25199
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_163
timestamp -25199
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_164
timestamp -25199
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_165
timestamp -25199
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_166
timestamp -25199
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_167
timestamp -25199
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_168
timestamp -25199
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_169
timestamp -25199
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_170
timestamp -25199
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_171
timestamp -25199
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_172
timestamp -25199
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_173
timestamp -25199
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_174
timestamp -25199
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_175
timestamp -25199
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_176
timestamp -25199
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_177
timestamp -25199
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_178
timestamp -25199
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_179
timestamp -25199
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_180
timestamp -25199
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_181
timestamp -25199
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_182
timestamp -25199
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_183
timestamp -25199
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_184
timestamp -25199
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_185
timestamp -25199
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_186
timestamp -25199
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_187
timestamp -25199
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_188
timestamp -25199
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_189
timestamp -25199
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_190
timestamp -25199
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_191
timestamp -25199
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_192
timestamp -25199
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_193
timestamp -25199
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_194
timestamp -25199
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_195
timestamp -25199
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_196
timestamp -25199
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_197
timestamp -25199
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_198
timestamp -25199
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_199
timestamp -25199
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_200
timestamp -25199
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_201
timestamp -25199
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_202
timestamp -25199
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_203
timestamp -25199
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_204
timestamp -25199
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_205
timestamp -25199
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_206
timestamp -25199
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_207
timestamp -25199
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_208
timestamp -25199
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_209
timestamp -25199
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_210
timestamp -25199
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_211
timestamp -25199
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_212
timestamp -25199
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_213
timestamp -25199
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_214
timestamp -25199
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_215
timestamp -25199
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_216
timestamp -25199
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_217
timestamp -25199
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_218
timestamp -25199
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_219
timestamp -25199
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_220
timestamp -25199
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_221
timestamp -25199
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_222
timestamp -25199
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_223
timestamp -25199
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_224
timestamp -25199
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_225
timestamp -25199
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_226
timestamp -25199
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_227
timestamp -25199
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_228
timestamp -25199
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_229
timestamp -25199
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_230
timestamp -25199
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_231
timestamp -25199
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_232
timestamp -25199
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_233
timestamp -25199
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_234
timestamp -25199
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_235
timestamp -25199
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_236
timestamp -25199
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_237
timestamp -25199
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_238
timestamp -25199
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_239
timestamp -25199
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_240
timestamp -25199
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_241
timestamp -25199
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_242
timestamp -25199
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_243
timestamp -25199
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_244
timestamp -25199
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_245
timestamp -25199
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_246
timestamp -25199
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_247
timestamp -25199
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_248
timestamp -25199
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_249
timestamp -25199
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_250
timestamp -25199
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_251
timestamp -25199
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_252
timestamp -25199
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_253
timestamp -25199
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_254
timestamp -25199
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_255
timestamp -25199
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_256
timestamp -25199
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_257
timestamp -25199
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_258
timestamp -25199
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_259
timestamp -25199
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_260
timestamp -25199
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_261
timestamp -25199
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_262
timestamp -25199
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_263
timestamp -25199
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_264
timestamp -25199
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_265
timestamp -25199
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_266
timestamp -25199
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_267
timestamp -25199
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_268
timestamp -25199
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_269
timestamp -25199
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_270
timestamp -25199
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_271
timestamp -25199
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_272
timestamp -25199
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_273
timestamp -25199
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_274
timestamp -25199
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_275
timestamp -25199
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_276
timestamp -25199
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_277
timestamp -25199
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_278
timestamp -25199
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_279
timestamp -25199
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_280
timestamp -25199
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_281
timestamp -25199
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_282
timestamp -25199
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_283
timestamp -25199
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_284
timestamp -25199
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_285
timestamp -25199
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_286
timestamp -25199
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_287
timestamp -25199
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_288
timestamp -25199
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_289
timestamp -25199
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_290
timestamp -25199
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_291
timestamp -25199
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_292
timestamp -25199
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_293
timestamp -25199
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_294
timestamp -25199
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_295
timestamp -25199
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_296
timestamp -25199
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_297
timestamp -25199
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_298
timestamp -25199
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_299
timestamp -25199
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_300
timestamp -25199
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_301
timestamp -25199
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_302
timestamp -25199
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_303
timestamp -25199
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_304
timestamp -25199
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_305
timestamp -25199
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_306
timestamp -25199
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_307
timestamp -25199
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_308
timestamp -25199
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_309
timestamp -25199
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_310
timestamp -25199
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_311
timestamp -25199
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_312
timestamp -25199
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_313
timestamp -25199
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_314
timestamp -25199
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_315
timestamp -25199
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_316
timestamp -25199
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_317
timestamp -25199
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_318
timestamp -25199
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_319
timestamp -25199
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_320
timestamp -25199
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_321
timestamp -25199
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_322
timestamp -25199
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_323
timestamp -25199
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_324
timestamp -25199
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_325
timestamp -25199
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_326
timestamp -25199
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_327
timestamp -25199
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_328
timestamp -25199
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_329
timestamp -25199
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_330
timestamp -25199
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_331
timestamp -25199
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_332
timestamp -25199
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_333
timestamp -25199
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_334
timestamp -25199
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_335
timestamp -25199
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_336
timestamp -25199
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_337
timestamp -25199
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_338
timestamp -25199
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_339
timestamp -25199
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_340
timestamp -25199
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_341
timestamp -25199
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_342
timestamp -25199
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_343
timestamp -25199
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_344
timestamp -25199
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_345
timestamp -25199
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_346
timestamp -25199
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_347
timestamp -25199
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_348
timestamp -25199
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_349
timestamp -25199
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_350
timestamp -25199
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_351
timestamp -25199
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_352
timestamp -25199
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_353
timestamp -25199
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_354
timestamp -25199
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_355
timestamp -25199
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_356
timestamp -25199
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_357
timestamp -25199
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_358
timestamp -25199
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_359
timestamp -25199
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_360
timestamp -25199
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_361
timestamp -25199
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_362
timestamp -25199
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_363
timestamp -25199
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_364
timestamp -25199
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_365
timestamp -25199
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_366
timestamp -25199
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_367
timestamp -25199
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_368
timestamp -25199
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_369
timestamp -25199
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_370
timestamp -25199
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_371
timestamp -25199
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_372
timestamp -25199
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_373
timestamp -25199
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_374
timestamp -25199
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_375
timestamp -25199
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_376
timestamp -25199
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_377
timestamp -25199
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_378
timestamp -25199
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_379
timestamp -25199
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_380
timestamp -25199
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_381
timestamp -25199
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_382
timestamp -25199
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_383
timestamp -25199
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_384
timestamp -25199
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_385
timestamp -25199
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_386
timestamp -25199
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_387
timestamp -25199
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_388
timestamp -25199
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_389
timestamp -25199
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_390
timestamp -25199
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_391
timestamp -25199
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_392
timestamp -25199
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_393
timestamp -25199
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_394
timestamp -25199
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_395
timestamp -25199
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_396
timestamp -25199
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_397
timestamp -25199
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_398
timestamp -25199
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_399
timestamp -25199
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_400
timestamp -25199
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_401
timestamp -25199
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_402
timestamp -25199
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_403
timestamp -25199
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_404
timestamp -25199
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_405
timestamp -25199
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_406
timestamp -25199
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_407
timestamp -25199
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_408
timestamp -25199
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_409
timestamp -25199
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_410
timestamp -25199
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_411
timestamp -25199
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_412
timestamp -25199
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_413
timestamp -25199
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_414
timestamp -25199
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_415
timestamp -25199
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_416
timestamp -25199
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_417
timestamp -25199
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_418
timestamp -25199
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_419
timestamp -25199
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_420
timestamp -25199
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_421
timestamp -25199
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_422
timestamp -25199
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_423
timestamp -25199
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_424
timestamp -25199
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_425
timestamp -25199
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_426
timestamp -25199
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_427
timestamp -25199
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_428
timestamp -25199
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_429
timestamp -25199
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_430
timestamp -25199
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_431
timestamp -25199
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_432
timestamp -25199
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_433
timestamp -25199
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_434
timestamp -25199
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_435
timestamp -25199
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_436
timestamp -25199
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_437
timestamp -25199
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_438
timestamp -25199
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_439
timestamp -25199
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_440
timestamp -25199
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_441
timestamp -25199
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_442
timestamp -25199
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_443
timestamp -25199
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_444
timestamp -25199
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_445
timestamp -25199
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_446
timestamp -25199
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_447
timestamp -25199
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_448
timestamp -25199
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_449
timestamp -25199
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_450
timestamp -25199
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_451
timestamp -25199
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_452
timestamp -25199
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_453
timestamp -25199
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_454
timestamp -25199
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_455
timestamp -25199
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_456
timestamp -25199
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_457
timestamp -25199
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_458
timestamp -25199
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_459
timestamp -25199
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_460
timestamp -25199
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_461
timestamp -25199
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_462
timestamp -25199
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_463
timestamp -25199
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_464
timestamp -25199
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_465
timestamp -25199
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_466
timestamp -25199
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_467
timestamp -25199
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_468
timestamp -25199
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_469
timestamp -25199
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_470
timestamp -25199
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_471
timestamp -25199
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_472
timestamp -25199
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_473
timestamp -25199
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_474
timestamp -25199
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_475
timestamp -25199
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_476
timestamp -25199
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_477
timestamp -25199
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_478
timestamp -25199
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_479
timestamp -25199
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_480
timestamp -25199
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_481
timestamp -25199
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_482
timestamp -25199
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_483
timestamp -25199
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_484
timestamp -25199
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_485
timestamp -25199
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_486
timestamp -25199
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_487
timestamp -25199
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_488
timestamp -25199
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_489
timestamp -25199
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_490
timestamp -25199
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_491
timestamp -25199
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_492
timestamp -25199
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_493
timestamp -25199
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_494
timestamp -25199
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_495
timestamp -25199
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_496
timestamp -25199
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_497
timestamp -25199
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_498
timestamp -25199
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_499
timestamp -25199
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_500
timestamp -25199
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_501
timestamp -25199
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_502
timestamp -25199
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_503
timestamp -25199
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_504
timestamp -25199
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_505
timestamp -25199
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_506
timestamp -25199
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_507
timestamp -25199
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_508
timestamp -25199
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_509
timestamp -25199
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_510
timestamp -25199
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_511
timestamp -25199
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_512
timestamp -25199
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_513
timestamp -25199
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_514
timestamp -25199
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_515
timestamp -25199
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_516
timestamp -25199
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_517
timestamp -25199
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_518
timestamp -25199
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_519
timestamp -25199
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_520
timestamp -25199
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_521
timestamp -25199
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_522
timestamp -25199
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_523
timestamp -25199
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_524
timestamp -25199
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_525
timestamp -25199
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_526
timestamp -25199
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_527
timestamp -25199
transform 1 0 3680 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_528
timestamp -25199
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_529
timestamp -25199
transform 1 0 8832 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_530
timestamp -25199
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_531
timestamp -25199
transform 1 0 13984 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_532
timestamp -25199
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_533
timestamp -25199
transform 1 0 19136 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_534
timestamp -25199
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_535
timestamp -25199
transform 1 0 24288 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_536
timestamp -25199
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_537
timestamp -25199
transform 1 0 29440 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_538
timestamp -25199
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_539
timestamp -25199
transform 1 0 34592 0 -1 35904
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 1096 800 1216 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 35673 4904 36473 5024 0 FreeSans 480 0 0 0 empty_o
port 1 nsew signal output
flabel metal3 s 35673 3000 36473 3120 0 FreeSans 480 0 0 0 full_o
port 2 nsew signal output
flabel metal3 s 35673 6808 36473 6928 0 FreeSans 480 0 0 0 rd_data_o[0]
port 3 nsew signal output
flabel metal3 s 35673 25848 36473 25968 0 FreeSans 480 0 0 0 rd_data_o[10]
port 4 nsew signal output
flabel metal3 s 35673 27752 36473 27872 0 FreeSans 480 0 0 0 rd_data_o[11]
port 5 nsew signal output
flabel metal3 s 35673 29656 36473 29776 0 FreeSans 480 0 0 0 rd_data_o[12]
port 6 nsew signal output
flabel metal3 s 35673 31560 36473 31680 0 FreeSans 480 0 0 0 rd_data_o[13]
port 7 nsew signal output
flabel metal3 s 35673 33464 36473 33584 0 FreeSans 480 0 0 0 rd_data_o[14]
port 8 nsew signal output
flabel metal3 s 35673 35368 36473 35488 0 FreeSans 480 0 0 0 rd_data_o[15]
port 9 nsew signal output
flabel metal3 s 35673 8712 36473 8832 0 FreeSans 480 0 0 0 rd_data_o[1]
port 10 nsew signal output
flabel metal3 s 35673 10616 36473 10736 0 FreeSans 480 0 0 0 rd_data_o[2]
port 11 nsew signal output
flabel metal3 s 35673 12520 36473 12640 0 FreeSans 480 0 0 0 rd_data_o[3]
port 12 nsew signal output
flabel metal3 s 35673 14424 36473 14544 0 FreeSans 480 0 0 0 rd_data_o[4]
port 13 nsew signal output
flabel metal3 s 35673 16328 36473 16448 0 FreeSans 480 0 0 0 rd_data_o[5]
port 14 nsew signal output
flabel metal3 s 35673 18232 36473 18352 0 FreeSans 480 0 0 0 rd_data_o[6]
port 15 nsew signal output
flabel metal3 s 35673 20136 36473 20256 0 FreeSans 480 0 0 0 rd_data_o[7]
port 16 nsew signal output
flabel metal3 s 35673 22040 36473 22160 0 FreeSans 480 0 0 0 rd_data_o[8]
port 17 nsew signal output
flabel metal3 s 35673 23944 36473 24064 0 FreeSans 480 0 0 0 rd_data_o[9]
port 18 nsew signal output
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 rd_en_i
port 19 nsew signal input
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 rst_n
port 20 nsew signal input
flabel metal4 s 4208 2128 4528 35952 0 FreeSans 1920 90 0 0 vccd1
port 21 nsew power bidirectional
flabel metal4 s 34928 2128 35248 35952 0 FreeSans 1920 90 0 0 vccd1
port 21 nsew power bidirectional
flabel metal4 s 4868 2128 5188 35952 0 FreeSans 1920 90 0 0 vssd1
port 22 nsew ground bidirectional
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 wr_data_i[0]
port 23 nsew signal input
flabel metal3 s 0 27752 800 27872 0 FreeSans 480 0 0 0 wr_data_i[10]
port 24 nsew signal input
flabel metal3 s 0 29656 800 29776 0 FreeSans 480 0 0 0 wr_data_i[11]
port 25 nsew signal input
flabel metal3 s 0 31560 800 31680 0 FreeSans 480 0 0 0 wr_data_i[12]
port 26 nsew signal input
flabel metal3 s 0 33464 800 33584 0 FreeSans 480 0 0 0 wr_data_i[13]
port 27 nsew signal input
flabel metal3 s 0 35368 800 35488 0 FreeSans 480 0 0 0 wr_data_i[14]
port 28 nsew signal input
flabel metal3 s 0 37272 800 37392 0 FreeSans 480 0 0 0 wr_data_i[15]
port 29 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 wr_data_i[1]
port 30 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 wr_data_i[2]
port 31 nsew signal input
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 wr_data_i[3]
port 32 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 wr_data_i[4]
port 33 nsew signal input
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 wr_data_i[5]
port 34 nsew signal input
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 wr_data_i[6]
port 35 nsew signal input
flabel metal3 s 0 22040 800 22160 0 FreeSans 480 0 0 0 wr_data_i[7]
port 36 nsew signal input
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 wr_data_i[8]
port 37 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 wr_data_i[9]
port 38 nsew signal input
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 wr_en_i
port 39 nsew signal input
rlabel metal1 18216 35360 18216 35360 0 vccd1
rlabel metal1 18216 35904 18216 35904 0 vssd1
rlabel metal2 29854 8024 29854 8024 0 _0000_
rlabel metal1 32522 8058 32522 8058 0 _0001_
rlabel metal1 27416 5610 27416 5610 0 _0002_
rlabel metal2 29854 3876 29854 3876 0 _0003_
rlabel metal2 33258 4386 33258 4386 0 _0004_
rlabel metal1 33718 6970 33718 6970 0 _0005_
rlabel metal2 33074 9180 33074 9180 0 _0006_
rlabel metal2 33534 10846 33534 10846 0 _0007_
rlabel metal1 32338 12410 32338 12410 0 _0008_
rlabel metal2 33994 14756 33994 14756 0 _0009_
rlabel metal2 32706 15572 32706 15572 0 _0010_
rlabel metal1 33442 17714 33442 17714 0 _0011_
rlabel metal2 33994 20196 33994 20196 0 _0012_
rlabel via1 33067 22202 33067 22202 0 _0013_
rlabel metal1 33534 23834 33534 23834 0 _0014_
rlabel metal2 33810 26078 33810 26078 0 _0015_
rlabel metal1 33580 27098 33580 27098 0 _0016_
rlabel metal1 33350 29682 33350 29682 0 _0017_
rlabel metal1 33902 31450 33902 31450 0 _0018_
rlabel metal1 32338 33082 32338 33082 0 _0019_
rlabel metal1 33258 32946 33258 32946 0 _0020_
rlabel metal2 33718 18462 33718 18462 0 _0021_
rlabel metal1 31280 16626 31280 16626 0 _0022_
rlabel metal2 31050 18972 31050 18972 0 _0023_
rlabel metal1 28566 16762 28566 16762 0 _0024_
rlabel metal1 22632 4250 22632 4250 0 _0025_
rlabel metal1 21482 5576 21482 5576 0 _0026_
rlabel metal1 24426 5100 24426 5100 0 _0027_
rlabel metal1 25990 6426 25990 6426 0 _0028_
rlabel metal1 17802 6970 17802 6970 0 _0029_
rlabel metal1 20741 6698 20741 6698 0 _0030_
rlabel metal1 19228 13498 19228 13498 0 _0031_
rlabel metal2 30130 12002 30130 12002 0 _0032_
rlabel via1 16794 14382 16794 14382 0 _0033_
rlabel via1 30677 15470 30677 15470 0 _0034_
rlabel metal1 16928 17850 16928 17850 0 _0035_
rlabel via1 29941 20910 29941 20910 0 _0036_
rlabel metal2 16698 21794 16698 21794 0 _0037_
rlabel metal2 30682 23970 30682 23970 0 _0038_
rlabel metal1 19637 27370 19637 27370 0 _0039_
rlabel via1 29674 26962 29674 26962 0 _0040_
rlabel metal2 30406 31518 30406 31518 0 _0041_
rlabel metal1 16146 32198 16146 32198 0 _0042_
rlabel metal1 29716 31994 29716 31994 0 _0043_
rlabel metal1 16728 33558 16728 33558 0 _0044_
rlabel metal1 17756 9146 17756 9146 0 _0045_
rlabel metal2 12374 8228 12374 8228 0 _0046_
rlabel metal1 11173 13294 11173 13294 0 _0047_
rlabel metal1 27278 8058 27278 8058 0 _0048_
rlabel metal2 11822 16694 11822 16694 0 _0049_
rlabel metal2 19918 17442 19918 17442 0 _0050_
rlabel metal1 11955 18734 11955 18734 0 _0051_
rlabel metal2 23322 18530 23322 18530 0 _0052_
rlabel metal1 10897 23766 10897 23766 0 _0053_
rlabel metal2 25530 22406 25530 22406 0 _0054_
rlabel metal1 17204 25466 17204 25466 0 _0055_
rlabel metal2 12190 24786 12190 24786 0 _0056_
rlabel metal2 27002 29410 27002 29410 0 _0057_
rlabel metal1 11035 31790 11035 31790 0 _0058_
rlabel metal2 20838 30464 20838 30464 0 _0059_
rlabel metal2 12834 30498 12834 30498 0 _0060_
rlabel metal1 16049 8466 16049 8466 0 _0061_
rlabel metal1 19775 7446 19775 7446 0 _0062_
rlabel metal2 2990 13090 2990 13090 0 _0063_
rlabel metal2 20378 12002 20378 12002 0 _0064_
rlabel metal2 4186 15266 4186 15266 0 _0065_
rlabel metal1 23041 16558 23041 16558 0 _0066_
rlabel metal1 3818 19414 3818 19414 0 _0067_
rlabel metal2 18170 21318 18170 21318 0 _0068_
rlabel metal2 3818 23222 3818 23222 0 _0069_
rlabel metal2 21482 26962 21482 26962 0 _0070_
rlabel metal1 18032 22746 18032 22746 0 _0071_
rlabel metal1 3813 27030 3813 27030 0 _0072_
rlabel metal2 22126 29342 22126 29342 0 _0073_
rlabel metal1 8827 29138 8827 29138 0 _0074_
rlabel metal1 19453 29614 19453 29614 0 _0075_
rlabel metal1 12834 29512 12834 29512 0 _0076_
rlabel metal1 16371 6766 16371 6766 0 _0077_
rlabel metal2 14214 6562 14214 6562 0 _0078_
rlabel metal1 14071 12886 14071 12886 0 _0079_
rlabel metal2 24978 10914 24978 10914 0 _0080_
rlabel metal2 12650 15266 12650 15266 0 _0081_
rlabel metal2 22218 17306 22218 17306 0 _0082_
rlabel metal2 14122 20060 14122 20060 0 _0083_
rlabel metal1 20700 19482 20700 19482 0 _0084_
rlabel metal2 12834 21794 12834 21794 0 _0085_
rlabel metal1 24789 23018 24789 23018 0 _0086_
rlabel metal1 16463 24106 16463 24106 0 _0087_
rlabel metal2 12558 26146 12558 26146 0 _0088_
rlabel metal1 26546 35054 26546 35054 0 _0089_
rlabel metal1 11776 33082 11776 33082 0 _0090_
rlabel metal1 18625 35054 18625 35054 0 _0091_
rlabel metal2 15594 34850 15594 34850 0 _0092_
rlabel metal2 7406 9350 7406 9350 0 _0093_
rlabel metal2 15778 10914 15778 10914 0 _0094_
rlabel metal1 8321 13226 8321 13226 0 _0095_
rlabel metal2 23506 12002 23506 12002 0 _0096_
rlabel metal1 7815 14994 7815 14994 0 _0097_
rlabel metal1 25893 15402 25893 15402 0 _0098_
rlabel metal1 16371 19754 16371 19754 0 _0099_
rlabel metal2 27646 21794 27646 21794 0 _0100_
rlabel metal2 9062 23222 9062 23222 0 _0101_
rlabel via1 21753 23086 21753 23086 0 _0102_
rlabel metal2 14674 25670 14674 25670 0 _0103_
rlabel metal2 10166 25058 10166 25058 0 _0104_
rlabel metal1 26787 33558 26787 33558 0 _0105_
rlabel metal2 15778 29410 15778 29410 0 _0106_
rlabel via1 27641 33966 27641 33966 0 _0107_
rlabel metal2 7406 33762 7406 33762 0 _0108_
rlabel via1 16049 10030 16049 10030 0 _0109_
rlabel metal1 20020 10642 20020 10642 0 _0110_
rlabel metal2 6394 14178 6394 14178 0 _0111_
rlabel metal1 29766 10710 29766 10710 0 _0112_
rlabel metal1 6762 15674 6762 15674 0 _0113_
rlabel metal2 28474 15878 28474 15878 0 _0114_
rlabel metal1 15359 18734 15359 18734 0 _0115_
rlabel metal2 19642 21318 19642 21318 0 _0116_
rlabel metal2 5842 21318 5842 21318 0 _0117_
rlabel metal1 28929 25194 28929 25194 0 _0118_
rlabel metal1 5653 27370 5653 27370 0 _0119_
rlabel metal1 8735 24854 8735 24854 0 _0120_
rlabel metal2 28566 29410 28566 29410 0 _0121_
rlabel metal1 9062 33626 9062 33626 0 _0122_
rlabel metal2 17802 31586 17802 31586 0 _0123_
rlabel metal2 13202 34374 13202 34374 0 _0124_
rlabel metal1 11132 9146 11132 9146 0 _0125_
rlabel metal2 4922 11526 4922 11526 0 _0126_
rlabel metal1 9747 13974 9747 13974 0 _0127_
rlabel via1 27273 12818 27273 12818 0 _0128_
rlabel metal2 15778 16966 15778 16966 0 _0129_
rlabel via1 30033 13906 30033 13906 0 _0130_
rlabel metal2 10350 18530 10350 18530 0 _0131_
rlabel metal1 24978 20298 24978 20298 0 _0132_
rlabel metal1 4779 23766 4779 23766 0 _0133_
rlabel metal1 30406 26010 30406 26010 0 _0134_
rlabel metal1 18165 25262 18165 25262 0 _0135_
rlabel metal2 27646 28322 27646 28322 0 _0136_
rlabel metal2 22126 34374 22126 34374 0 _0137_
rlabel metal2 9614 34850 9614 34850 0 _0138_
rlabel metal2 20194 34850 20194 34850 0 _0139_
rlabel metal2 5474 33286 5474 33286 0 _0140_
rlabel metal1 8597 7378 8597 7378 0 _0141_
rlabel metal1 20143 8874 20143 8874 0 _0142_
rlabel metal1 12742 13498 12742 13498 0 _0143_
rlabel metal1 22172 11322 22172 11322 0 _0144_
rlabel metal2 8050 16354 8050 16354 0 _0145_
rlabel metal2 18078 16966 18078 16966 0 _0146_
rlabel metal2 12466 20570 12466 20570 0 _0147_
rlabel metal2 27830 20706 27830 20706 0 _0148_
rlabel metal2 12742 22882 12742 22882 0 _0149_
rlabel metal2 27002 25058 27002 25058 0 _0150_
rlabel metal1 8132 26962 8132 26962 0 _0151_
rlabel metal1 7355 25262 7355 25262 0 _0152_
rlabel metal1 24656 34714 24656 34714 0 _0153_
rlabel metal2 8142 34850 8142 34850 0 _0154_
rlabel via1 27641 35054 27641 35054 0 _0155_
rlabel metal1 8643 32402 8643 32402 0 _0156_
rlabel metal2 8970 9350 8970 9350 0 _0157_
rlabel metal1 3772 11322 3772 11322 0 _0158_
rlabel metal1 17986 11322 17986 11322 0 _0159_
rlabel metal2 25530 13090 25530 13090 0 _0160_
rlabel metal1 9747 17238 9747 17238 0 _0161_
rlabel metal2 25254 14790 25254 14790 0 _0162_
rlabel metal2 5382 19618 5382 19618 0 _0163_
rlabel metal2 27002 20706 27002 20706 0 _0164_
rlabel metal2 14858 21726 14858 21726 0 _0165_
rlabel metal2 24610 26758 24610 26758 0 _0166_
rlabel metal1 14623 24786 14623 24786 0 _0167_
rlabel metal1 3399 24786 3399 24786 0 _0168_
rlabel metal1 23000 31994 23000 31994 0 _0169_
rlabel metal1 3859 32402 3859 32402 0 _0170_
rlabel metal2 21482 32402 21482 32402 0 _0171_
rlabel metal2 14490 32674 14490 32674 0 _0172_
rlabel metal1 7033 7378 7033 7378 0 _0173_
rlabel metal2 14214 7990 14214 7990 0 _0174_
rlabel metal2 12374 11526 12374 11526 0 _0175_
rlabel metal1 26583 8874 26583 8874 0 _0176_
rlabel metal1 13979 16150 13979 16150 0 _0177_
rlabel metal2 21850 15266 21850 15266 0 _0178_
rlabel metal1 8505 18326 8505 18326 0 _0179_
rlabel metal1 20480 18734 20480 18734 0 _0180_
rlabel metal1 7697 21590 7697 21590 0 _0181_
rlabel metal2 24886 25670 24886 25670 0 _0182_
rlabel metal2 19734 25058 19734 25058 0 _0183_
rlabel metal2 27370 26758 27370 26758 0 _0184_
rlabel metal1 23179 28526 23179 28526 0 _0185_
rlabel metal1 13887 29206 13887 29206 0 _0186_
rlabel metal2 20286 28934 20286 28934 0 _0187_
rlabel metal2 7406 29410 7406 29410 0 _0188_
rlabel viali 5561 8942 5561 8942 0 _0189_
rlabel metal1 3189 10710 3189 10710 0 _0190_
rlabel metal1 4048 12954 4048 12954 0 _0191_
rlabel metal1 29680 9554 29680 9554 0 _0192_
rlabel metal2 4094 16694 4094 16694 0 _0193_
rlabel metal2 20102 15878 20102 15878 0 _0194_
rlabel metal1 3864 18394 3864 18394 0 _0195_
rlabel metal2 30590 22406 30590 22406 0 _0196_
rlabel metal1 3496 21862 3496 21862 0 _0197_
rlabel metal1 29256 23290 29256 23290 0 _0198_
rlabel metal2 6854 27234 6854 27234 0 _0199_
rlabel metal2 6394 25058 6394 25058 0 _0200_
rlabel metal2 29762 28934 29762 28934 0 _0201_
rlabel metal1 3828 31314 3828 31314 0 _0202_
rlabel metal1 27043 31722 27043 31722 0 _0203_
rlabel metal1 6159 31790 6159 31790 0 _0204_
rlabel metal1 6711 11050 6711 11050 0 _0205_
rlabel metal1 13473 9962 13473 9962 0 _0206_
rlabel metal2 10994 11526 10994 11526 0 _0207_
rlabel metal1 21293 13226 21293 13226 0 _0208_
rlabel metal2 9982 15266 9982 15266 0 _0209_
rlabel metal2 17986 15266 17986 15266 0 _0210_
rlabel metal1 6527 18666 6527 18666 0 _0211_
rlabel metal1 22310 21896 22310 21896 0 _0212_
rlabel metal2 7222 23460 7222 23460 0 _0213_
rlabel metal2 21850 25058 21850 25058 0 _0214_
rlabel metal1 13795 27030 13795 27030 0 _0215_
rlabel metal2 12190 27812 12190 27812 0 _0216_
rlabel metal2 23322 34850 23322 34850 0 _0217_
rlabel via1 11357 34986 11357 34986 0 _0218_
rlabel via1 17705 33966 17705 33966 0 _0219_
rlabel via1 13749 34578 13749 34578 0 _0220_
rlabel metal2 10074 7174 10074 7174 0 _0221_
rlabel metal1 11592 6970 11592 6970 0 _0222_
rlabel metal1 16463 11118 16463 11118 0 _0223_
rlabel metal1 27508 10234 27508 10234 0 _0224_
rlabel metal2 14674 14790 14674 14790 0 _0225_
rlabel metal1 27048 14586 27048 14586 0 _0226_
rlabel metal2 10350 20706 10350 20706 0 _0227_
rlabel metal1 22259 19414 22259 19414 0 _0228_
rlabel metal2 14858 22882 14858 22882 0 _0229_
rlabel metal1 27232 23290 27232 23290 0 _0230_
rlabel metal2 18998 27234 18998 27234 0 _0231_
rlabel metal2 25622 27846 25622 27846 0 _0232_
rlabel metal1 24472 32266 24472 32266 0 _0233_
rlabel metal2 14582 30498 14582 30498 0 _0234_
rlabel metal2 19642 32674 19642 32674 0 _0235_
rlabel metal1 12742 31994 12742 31994 0 _0236_
rlabel via1 4089 8942 4089 8942 0 _0237_
rlabel metal1 3741 9622 3741 9622 0 _0238_
rlabel metal2 17342 13702 17342 13702 0 _0239_
rlabel metal1 23777 14314 23777 14314 0 _0240_
rlabel metal2 2898 15266 2898 15266 0 _0241_
rlabel metal1 19867 14382 19867 14382 0 _0242_
rlabel metal1 8689 20502 8689 20502 0 _0243_
rlabel metal1 23961 21590 23961 21590 0 _0244_
rlabel metal2 10442 22236 10442 22236 0 _0245_
rlabel metal2 23138 25058 23138 25058 0 _0246_
rlabel metal2 16790 27846 16790 27846 0 _0247_
rlabel metal2 2622 27234 2622 27234 0 _0248_
rlabel metal2 24702 29410 24702 29410 0 _0249_
rlabel metal2 3082 29410 3082 29410 0 _0250_
rlabel metal2 17434 29410 17434 29410 0 _0251_
rlabel metal1 6348 29002 6348 29002 0 _0252_
rlabel metal2 7682 11526 7682 11526 0 _0253_
rlabel metal2 20654 9826 20654 9826 0 _0254_
rlabel metal2 6394 13090 6394 13090 0 _0255_
rlabel metal2 29118 11526 29118 11526 0 _0256_
rlabel metal2 14674 17442 14674 17442 0 _0257_
rlabel metal2 28474 13736 28474 13736 0 _0258_
rlabel via1 13381 18326 13381 18326 0 _0259_
rlabel metal1 23000 20570 23000 20570 0 _0260_
rlabel metal1 4140 21114 4140 21114 0 _0261_
rlabel metal2 22862 26758 22862 26758 0 _0262_
rlabel metal2 15134 26962 15134 26962 0 _0263_
rlabel metal2 4554 25058 4554 25058 0 _0264_
rlabel metal2 25162 31110 25162 31110 0 _0265_
rlabel metal2 4278 29410 4278 29410 0 _0266_
rlabel metal1 28428 30906 28428 30906 0 _0267_
rlabel metal1 9011 31382 9011 31382 0 _0268_
rlabel metal1 9384 11322 9384 11322 0 _0269_
rlabel metal1 11806 9622 11806 9622 0 _0270_
rlabel metal2 15686 13090 15686 13090 0 _0271_
rlabel metal1 23271 13974 23271 13974 0 _0272_
rlabel metal1 6021 16558 6021 16558 0 _0273_
rlabel metal1 23961 16082 23961 16082 0 _0274_
rlabel metal2 7958 19142 7958 19142 0 _0275_
rlabel metal2 18262 19346 18262 19346 0 _0276_
rlabel metal1 5929 23086 5929 23086 0 _0277_
rlabel metal1 22954 23290 22954 23290 0 _0278_
rlabel metal2 19366 23256 19366 23256 0 _0279_
rlabel metal2 10166 27234 10166 27234 0 _0280_
rlabel metal2 22862 30498 22862 30498 0 _0281_
rlabel metal2 10166 29410 10166 29410 0 _0282_
rlabel metal2 19274 31076 19274 31076 0 _0283_
rlabel metal2 6302 31110 6302 31110 0 _0284_
rlabel metal1 21482 15334 21482 15334 0 _0285_
rlabel metal1 22218 13906 22218 13906 0 _0286_
rlabel metal1 25622 9520 25622 9520 0 _0287_
rlabel metal1 27278 9622 27278 9622 0 _0288_
rlabel metal2 24242 12308 24242 12308 0 _0289_
rlabel metal1 22816 10098 22816 10098 0 _0290_
rlabel metal1 23460 14994 23460 14994 0 _0291_
rlabel metal1 34270 5678 34270 5678 0 _0292_
rlabel metal1 25070 6970 25070 6970 0 _0293_
rlabel metal1 29440 18394 29440 18394 0 _0294_
rlabel metal2 32522 5814 32522 5814 0 _0295_
rlabel metal1 32200 6426 32200 6426 0 _0296_
rlabel metal1 33120 7378 33120 7378 0 _0297_
rlabel metal2 32614 6256 32614 6256 0 _0298_
rlabel metal2 32890 6239 32890 6239 0 _0299_
rlabel metal1 32522 6800 32522 6800 0 _0300_
rlabel metal1 28980 7446 28980 7446 0 _0301_
rlabel metal1 30406 3604 30406 3604 0 _0302_
rlabel metal1 31418 6766 31418 6766 0 _0303_
rlabel metal1 32062 6664 32062 6664 0 _0304_
rlabel metal1 31418 6324 31418 6324 0 _0305_
rlabel metal2 31326 6868 31326 6868 0 _0306_
rlabel metal2 31602 7616 31602 7616 0 _0307_
rlabel metal1 30222 6256 30222 6256 0 _0308_
rlabel metal1 29992 6834 29992 6834 0 _0309_
rlabel metal2 28842 6630 28842 6630 0 _0310_
rlabel metal1 29670 4658 29670 4658 0 _0311_
rlabel metal2 28750 4828 28750 4828 0 _0312_
rlabel metal1 29670 3570 29670 3570 0 _0313_
rlabel metal1 30452 5338 30452 5338 0 _0314_
rlabel metal2 32062 5202 32062 5202 0 _0315_
rlabel metal1 31878 4658 31878 4658 0 _0316_
rlabel metal1 32614 4250 32614 4250 0 _0317_
rlabel metal1 27232 19482 27232 19482 0 _0318_
rlabel metal1 26312 17850 26312 17850 0 _0319_
rlabel via2 25990 17867 25990 17867 0 _0320_
rlabel metal1 31372 15062 31372 15062 0 _0321_
rlabel via1 28661 14382 28661 14382 0 _0322_
rlabel metal1 22816 16082 22816 16082 0 _0323_
rlabel metal1 23644 17850 23644 17850 0 _0324_
rlabel metal1 30268 18598 30268 18598 0 _0325_
rlabel metal2 29946 17272 29946 17272 0 _0326_
rlabel metal1 27002 18768 27002 18768 0 _0327_
rlabel metal1 26864 15538 26864 15538 0 _0328_
rlabel metal1 26772 16558 26772 16558 0 _0329_
rlabel metal1 25438 18870 25438 18870 0 _0330_
rlabel metal1 25116 17238 25116 17238 0 _0331_
rlabel metal2 30498 15929 30498 15929 0 _0332_
rlabel metal1 28796 17646 28796 17646 0 _0333_
rlabel metal2 24426 17884 24426 17884 0 _0334_
rlabel metal1 25668 18054 25668 18054 0 _0335_
rlabel metal1 7176 10030 7176 10030 0 _0336_
rlabel metal2 10028 8942 10028 8942 0 _0337_
rlabel metal2 10718 11594 10718 11594 0 _0338_
rlabel metal2 17342 8874 17342 8874 0 _0339_
rlabel metal1 18032 8058 18032 8058 0 _0340_
rlabel metal1 10580 8602 10580 8602 0 _0341_
rlabel metal2 10074 9520 10074 9520 0 _0342_
rlabel metal1 9982 8976 9982 8976 0 _0343_
rlabel metal2 15594 8806 15594 8806 0 _0344_
rlabel metal2 34086 6817 34086 6817 0 _0345_
rlabel metal1 20470 8432 20470 8432 0 _0346_
rlabel metal1 4830 10642 4830 10642 0 _0347_
rlabel metal2 13938 11492 13938 11492 0 _0348_
rlabel metal1 21436 8602 21436 8602 0 _0349_
rlabel metal1 13662 9520 13662 9520 0 _0350_
rlabel metal1 13846 8942 13846 8942 0 _0351_
rlabel metal2 14950 9248 14950 9248 0 _0352_
rlabel metal1 15042 9554 15042 9554 0 _0353_
rlabel metal2 20010 9248 20010 9248 0 _0354_
rlabel metal2 34086 9163 34086 9163 0 _0355_
rlabel metal1 8786 12852 8786 12852 0 _0356_
rlabel metal1 18078 12750 18078 12750 0 _0357_
rlabel metal1 13432 13906 13432 13906 0 _0358_
rlabel metal1 18998 12784 18998 12784 0 _0359_
rlabel metal2 13294 13702 13294 13702 0 _0360_
rlabel metal2 7774 14212 7774 14212 0 _0361_
rlabel metal2 12282 13872 12282 13872 0 _0362_
rlabel metal1 10764 12954 10764 12954 0 _0363_
rlabel metal2 19090 12903 19090 12903 0 _0364_
rlabel metal2 34178 11169 34178 11169 0 _0365_
rlabel metal1 21873 12682 21873 12682 0 _0366_
rlabel metal2 26450 13668 26450 13668 0 _0367_
rlabel metal1 24426 12682 24426 12682 0 _0368_
rlabel metal1 26864 13158 26864 13158 0 _0369_
rlabel metal1 28934 9146 28934 9146 0 _0370_
rlabel metal1 28612 9894 28612 9894 0 _0371_
rlabel metal1 26634 11322 26634 11322 0 _0372_
rlabel metal2 26358 11764 26358 11764 0 _0373_
rlabel metal1 30222 12172 30222 12172 0 _0374_
rlabel metal2 31418 12036 31418 12036 0 _0375_
rlabel metal2 7590 15878 7590 15878 0 _0376_
rlabel metal1 9660 15470 9660 15470 0 _0377_
rlabel metal1 15410 16082 15410 16082 0 _0378_
rlabel metal2 15870 15674 15870 15674 0 _0379_
rlabel metal2 11546 15062 11546 15062 0 _0380_
rlabel metal2 7774 17476 7774 17476 0 _0381_
rlabel metal1 11546 14926 11546 14926 0 _0382_
rlabel metal1 11454 15062 11454 15062 0 _0383_
rlabel metal2 13754 15198 13754 15198 0 _0384_
rlabel metal1 32936 14586 32936 14586 0 _0385_
rlabel metal1 21942 16116 21942 16116 0 _0386_
rlabel metal1 20194 14994 20194 14994 0 _0387_
rlabel metal2 21482 15606 21482 15606 0 _0388_
rlabel metal1 22862 15946 22862 15946 0 _0389_
rlabel metal1 29118 15028 29118 15028 0 _0390_
rlabel metal2 29762 15946 29762 15946 0 _0391_
rlabel metal1 26910 16082 26910 16082 0 _0392_
rlabel metal1 28612 16218 28612 16218 0 _0393_
rlabel metal1 32338 15096 32338 15096 0 _0394_
rlabel metal1 32016 14994 32016 14994 0 _0395_
rlabel metal2 16698 19414 16698 19414 0 _0396_
rlabel metal2 17158 18938 17158 18938 0 _0397_
rlabel metal1 10304 19346 10304 19346 0 _0398_
rlabel metal1 10074 19176 10074 19176 0 _0399_
rlabel metal1 5796 19346 5796 19346 0 _0400_
rlabel metal1 10166 19312 10166 19312 0 _0401_
rlabel metal1 12926 19448 12926 19448 0 _0402_
rlabel metal1 10350 19414 10350 19414 0 _0403_
rlabel metal2 12834 19618 12834 19618 0 _0404_
rlabel via2 34178 18717 34178 18717 0 _0405_
rlabel metal1 29302 21522 29302 21522 0 _0406_
rlabel metal1 22402 21454 22402 21454 0 _0407_
rlabel metal2 29854 20910 29854 20910 0 _0408_
rlabel metal1 24288 20434 24288 20434 0 _0409_
rlabel metal1 23874 20230 23874 20230 0 _0410_
rlabel metal1 24104 19482 24104 19482 0 _0411_
rlabel metal1 21068 19822 21068 19822 0 _0412_
rlabel metal2 24058 20230 24058 20230 0 _0413_
rlabel metal1 29946 20332 29946 20332 0 _0414_
rlabel metal1 34178 19856 34178 19856 0 _0415_
rlabel metal1 14260 22746 14260 22746 0 _0416_
rlabel metal1 16882 22644 16882 22644 0 _0417_
rlabel metal1 7820 21114 7820 21114 0 _0418_
rlabel metal1 8188 22610 8188 22610 0 _0419_
rlabel metal1 7958 22440 7958 22440 0 _0420_
rlabel metal1 5382 21862 5382 21862 0 _0421_
rlabel metal1 10442 23052 10442 23052 0 _0422_
rlabel metal1 8970 22678 8970 22678 0 _0423_
rlabel metal1 9039 22474 9039 22474 0 _0424_
rlabel metal2 17434 22304 17434 22304 0 _0425_
rlabel metal1 30268 24378 30268 24378 0 _0426_
rlabel metal2 30866 24956 30866 24956 0 _0427_
rlabel metal1 27554 24208 27554 24208 0 _0428_
rlabel metal2 26910 24548 26910 24548 0 _0429_
rlabel metal1 25438 26316 25438 26316 0 _0430_
rlabel metal1 26450 24616 26450 24616 0 _0431_
rlabel metal1 22862 24310 22862 24310 0 _0432_
rlabel metal1 26450 24752 26450 24752 0 _0433_
rlabel metal1 30958 24684 30958 24684 0 _0434_
rlabel metal2 31418 24140 31418 24140 0 _0435_
rlabel metal2 16054 25908 16054 25908 0 _0436_
rlabel metal2 9062 27676 9062 27676 0 _0437_
rlabel metal1 19734 24378 19734 24378 0 _0438_
rlabel metal1 20240 26010 20240 26010 0 _0439_
rlabel metal2 17526 26350 17526 26350 0 _0440_
rlabel metal1 16882 26962 16882 26962 0 _0441_
rlabel metal2 17710 26656 17710 26656 0 _0442_
rlabel metal2 15870 26962 15870 26962 0 _0443_
rlabel metal1 19090 26554 19090 26554 0 _0444_
rlabel metal2 31878 26962 31878 26962 0 _0445_
rlabel metal2 27462 27642 27462 27642 0 _0446_
rlabel metal1 28842 26384 28842 26384 0 _0447_
rlabel metal2 11546 26554 11546 26554 0 _0448_
rlabel metal1 11960 26554 11960 26554 0 _0449_
rlabel metal2 4830 26860 4830 26860 0 _0450_
rlabel metal1 7820 26010 7820 26010 0 _0451_
rlabel metal2 9522 25670 9522 25670 0 _0452_
rlabel metal2 10626 26146 10626 26146 0 _0453_
rlabel via2 11730 26469 11730 26469 0 _0454_
rlabel metal2 33994 26758 33994 26758 0 _0455_
rlabel metal1 28796 29818 28796 29818 0 _0456_
rlabel metal1 28336 30090 28336 30090 0 _0457_
rlabel metal2 23690 30260 23690 30260 0 _0458_
rlabel metal1 25484 30838 25484 30838 0 _0459_
rlabel metal2 25898 33354 25898 33354 0 _0460_
rlabel metal2 26082 32368 26082 32368 0 _0461_
rlabel metal2 26496 32844 26496 32844 0 _0462_
rlabel metal1 25990 31450 25990 31450 0 _0463_
rlabel metal1 27140 31994 27140 31994 0 _0464_
rlabel metal1 33442 30226 33442 30226 0 _0465_
rlabel metal1 15134 29818 15134 29818 0 _0466_
rlabel metal1 16514 30090 16514 30090 0 _0467_
rlabel metal1 11086 30090 11086 30090 0 _0468_
rlabel metal1 11178 31144 11178 31144 0 _0469_
rlabel metal2 10258 33796 10258 33796 0 _0470_
rlabel metal2 11132 31314 11132 31314 0 _0471_
rlabel metal2 4830 30532 4830 30532 0 _0472_
rlabel metal1 8188 30838 8188 30838 0 _0473_
rlabel metal1 11914 31178 11914 31178 0 _0474_
rlabel metal1 34178 31212 34178 31212 0 _0475_
rlabel metal1 21344 33490 21344 33490 0 _0476_
rlabel metal1 28152 32538 28152 32538 0 _0477_
rlabel metal1 29486 33456 29486 33456 0 _0478_
rlabel metal2 21114 32368 21114 32368 0 _0479_
rlabel metal1 18676 30090 18676 30090 0 _0480_
rlabel metal1 20286 33422 20286 33422 0 _0481_
rlabel metal1 21436 32402 21436 32402 0 _0482_
rlabel metal2 21022 33014 21022 33014 0 _0483_
rlabel metal1 25806 33422 25806 33422 0 _0484_
rlabel metal1 32430 32844 32430 32844 0 _0485_
rlabel metal1 14996 33490 14996 33490 0 _0486_
rlabel metal2 17434 33082 17434 33082 0 _0487_
rlabel metal1 7498 31994 7498 31994 0 _0488_
rlabel metal1 10166 32980 10166 32980 0 _0489_
rlabel metal1 8878 31790 8878 31790 0 _0490_
rlabel metal2 9614 32538 9614 32538 0 _0491_
rlabel metal1 13432 30090 13432 30090 0 _0492_
rlabel metal1 12581 32878 12581 32878 0 _0493_
rlabel metal1 14030 32878 14030 32878 0 _0494_
rlabel metal2 34178 33014 34178 33014 0 _0495_
rlabel metal1 31326 18122 31326 18122 0 _0496_
rlabel metal1 31372 17646 31372 17646 0 _0497_
rlabel metal1 28704 16558 28704 16558 0 _0498_
rlabel metal1 23184 7378 23184 7378 0 _0499_
rlabel metal1 23736 5746 23736 5746 0 _0500_
rlabel metal2 23782 5882 23782 5882 0 _0501_
rlabel metal1 25622 6222 25622 6222 0 _0502_
rlabel metal1 23828 7514 23828 7514 0 _0503_
rlabel metal2 25346 9350 25346 9350 0 _0504_
rlabel metal1 22402 7752 22402 7752 0 _0505_
rlabel metal2 24426 9316 24426 9316 0 _0506_
rlabel metal1 23276 7514 23276 7514 0 _0507_
rlabel metal1 23598 9996 23598 9996 0 _0508_
rlabel metal1 18630 21964 18630 21964 0 _0509_
rlabel metal1 23644 7514 23644 7514 0 _0510_
rlabel metal1 24702 10030 24702 10030 0 _0511_
rlabel metal1 25024 12750 25024 12750 0 _0512_
rlabel metal1 25254 10234 25254 10234 0 _0513_
rlabel metal2 27968 12852 27968 12852 0 _0514_
rlabel metal1 20470 9486 20470 9486 0 _0515_
rlabel metal2 23230 8194 23230 8194 0 _0516_
rlabel metal1 25714 13974 25714 13974 0 _0517_
rlabel metal2 26358 26469 26358 26469 0 _0518_
rlabel metal3 9422 1156 9422 1156 0 clk
rlabel metal1 13616 16558 13616 16558 0 clknet_0_clk
rlabel metal1 15134 15402 15134 15402 0 clknet_2_0__leaf_clk
rlabel metal1 14214 21114 14214 21114 0 clknet_2_1__leaf_clk
rlabel metal1 32154 15402 32154 15402 0 clknet_2_2__leaf_clk
rlabel metal1 25576 21998 25576 21998 0 clknet_2_3__leaf_clk
rlabel metal1 2346 19380 2346 19380 0 clknet_leaf_0_clk
rlabel metal1 20838 22100 20838 22100 0 clknet_leaf_10_clk
rlabel metal2 21850 29920 21850 29920 0 clknet_leaf_11_clk
rlabel metal1 21850 34612 21850 34612 0 clknet_leaf_12_clk
rlabel metal2 32154 33150 32154 33150 0 clknet_leaf_13_clk
rlabel metal1 33028 25806 33028 25806 0 clknet_leaf_14_clk
rlabel metal1 32982 22066 32982 22066 0 clknet_leaf_15_clk
rlabel metal1 25346 20910 25346 20910 0 clknet_leaf_16_clk
rlabel metal2 20654 17680 20654 17680 0 clknet_leaf_17_clk
rlabel metal2 27002 13872 27002 13872 0 clknet_leaf_18_clk
rlabel metal1 32476 17646 32476 17646 0 clknet_leaf_19_clk
rlabel metal2 13110 16558 13110 16558 0 clknet_leaf_1_clk
rlabel metal2 32798 8126 32798 8126 0 clknet_leaf_20_clk
rlabel metal1 32706 4556 32706 4556 0 clknet_leaf_21_clk
rlabel metal2 18906 8160 18906 8160 0 clknet_leaf_22_clk
rlabel metal1 19964 13294 19964 13294 0 clknet_leaf_23_clk
rlabel metal2 17526 17374 17526 17374 0 clknet_leaf_24_clk
rlabel metal1 13156 12750 13156 12750 0 clknet_leaf_25_clk
rlabel metal2 15962 7072 15962 7072 0 clknet_leaf_26_clk
rlabel metal1 3864 8942 3864 8942 0 clknet_leaf_27_clk
rlabel metal2 5566 13804 5566 13804 0 clknet_leaf_28_clk
rlabel metal1 13570 20468 13570 20468 0 clknet_leaf_2_clk
rlabel metal1 7866 21556 7866 21556 0 clknet_leaf_3_clk
rlabel metal1 2438 23732 2438 23732 0 clknet_leaf_4_clk
rlabel metal2 2254 28560 2254 28560 0 clknet_leaf_5_clk
rlabel metal2 4830 32946 4830 32946 0 clknet_leaf_6_clk
rlabel metal1 7774 32436 7774 32436 0 clknet_leaf_7_clk
rlabel metal2 15134 34850 15134 34850 0 clknet_leaf_8_clk
rlabel metal2 18078 25636 18078 25636 0 clknet_leaf_9_clk
rlabel metal2 31326 8262 31326 8262 0 count\[0\]
rlabel metal2 31786 6477 31786 6477 0 count\[1\]
rlabel metal2 28842 6086 28842 6086 0 count\[2\]
rlabel metal2 30866 3706 30866 3706 0 count\[3\]
rlabel metal2 34454 4318 34454 4318 0 count\[4\]
rlabel metal1 35098 5134 35098 5134 0 empty_o
rlabel metal2 34362 3247 34362 3247 0 full_o
rlabel metal1 18630 7514 18630 7514 0 mem\[0\]\[0\]
rlabel metal1 20424 27642 20424 27642 0 mem\[0\]\[10\]
rlabel metal1 29302 27098 29302 27098 0 mem\[0\]\[11\]
rlabel metal1 31142 31450 31142 31450 0 mem\[0\]\[12\]
rlabel metal1 16928 31994 16928 31994 0 mem\[0\]\[13\]
rlabel metal1 30406 33082 30406 33082 0 mem\[0\]\[14\]
rlabel metal1 17894 33354 17894 33354 0 mem\[0\]\[15\]
rlabel metal2 21298 8398 21298 8398 0 mem\[0\]\[1\]
rlabel metal2 19734 13430 19734 13430 0 mem\[0\]\[2\]
rlabel metal2 30958 11900 30958 11900 0 mem\[0\]\[3\]
rlabel metal1 16192 15470 16192 15470 0 mem\[0\]\[4\]
rlabel metal1 31234 16082 31234 16082 0 mem\[0\]\[5\]
rlabel metal1 17710 18054 17710 18054 0 mem\[0\]\[6\]
rlabel metal1 30682 21114 30682 21114 0 mem\[0\]\[7\]
rlabel metal1 17204 21658 17204 21658 0 mem\[0\]\[8\]
rlabel metal2 31786 24582 31786 24582 0 mem\[0\]\[9\]
rlabel via1 6394 9554 6394 9554 0 mem\[10\]\[0\]
rlabel metal1 7544 27642 7544 27642 0 mem\[10\]\[10\]
rlabel metal1 6762 25160 6762 25160 0 mem\[10\]\[11\]
rlabel metal1 30360 29274 30360 29274 0 mem\[10\]\[12\]
rlabel metal2 5198 31076 5198 31076 0 mem\[10\]\[13\]
rlabel metal2 28566 32096 28566 32096 0 mem\[10\]\[14\]
rlabel metal1 6900 31994 6900 31994 0 mem\[10\]\[15\]
rlabel metal1 3726 10540 3726 10540 0 mem\[10\]\[1\]
rlabel metal1 4784 13158 4784 13158 0 mem\[10\]\[2\]
rlabel metal2 28934 9792 28934 9792 0 mem\[10\]\[3\]
rlabel metal1 4922 17272 4922 17272 0 mem\[10\]\[4\]
rlabel metal1 20608 15402 20608 15402 0 mem\[10\]\[5\]
rlabel metal1 4692 18598 4692 18598 0 mem\[10\]\[6\]
rlabel metal1 28842 22032 28842 22032 0 mem\[10\]\[7\]
rlabel metal2 4186 21760 4186 21760 0 mem\[10\]\[8\]
rlabel metal1 29854 23834 29854 23834 0 mem\[10\]\[9\]
rlabel metal2 7406 11696 7406 11696 0 mem\[11\]\[0\]
rlabel metal1 15410 27098 15410 27098 0 mem\[11\]\[10\]
rlabel metal2 11822 27642 11822 27642 0 mem\[11\]\[11\]
rlabel metal1 23644 34714 23644 34714 0 mem\[11\]\[12\]
rlabel metal1 11454 35666 11454 35666 0 mem\[11\]\[13\]
rlabel metal1 18584 34170 18584 34170 0 mem\[11\]\[14\]
rlabel metal1 14674 34714 14674 34714 0 mem\[11\]\[15\]
rlabel metal2 13938 10642 13938 10642 0 mem\[11\]\[1\]
rlabel metal2 11362 12036 11362 12036 0 mem\[11\]\[2\]
rlabel metal2 22218 13158 22218 13158 0 mem\[11\]\[3\]
rlabel metal2 10810 15232 10810 15232 0 mem\[11\]\[4\]
rlabel metal1 18952 15674 18952 15674 0 mem\[11\]\[5\]
rlabel metal2 7038 19176 7038 19176 0 mem\[11\]\[6\]
rlabel metal1 22448 21998 22448 21998 0 mem\[11\]\[7\]
rlabel metal1 8418 23120 8418 23120 0 mem\[11\]\[8\]
rlabel metal1 22264 24922 22264 24922 0 mem\[11\]\[9\]
rlabel metal1 10488 7514 10488 7514 0 mem\[12\]\[0\]
rlabel metal2 17526 27166 17526 27166 0 mem\[12\]\[10\]
rlabel metal2 26450 27642 26450 27642 0 mem\[12\]\[11\]
rlabel metal2 25806 32640 25806 32640 0 mem\[12\]\[12\]
rlabel via1 15594 30226 15594 30226 0 mem\[12\]\[13\]
rlabel metal1 20332 32742 20332 32742 0 mem\[12\]\[14\]
rlabel metal1 13386 32538 13386 32538 0 mem\[12\]\[15\]
rlabel metal1 12834 7514 12834 7514 0 mem\[12\]\[1\]
rlabel metal1 17112 11866 17112 11866 0 mem\[12\]\[2\]
rlabel metal2 27002 10880 27002 10880 0 mem\[12\]\[3\]
rlabel metal1 15594 15130 15594 15130 0 mem\[12\]\[4\]
rlabel metal2 28014 14586 28014 14586 0 mem\[12\]\[5\]
rlabel metal1 10948 20570 10948 20570 0 mem\[12\]\[6\]
rlabel metal1 23000 19482 23000 19482 0 mem\[12\]\[7\]
rlabel metal2 15686 22848 15686 22848 0 mem\[12\]\[8\]
rlabel metal1 27370 23086 27370 23086 0 mem\[12\]\[9\]
rlabel metal1 5336 9622 5336 9622 0 mem\[13\]\[0\]
rlabel metal1 17618 27438 17618 27438 0 mem\[13\]\[10\]
rlabel metal1 3864 27574 3864 27574 0 mem\[13\]\[11\]
rlabel metal1 26450 29818 26450 29818 0 mem\[13\]\[12\]
rlabel metal2 3634 30022 3634 30022 0 mem\[13\]\[13\]
rlabel metal2 18354 29376 18354 29376 0 mem\[13\]\[14\]
rlabel metal1 6808 29478 6808 29478 0 mem\[13\]\[15\]
rlabel metal1 4232 10030 4232 10030 0 mem\[13\]\[1\]
rlabel metal1 17848 13294 17848 13294 0 mem\[13\]\[2\]
rlabel metal1 24518 14382 24518 14382 0 mem\[13\]\[3\]
rlabel metal1 3818 15334 3818 15334 0 mem\[13\]\[4\]
rlabel via1 20930 14994 20930 14994 0 mem\[13\]\[5\]
rlabel metal1 9430 20570 9430 20570 0 mem\[13\]\[6\]
rlabel metal1 24932 21386 24932 21386 0 mem\[13\]\[7\]
rlabel metal1 11040 21998 11040 21998 0 mem\[13\]\[8\]
rlabel via1 24058 24786 24058 24786 0 mem\[13\]\[9\]
rlabel metal2 8418 11322 8418 11322 0 mem\[14\]\[0\]
rlabel metal2 15962 26826 15962 26826 0 mem\[14\]\[10\]
rlabel metal1 5244 25466 5244 25466 0 mem\[14\]\[11\]
rlabel metal2 25990 30906 25990 30906 0 mem\[14\]\[12\]
rlabel metal2 4646 29682 4646 29682 0 mem\[14\]\[13\]
rlabel metal1 28888 31450 28888 31450 0 mem\[14\]\[14\]
rlabel metal1 9430 31450 9430 31450 0 mem\[14\]\[15\]
rlabel via1 21390 9894 21390 9894 0 mem\[14\]\[1\]
rlabel metal2 6946 13736 6946 13736 0 mem\[14\]\[2\]
rlabel metal1 27002 11594 27002 11594 0 mem\[14\]\[3\]
rlabel metal2 14306 17408 14306 17408 0 mem\[14\]\[4\]
rlabel metal2 28290 14178 28290 14178 0 mem\[14\]\[5\]
rlabel metal1 14536 19346 14536 19346 0 mem\[14\]\[6\]
rlabel metal1 22724 20570 22724 20570 0 mem\[14\]\[7\]
rlabel metal2 4738 21760 4738 21760 0 mem\[14\]\[8\]
rlabel metal2 23690 26554 23690 26554 0 mem\[14\]\[9\]
rlabel metal2 9798 11322 9798 11322 0 mem\[15\]\[0\]
rlabel metal1 19964 23834 19964 23834 0 mem\[15\]\[10\]
rlabel metal1 11316 27098 11316 27098 0 mem\[15\]\[11\]
rlabel metal1 24104 30566 24104 30566 0 mem\[15\]\[12\]
rlabel metal1 10810 29818 10810 29818 0 mem\[15\]\[13\]
rlabel metal2 20010 30906 20010 30906 0 mem\[15\]\[14\]
rlabel metal1 7268 31450 7268 31450 0 mem\[15\]\[15\]
rlabel metal1 13202 9690 13202 9690 0 mem\[15\]\[1\]
rlabel metal2 16054 13056 16054 13056 0 mem\[15\]\[2\]
rlabel metal1 24610 13974 24610 13974 0 mem\[15\]\[3\]
rlabel metal2 6762 16966 6762 16966 0 mem\[15\]\[4\]
rlabel metal1 24656 15946 24656 15946 0 mem\[15\]\[5\]
rlabel metal1 8556 19142 8556 19142 0 mem\[15\]\[6\]
rlabel metal1 18860 19686 18860 19686 0 mem\[15\]\[7\]
rlabel metal1 6670 23222 6670 23222 0 mem\[15\]\[8\]
rlabel metal1 24150 23834 24150 23834 0 mem\[15\]\[9\]
rlabel metal2 18814 9690 18814 9690 0 mem\[1\]\[0\]
rlabel metal1 16790 26010 16790 26010 0 mem\[1\]\[10\]
rlabel metal2 13018 26214 13018 26214 0 mem\[1\]\[11\]
rlabel metal1 27416 29818 27416 29818 0 mem\[1\]\[12\]
rlabel metal1 11822 31654 11822 31654 0 mem\[1\]\[13\]
rlabel metal2 21298 30872 21298 30872 0 mem\[1\]\[14\]
rlabel metal1 13800 30294 13800 30294 0 mem\[1\]\[15\]
rlabel metal1 13018 8262 13018 8262 0 mem\[1\]\[1\]
rlabel metal1 11592 14042 11592 14042 0 mem\[1\]\[2\]
rlabel metal2 28382 8092 28382 8092 0 mem\[1\]\[3\]
rlabel metal2 11178 17442 11178 17442 0 mem\[1\]\[4\]
rlabel metal1 21114 17170 21114 17170 0 mem\[1\]\[5\]
rlabel metal1 13110 19414 13110 19414 0 mem\[1\]\[6\]
rlabel metal1 23920 18938 23920 18938 0 mem\[1\]\[7\]
rlabel metal1 11362 23596 11362 23596 0 mem\[1\]\[8\]
rlabel metal1 26174 22746 26174 22746 0 mem\[1\]\[9\]
rlabel metal1 16836 8602 16836 8602 0 mem\[2\]\[0\]
rlabel metal1 18630 23494 18630 23494 0 mem\[2\]\[10\]
rlabel metal2 4370 27200 4370 27200 0 mem\[2\]\[11\]
rlabel metal1 22816 29614 22816 29614 0 mem\[2\]\[12\]
rlabel metal1 9890 30226 9890 30226 0 mem\[2\]\[13\]
rlabel metal2 20654 29988 20654 29988 0 mem\[2\]\[14\]
rlabel metal1 13708 29614 13708 29614 0 mem\[2\]\[15\]
rlabel metal1 20746 7514 20746 7514 0 mem\[2\]\[1\]
rlabel metal1 3864 13498 3864 13498 0 mem\[2\]\[2\]
rlabel metal1 21160 12410 21160 12410 0 mem\[2\]\[3\]
rlabel metal1 4922 15334 4922 15334 0 mem\[2\]\[4\]
rlabel metal1 24518 16694 24518 16694 0 mem\[2\]\[5\]
rlabel metal1 4278 19244 4278 19244 0 mem\[2\]\[6\]
rlabel metal1 19780 21658 19780 21658 0 mem\[2\]\[7\]
rlabel metal1 4416 22746 4416 22746 0 mem\[2\]\[8\]
rlabel metal1 22356 27642 22356 27642 0 mem\[2\]\[9\]
rlabel metal1 17710 7752 17710 7752 0 mem\[3\]\[0\]
rlabel metal2 17158 25568 17158 25568 0 mem\[3\]\[10\]
rlabel metal2 12742 26486 12742 26486 0 mem\[3\]\[11\]
rlabel metal1 25760 35258 25760 35258 0 mem\[3\]\[12\]
rlabel metal1 12006 32878 12006 32878 0 mem\[3\]\[13\]
rlabel metal2 19090 35428 19090 35428 0 mem\[3\]\[14\]
rlabel metal2 16054 34816 16054 34816 0 mem\[3\]\[15\]
rlabel metal2 14674 7684 14674 7684 0 mem\[3\]\[1\]
rlabel metal1 14398 13362 14398 13362 0 mem\[3\]\[2\]
rlabel metal1 25944 11322 25944 11322 0 mem\[3\]\[3\]
rlabel metal2 12558 14926 12558 14926 0 mem\[3\]\[4\]
rlabel metal2 22126 17374 22126 17374 0 mem\[3\]\[5\]
rlabel metal1 14628 19686 14628 19686 0 mem\[3\]\[6\]
rlabel metal1 21666 19788 21666 19788 0 mem\[3\]\[7\]
rlabel metal1 13708 21862 13708 21862 0 mem\[3\]\[8\]
rlabel metal1 26174 24072 26174 24072 0 mem\[3\]\[9\]
rlabel metal1 8050 9690 8050 9690 0 mem\[4\]\[0\]
rlabel metal1 15686 25262 15686 25262 0 mem\[4\]\[10\]
rlabel metal1 10442 24922 10442 24922 0 mem\[4\]\[11\]
rlabel metal1 26450 32810 26450 32810 0 mem\[4\]\[12\]
rlabel metal1 16008 29274 16008 29274 0 mem\[4\]\[13\]
rlabel metal1 28428 34170 28428 34170 0 mem\[4\]\[14\]
rlabel metal1 7728 33626 7728 33626 0 mem\[4\]\[15\]
rlabel metal1 15318 11322 15318 11322 0 mem\[4\]\[1\]
rlabel metal1 8924 12818 8924 12818 0 mem\[4\]\[2\]
rlabel metal1 23920 12410 23920 12410 0 mem\[4\]\[3\]
rlabel metal1 9016 15130 9016 15130 0 mem\[4\]\[4\]
rlabel metal1 26634 15674 26634 15674 0 mem\[4\]\[5\]
rlabel metal1 17112 20026 17112 20026 0 mem\[4\]\[6\]
rlabel metal2 28566 21828 28566 21828 0 mem\[4\]\[7\]
rlabel metal2 10258 22916 10258 22916 0 mem\[4\]\[8\]
rlabel metal2 22310 23324 22310 23324 0 mem\[4\]\[9\]
rlabel metal1 17112 10234 17112 10234 0 mem\[5\]\[0\]
rlabel metal1 6440 28050 6440 28050 0 mem\[5\]\[10\]
rlabel viali 10074 25874 10074 25874 0 mem\[5\]\[11\]
rlabel metal1 29762 29750 29762 29750 0 mem\[5\]\[12\]
rlabel metal1 9246 33524 9246 33524 0 mem\[5\]\[13\]
rlabel metal2 18170 30804 18170 30804 0 mem\[5\]\[14\]
rlabel metal1 13478 33966 13478 33966 0 mem\[5\]\[15\]
rlabel metal1 19734 10778 19734 10778 0 mem\[5\]\[1\]
rlabel metal2 6762 14144 6762 14144 0 mem\[5\]\[2\]
rlabel metal1 29394 10438 29394 10438 0 mem\[5\]\[3\]
rlabel metal1 7498 15538 7498 15538 0 mem\[5\]\[4\]
rlabel metal1 29026 15402 29026 15402 0 mem\[5\]\[5\]
rlabel metal2 16330 19142 16330 19142 0 mem\[5\]\[6\]
rlabel metal2 20470 21114 20470 21114 0 mem\[5\]\[7\]
rlabel metal2 6210 21114 6210 21114 0 mem\[5\]\[8\]
rlabel metal1 29670 25262 29670 25262 0 mem\[5\]\[9\]
rlabel metal1 10074 9350 10074 9350 0 mem\[6\]\[0\]
rlabel metal2 19090 25670 19090 25670 0 mem\[6\]\[10\]
rlabel metal2 28014 28288 28014 28288 0 mem\[6\]\[11\]
rlabel metal2 23230 34170 23230 34170 0 mem\[6\]\[12\]
rlabel metal1 10442 34714 10442 34714 0 mem\[6\]\[13\]
rlabel metal1 20792 34714 20792 34714 0 mem\[6\]\[14\]
rlabel metal1 6486 32810 6486 32810 0 mem\[6\]\[15\]
rlabel metal2 5290 11322 5290 11322 0 mem\[6\]\[1\]
rlabel viali 10902 14382 10902 14382 0 mem\[6\]\[2\]
rlabel metal1 28106 12954 28106 12954 0 mem\[6\]\[3\]
rlabel metal1 16330 16558 16330 16558 0 mem\[6\]\[4\]
rlabel metal1 29946 14382 29946 14382 0 mem\[6\]\[5\]
rlabel metal1 10948 18598 10948 18598 0 mem\[6\]\[6\]
rlabel metal2 25346 20672 25346 20672 0 mem\[6\]\[7\]
rlabel metal2 5290 23086 5290 23086 0 mem\[6\]\[8\]
rlabel metal1 31096 26010 31096 26010 0 mem\[6\]\[9\]
rlabel metal1 9614 7854 9614 7854 0 mem\[7\]\[0\]
rlabel metal1 9200 27438 9200 27438 0 mem\[7\]\[10\]
rlabel metal2 8234 25670 8234 25670 0 mem\[7\]\[11\]
rlabel metal1 25392 34714 25392 34714 0 mem\[7\]\[12\]
rlabel metal1 9108 34578 9108 34578 0 mem\[7\]\[13\]
rlabel metal2 28750 35462 28750 35462 0 mem\[7\]\[14\]
rlabel metal1 9384 32538 9384 32538 0 mem\[7\]\[15\]
rlabel metal1 21022 8942 21022 8942 0 mem\[7\]\[1\]
rlabel metal2 13754 13498 13754 13498 0 mem\[7\]\[2\]
rlabel via1 23322 12818 23322 12818 0 mem\[7\]\[3\]
rlabel via1 8970 16082 8970 16082 0 mem\[7\]\[4\]
rlabel metal1 18676 16558 18676 16558 0 mem\[7\]\[5\]
rlabel metal1 13156 20434 13156 20434 0 mem\[7\]\[6\]
rlabel metal2 28934 20672 28934 20672 0 mem\[7\]\[7\]
rlabel metal2 13570 22780 13570 22780 0 mem\[7\]\[8\]
rlabel metal2 27370 25024 27370 25024 0 mem\[7\]\[9\]
rlabel metal1 10166 9690 10166 9690 0 mem\[8\]\[0\]
rlabel metal1 15364 24922 15364 24922 0 mem\[8\]\[10\]
rlabel metal1 4048 25942 4048 25942 0 mem\[8\]\[11\]
rlabel metal2 23506 31280 23506 31280 0 mem\[8\]\[12\]
rlabel via1 4922 30702 4922 30702 0 mem\[8\]\[13\]
rlabel metal2 21298 32572 21298 32572 0 mem\[8\]\[14\]
rlabel metal1 15180 32742 15180 32742 0 mem\[8\]\[15\]
rlabel metal1 4416 11118 4416 11118 0 mem\[8\]\[1\]
rlabel metal1 18722 11866 18722 11866 0 mem\[8\]\[2\]
rlabel metal2 26358 13056 26358 13056 0 mem\[8\]\[3\]
rlabel viali 10902 17646 10902 17646 0 mem\[8\]\[4\]
rlabel metal1 26588 15130 26588 15130 0 mem\[8\]\[5\]
rlabel viali 6486 19346 6486 19346 0 mem\[8\]\[6\]
rlabel metal2 27462 21352 27462 21352 0 mem\[8\]\[7\]
rlabel metal1 15916 21658 15916 21658 0 mem\[8\]\[8\]
rlabel viali 25530 26350 25530 26350 0 mem\[8\]\[9\]
rlabel metal1 7866 7854 7866 7854 0 mem\[9\]\[0\]
rlabel metal1 20056 24922 20056 24922 0 mem\[9\]\[10\]
rlabel metal2 27002 27200 27002 27200 0 mem\[9\]\[11\]
rlabel metal2 23690 28934 23690 28934 0 mem\[9\]\[12\]
rlabel metal1 14628 29138 14628 29138 0 mem\[9\]\[13\]
rlabel metal2 21114 28764 21114 28764 0 mem\[9\]\[14\]
rlabel metal1 8326 29478 8326 29478 0 mem\[9\]\[15\]
rlabel metal1 14766 8602 14766 8602 0 mem\[9\]\[1\]
rlabel metal2 13202 12002 13202 12002 0 mem\[9\]\[2\]
rlabel metal1 27324 8942 27324 8942 0 mem\[9\]\[3\]
rlabel metal1 14720 16082 14720 16082 0 mem\[9\]\[4\]
rlabel metal1 22632 15674 22632 15674 0 mem\[9\]\[5\]
rlabel metal1 9246 18666 9246 18666 0 mem\[9\]\[6\]
rlabel via1 19550 19346 19550 19346 0 mem\[9\]\[7\]
rlabel metal2 7498 21114 7498 21114 0 mem\[9\]\[8\]
rlabel metal1 25484 25670 25484 25670 0 mem\[9\]\[9\]
rlabel metal1 1748 7242 1748 7242 0 net1
rlabel metal2 3174 10863 3174 10863 0 net10
rlabel metal1 30084 14858 30084 14858 0 net100
rlabel metal2 20562 29767 20562 29767 0 net101
rlabel metal1 20654 22644 20654 22644 0 net102
rlabel metal1 15778 16150 15778 16150 0 net103
rlabel metal1 13156 32946 13156 32946 0 net104
rlabel metal1 28658 14790 28658 14790 0 net105
rlabel metal1 15318 33456 15318 33456 0 net106
rlabel metal1 6164 25670 6164 25670 0 net107
rlabel metal1 19366 13430 19366 13430 0 net108
rlabel metal1 17020 17714 17020 17714 0 net109
rlabel metal1 14490 14484 14490 14484 0 net11
rlabel metal1 17572 19142 17572 19142 0 net110
rlabel metal1 20194 24684 20194 24684 0 net111
rlabel via1 28752 33490 28752 33490 0 net112
rlabel metal1 27554 21080 27554 21080 0 net113
rlabel metal1 10810 19380 10810 19380 0 net114
rlabel metal1 20562 25670 20562 25670 0 net115
rlabel via2 17250 16541 17250 16541 0 net116
rlabel metal1 14950 13838 14950 13838 0 net117
rlabel metal1 15617 33490 15617 33490 0 net118
rlabel metal2 21758 19074 21758 19074 0 net119
rlabel metal1 1702 14858 1702 14858 0 net12
rlabel metal2 31970 6698 31970 6698 0 net120
rlabel metal1 34408 6766 34408 6766 0 net121
rlabel metal1 32660 18802 32660 18802 0 net122
rlabel metal1 34362 23698 34362 23698 0 net123
rlabel metal2 34454 32402 34454 32402 0 net124
rlabel metal2 33442 6562 33442 6562 0 net125
rlabel metal1 32062 6970 32062 6970 0 net126
rlabel metal1 33028 6766 33028 6766 0 net127
rlabel metal1 17250 32844 17250 32844 0 net128
rlabel metal2 28750 26826 28750 26826 0 net129
rlabel metal2 1610 16252 1610 16252 0 net13
rlabel metal1 32154 7514 32154 7514 0 net130
rlabel metal2 5612 21828 5612 21828 0 net131
rlabel metal1 19642 12682 19642 12682 0 net132
rlabel metal1 8832 29682 8832 29682 0 net133
rlabel metal1 17066 12920 17066 12920 0 net134
rlabel metal1 19504 24174 19504 24174 0 net135
rlabel metal1 20746 20298 20746 20298 0 net136
rlabel metal1 7590 17238 7590 17238 0 net137
rlabel metal1 8234 25670 8234 25670 0 net138
rlabel metal1 8924 17306 8924 17306 0 net139
rlabel metal2 1794 18224 1794 18224 0 net14
rlabel metal1 13064 15334 13064 15334 0 net140
rlabel metal2 14766 34068 14766 34068 0 net141
rlabel metal1 21528 12818 21528 12818 0 net142
rlabel metal1 14214 16762 14214 16762 0 net143
rlabel metal2 20010 20927 20010 20927 0 net144
rlabel metal1 23552 29614 23552 29614 0 net145
rlabel metal1 20194 20468 20194 20468 0 net146
rlabel metal1 15042 19278 15042 19278 0 net147
rlabel metal1 5428 26554 5428 26554 0 net148
rlabel metal1 22977 21522 22977 21522 0 net149
rlabel metal2 3818 20026 3818 20026 0 net15
rlabel via2 15318 16677 15318 16677 0 net150
rlabel metal1 19872 18666 19872 18666 0 net151
rlabel metal1 19044 32742 19044 32742 0 net152
rlabel metal1 32292 14790 32292 14790 0 net153
rlabel metal1 11362 19346 11362 19346 0 net154
rlabel metal1 13432 32878 13432 32878 0 net155
rlabel metal1 19458 16422 19458 16422 0 net156
rlabel metal1 20746 9928 20746 9928 0 net157
rlabel metal1 20654 28968 20654 28968 0 net158
rlabel metal1 21206 31314 21206 31314 0 net159
rlabel via2 1886 22491 1886 22491 0 net16
rlabel metal1 25530 19482 25530 19482 0 net160
rlabel metal1 22540 6630 22540 6630 0 net161
rlabel metal1 23414 8058 23414 8058 0 net162
rlabel metal2 23322 4624 23322 4624 0 net163
rlabel viali 22954 8943 22954 8943 0 net164
rlabel metal1 26266 18156 26266 18156 0 net165
rlabel metal1 27094 17578 27094 17578 0 net166
rlabel metal1 25530 19380 25530 19380 0 net167
rlabel metal1 27830 18768 27830 18768 0 net168
rlabel metal1 30406 19346 30406 19346 0 net169
rlabel metal1 1610 24072 1610 24072 0 net17
rlabel metal1 27186 19346 27186 19346 0 net170
rlabel metal2 25162 18020 25162 18020 0 net171
rlabel metal1 25576 19278 25576 19278 0 net172
rlabel metal1 28428 18734 28428 18734 0 net173
rlabel metal1 31970 18224 31970 18224 0 net174
rlabel metal2 26450 18972 26450 18972 0 net175
rlabel metal1 26403 19346 26403 19346 0 net176
rlabel metal2 32798 18938 32798 18938 0 net177
rlabel metal1 32384 19346 32384 19346 0 net178
rlabel metal1 9890 31450 9890 31450 0 net179
rlabel via2 1886 26299 1886 26299 0 net18
rlabel metal1 14628 32334 14628 32334 0 net180
rlabel metal2 7866 33082 7866 33082 0 net181
rlabel metal1 19412 34510 19412 34510 0 net182
rlabel metal1 18768 34102 18768 34102 0 net183
rlabel metal1 21574 31858 21574 31858 0 net184
rlabel metal1 19090 35462 19090 35462 0 net185
rlabel metal1 4554 31858 4554 31858 0 net186
rlabel via2 12098 32725 12098 32725 0 net187
rlabel metal1 15410 30362 15410 30362 0 net188
rlabel metal1 13570 30600 13570 30600 0 net189
rlabel metal2 1886 4896 1886 4896 0 net19
rlabel metal1 25668 30634 25668 30634 0 net190
rlabel metal1 23874 34578 23874 34578 0 net191
rlabel metal1 27508 33558 27508 33558 0 net192
rlabel metal1 8372 25942 8372 25942 0 net193
rlabel metal2 12926 26656 12926 26656 0 net194
rlabel metal2 29946 27608 29946 27608 0 net195
rlabel metal1 20148 24786 20148 24786 0 net196
rlabel metal1 17020 27302 17020 27302 0 net197
rlabel metal1 16054 28526 16054 28526 0 net198
rlabel metal1 8372 27506 8372 27506 0 net199
rlabel metal1 1610 3400 1610 3400 0 net2
rlabel metal1 34546 5168 34546 5168 0 net20
rlabel metal1 7820 11186 7820 11186 0 net200
rlabel metal1 9522 7718 9522 7718 0 net201
rlabel metal1 17020 8466 17020 8466 0 net202
rlabel metal2 25438 6630 25438 6630 0 net203
rlabel metal1 26043 5270 26043 5270 0 net204
rlabel metal1 33350 4488 33350 4488 0 net205
rlabel metal1 32614 5576 32614 5576 0 net206
rlabel metal1 33343 17578 33343 17578 0 net207
rlabel metal1 33028 12138 33028 12138 0 net208
rlabel metal2 32246 19278 32246 19278 0 net209
rlabel metal2 34086 4250 34086 4250 0 net21
rlabel metal2 33534 33150 33534 33150 0 net210
rlabel metal1 32660 20026 32660 20026 0 net211
rlabel metal1 21758 26350 21758 26350 0 net212
rlabel metal1 25622 21930 25622 21930 0 net213
rlabel metal1 29762 25330 29762 25330 0 net214
rlabel metal1 5474 20842 5474 20842 0 net215
rlabel metal1 8372 21658 8372 21658 0 net216
rlabel metal1 15640 21930 15640 21930 0 net217
rlabel metal1 14398 22542 14398 22542 0 net218
rlabel metal2 18722 19108 18722 19108 0 net219
rlabel metal1 34638 7174 34638 7174 0 net22
rlabel metal1 23460 21930 23460 21930 0 net220
rlabel metal1 18354 22032 18354 22032 0 net221
rlabel metal2 9430 19788 9430 19788 0 net222
rlabel metal1 17020 17646 17020 17646 0 net223
rlabel metal2 15962 19890 15962 19890 0 net224
rlabel metal2 12374 19550 12374 19550 0 net225
rlabel metal1 19182 17272 19182 17272 0 net226
rlabel metal2 22678 16694 22678 16694 0 net227
rlabel metal1 30498 14484 30498 14484 0 net228
rlabel metal1 19366 17510 19366 17510 0 net229
rlabel metal1 34592 26282 34592 26282 0 net23
rlabel metal1 7222 15402 7222 15402 0 net230
rlabel metal1 16652 15130 16652 15130 0 net231
rlabel metal2 15042 15266 15042 15266 0 net232
rlabel metal1 14122 16524 14122 16524 0 net233
rlabel metal2 20746 11696 20746 11696 0 net234
rlabel metal1 30360 10778 30360 10778 0 net235
rlabel metal1 26174 12682 26174 12682 0 net236
rlabel metal1 21850 12818 21850 12818 0 net237
rlabel metal1 15134 13158 15134 13158 0 net238
rlabel metal1 17664 13158 17664 13158 0 net239
rlabel metal2 34546 27846 34546 27846 0 net24
rlabel metal1 9476 13226 9476 13226 0 net240
rlabel metal1 13294 7718 13294 7718 0 net241
rlabel metal1 20700 10574 20700 10574 0 net242
rlabel via2 19642 11067 19642 11067 0 net243
rlabel metal1 34086 30294 34086 30294 0 net25
rlabel metal2 34546 31484 34546 31484 0 net26
rlabel metal1 33534 33286 33534 33286 0 net27
rlabel metal1 34454 33626 34454 33626 0 net28
rlabel metal1 34408 9146 34408 9146 0 net29
rlabel metal2 5106 10404 5106 10404 0 net3
rlabel metal1 34684 11050 34684 11050 0 net30
rlabel metal2 33902 12444 33902 12444 0 net31
rlabel metal1 34914 14790 34914 14790 0 net32
rlabel metal1 33810 15878 33810 15878 0 net33
rlabel metal2 34546 18428 34546 18428 0 net34
rlabel metal1 34868 20230 34868 20230 0 net35
rlabel metal2 34546 22406 34546 22406 0 net36
rlabel metal2 34546 23868 34546 23868 0 net37
rlabel metal1 16882 12682 16882 12682 0 net38
rlabel metal1 19918 22508 19918 22508 0 net39
rlabel metal1 6026 28118 6026 28118 0 net4
rlabel metal2 18906 18428 18906 18428 0 net40
rlabel metal1 14352 19278 14352 19278 0 net41
rlabel metal1 4922 29104 4922 29104 0 net42
rlabel metal1 21574 9486 21574 9486 0 net43
rlabel metal1 15778 18054 15778 18054 0 net44
rlabel metal1 3634 14926 3634 14926 0 net45
rlabel metal1 18032 13362 18032 13362 0 net46
rlabel metal1 15502 22032 15502 22032 0 net47
rlabel metal1 16100 14314 16100 14314 0 net48
rlabel metal2 15870 21080 15870 21080 0 net49
rlabel metal2 2898 29070 2898 29070 0 net5
rlabel metal1 25622 32334 25622 32334 0 net50
rlabel via2 15870 23613 15870 23613 0 net51
rlabel metal1 7820 18054 7820 18054 0 net52
rlabel metal1 14352 35122 14352 35122 0 net53
rlabel metal1 19826 34476 19826 34476 0 net54
rlabel metal1 4876 18190 4876 18190 0 net55
rlabel metal1 5934 31246 5934 31246 0 net56
rlabel via2 30774 21301 30774 21301 0 net57
rlabel metal2 16238 19108 16238 19108 0 net58
rlabel metal1 20838 28628 20838 28628 0 net59
rlabel metal1 2070 31790 2070 31790 0 net6
rlabel metal1 15962 15606 15962 15606 0 net60
rlabel metal1 20608 16966 20608 16966 0 net61
rlabel metal1 16146 21114 16146 21114 0 net62
rlabel metal1 17526 21318 17526 21318 0 net63
rlabel metal1 13202 20366 13202 20366 0 net64
rlabel metal2 17250 34952 17250 34952 0 net65
rlabel metal1 19458 16626 19458 16626 0 net66
rlabel metal1 15870 16626 15870 16626 0 net67
rlabel metal1 27922 13498 27922 13498 0 net68
rlabel via2 20838 34493 20838 34493 0 net69
rlabel metal1 2852 33830 2852 33830 0 net7
rlabel metal1 14812 12614 14812 12614 0 net70
rlabel metal1 20930 10540 20930 10540 0 net71
rlabel metal1 9890 26554 9890 26554 0 net72
rlabel metal1 18262 10642 18262 10642 0 net73
rlabel metal2 17204 20366 17204 20366 0 net74
rlabel metal1 14398 33456 14398 33456 0 net75
rlabel metal1 27692 33422 27692 33422 0 net76
rlabel metal1 21942 24106 21942 24106 0 net77
rlabel metal1 14904 19890 14904 19890 0 net78
rlabel metal1 16330 34510 16330 34510 0 net79
rlabel metal1 1610 35564 1610 35564 0 net8
rlabel metal1 19918 35564 19918 35564 0 net80
rlabel metal1 18722 21012 18722 21012 0 net81
rlabel metal1 18630 22576 18630 22576 0 net82
rlabel metal1 17020 8398 17020 8398 0 net83
rlabel metal1 12834 19686 12834 19686 0 net84
rlabel metal2 12742 31799 12742 31799 0 net85
rlabel metal1 20148 17102 20148 17102 0 net86
rlabel metal2 17618 14110 17618 14110 0 net87
rlabel metal2 17342 21148 17342 21148 0 net88
rlabel metal1 30590 31858 30590 31858 0 net89
rlabel metal2 3634 34748 3634 34748 0 net9
rlabel metal1 30544 16014 30544 16014 0 net90
rlabel metal1 16698 14348 16698 14348 0 net91
rlabel metal1 5152 28118 5152 28118 0 net92
rlabel metal2 19918 26928 19918 26928 0 net93
rlabel metal1 21068 21046 21068 21046 0 net94
rlabel metal2 14674 13277 14674 13277 0 net95
rlabel metal1 18906 16184 18906 16184 0 net96
rlabel metal1 13984 22678 13984 22678 0 net97
rlabel metal1 29716 17646 29716 17646 0 net98
rlabel metal1 17572 19482 17572 19482 0 net99
rlabel metal3 35244 6868 35244 6868 0 rd_data_o[0]
rlabel metal3 35290 25908 35290 25908 0 rd_data_o[10]
rlabel metal1 35098 27982 35098 27982 0 rd_data_o[11]
rlabel metal1 34454 30634 34454 30634 0 rd_data_o[12]
rlabel metal2 34822 31501 34822 31501 0 rd_data_o[13]
rlabel metal2 34362 33711 34362 33711 0 rd_data_o[14]
rlabel via2 34362 35581 34362 35581 0 rd_data_o[15]
rlabel metal2 34822 8653 34822 8653 0 rd_data_o[1]
rlabel metal2 34822 11169 34822 11169 0 rd_data_o[2]
rlabel metal1 35098 12750 35098 12750 0 rd_data_o[3]
rlabel metal1 34500 15402 34500 15402 0 rd_data_o[4]
rlabel metal2 34362 16439 34362 16439 0 rd_data_o[5]
rlabel via2 34822 18275 34822 18275 0 rd_data_o[6]
rlabel metal1 34822 20842 34822 20842 0 rd_data_o[7]
rlabel metal2 34822 22321 34822 22321 0 rd_data_o[8]
rlabel metal2 34822 23885 34822 23885 0 rd_data_o[9]
rlabel metal3 1004 6868 1004 6868 0 rd_en_i
rlabel metal1 32200 18394 32200 18394 0 rd_ptr\[0\]
rlabel metal2 31694 17340 31694 17340 0 rd_ptr\[1\]
rlabel metal2 32522 19380 32522 19380 0 rd_ptr\[2\]
rlabel metal2 30130 17748 30130 17748 0 rd_ptr\[3\]
rlabel metal1 1380 3502 1380 3502 0 rst_n
rlabel metal1 1380 8942 1380 8942 0 wr_data_i[0]
rlabel metal1 1380 28050 1380 28050 0 wr_data_i[10]
rlabel metal1 1380 30226 1380 30226 0 wr_data_i[11]
rlabel metal2 1426 31535 1426 31535 0 wr_data_i[12]
rlabel metal1 1380 33966 1380 33966 0 wr_data_i[13]
rlabel metal1 1380 35258 1380 35258 0 wr_data_i[14]
rlabel metal3 958 37332 958 37332 0 wr_data_i[15]
rlabel metal1 1380 11118 1380 11118 0 wr_data_i[1]
rlabel metal1 1380 12818 1380 12818 0 wr_data_i[2]
rlabel metal1 1380 14994 1380 14994 0 wr_data_i[3]
rlabel metal2 1426 16473 1426 16473 0 wr_data_i[4]
rlabel metal1 1380 18734 1380 18734 0 wr_data_i[5]
rlabel metal1 1380 20434 1380 20434 0 wr_data_i[6]
rlabel metal1 1426 22610 1426 22610 0 wr_data_i[7]
rlabel metal1 1334 24174 1334 24174 0 wr_data_i[8]
rlabel metal3 1004 25908 1004 25908 0 wr_data_i[9]
rlabel metal1 1426 5202 1426 5202 0 wr_en_i
rlabel metal2 23598 7378 23598 7378 0 wr_ptr\[0\]
rlabel metal1 23782 6732 23782 6732 0 wr_ptr\[1\]
rlabel metal2 24794 6052 24794 6052 0 wr_ptr\[2\]
rlabel metal2 26082 7174 26082 7174 0 wr_ptr\[3\]
<< properties >>
string FIXED_BBOX 0 0 36473 38617
<< end >>
