VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO acsu
  CLASS BLOCK ;
  FOREIGN acsu ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN bm_s0_s0_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END bm_s0_s0_i[0]
  PIN bm_s0_s0_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END bm_s0_s0_i[1]
  PIN bm_s0_s2_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END bm_s0_s2_i[0]
  PIN bm_s0_s2_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END bm_s0_s2_i[1]
  PIN bm_s1_s0_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END bm_s1_s0_i[0]
  PIN bm_s1_s0_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END bm_s1_s0_i[1]
  PIN bm_s1_s2_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END bm_s1_s2_i[0]
  PIN bm_s1_s2_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END bm_s1_s2_i[1]
  PIN bm_s2_s1_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END bm_s2_s1_i[0]
  PIN bm_s2_s1_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END bm_s2_s1_i[1]
  PIN bm_s2_s3_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END bm_s2_s3_i[0]
  PIN bm_s2_s3_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END bm_s2_s3_i[1]
  PIN bm_s3_s1_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END bm_s3_s1_i[0]
  PIN bm_s3_s1_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END bm_s3_s1_i[1]
  PIN bm_s3_s3_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END bm_s3_s3_i[0]
  PIN bm_s3_s3_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END bm_s3_s3_i[1]
  PIN dec_bits_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 96.000 12.280 100.000 12.880 ;
    END
  END dec_bits_o[0]
  PIN dec_bits_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 96.000 36.760 100.000 37.360 ;
    END
  END dec_bits_o[1]
  PIN dec_bits_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 96.000 61.240 100.000 61.840 ;
    END
  END dec_bits_o[2]
  PIN dec_bits_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 96.000 85.720 100.000 86.320 ;
    END
  END dec_bits_o[3]
  PIN pm_s0_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 6.990 96.000 7.270 100.000 ;
    END
  END pm_s0_i[0]
  PIN pm_s0_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 9.750 96.000 10.030 100.000 ;
    END
  END pm_s0_i[1]
  PIN pm_s0_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 12.510 96.000 12.790 100.000 ;
    END
  END pm_s0_i[2]
  PIN pm_s0_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 15.270 96.000 15.550 100.000 ;
    END
  END pm_s0_i[3]
  PIN pm_s0_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 18.030 96.000 18.310 100.000 ;
    END
  END pm_s0_i[4]
  PIN pm_s0_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 20.790 96.000 21.070 100.000 ;
    END
  END pm_s0_i[5]
  PIN pm_s0_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 23.550 96.000 23.830 100.000 ;
    END
  END pm_s0_i[6]
  PIN pm_s0_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 26.310 96.000 26.590 100.000 ;
    END
  END pm_s0_i[7]
  PIN pm_s0_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END pm_s0_o[0]
  PIN pm_s0_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END pm_s0_o[1]
  PIN pm_s0_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END pm_s0_o[2]
  PIN pm_s0_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END pm_s0_o[3]
  PIN pm_s0_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END pm_s0_o[4]
  PIN pm_s0_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END pm_s0_o[5]
  PIN pm_s0_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END pm_s0_o[6]
  PIN pm_s0_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END pm_s0_o[7]
  PIN pm_s1_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 29.070 96.000 29.350 100.000 ;
    END
  END pm_s1_i[0]
  PIN pm_s1_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 31.830 96.000 32.110 100.000 ;
    END
  END pm_s1_i[1]
  PIN pm_s1_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 34.590 96.000 34.870 100.000 ;
    END
  END pm_s1_i[2]
  PIN pm_s1_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 37.350 96.000 37.630 100.000 ;
    END
  END pm_s1_i[3]
  PIN pm_s1_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 40.110 96.000 40.390 100.000 ;
    END
  END pm_s1_i[4]
  PIN pm_s1_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 42.870 96.000 43.150 100.000 ;
    END
  END pm_s1_i[5]
  PIN pm_s1_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 45.630 96.000 45.910 100.000 ;
    END
  END pm_s1_i[6]
  PIN pm_s1_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 48.390 96.000 48.670 100.000 ;
    END
  END pm_s1_i[7]
  PIN pm_s1_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END pm_s1_o[0]
  PIN pm_s1_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END pm_s1_o[1]
  PIN pm_s1_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END pm_s1_o[2]
  PIN pm_s1_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END pm_s1_o[3]
  PIN pm_s1_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END pm_s1_o[4]
  PIN pm_s1_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END pm_s1_o[5]
  PIN pm_s1_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END pm_s1_o[6]
  PIN pm_s1_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END pm_s1_o[7]
  PIN pm_s2_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 51.150 96.000 51.430 100.000 ;
    END
  END pm_s2_i[0]
  PIN pm_s2_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 53.910 96.000 54.190 100.000 ;
    END
  END pm_s2_i[1]
  PIN pm_s2_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 56.670 96.000 56.950 100.000 ;
    END
  END pm_s2_i[2]
  PIN pm_s2_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 59.430 96.000 59.710 100.000 ;
    END
  END pm_s2_i[3]
  PIN pm_s2_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 62.190 96.000 62.470 100.000 ;
    END
  END pm_s2_i[4]
  PIN pm_s2_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 64.950 96.000 65.230 100.000 ;
    END
  END pm_s2_i[5]
  PIN pm_s2_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 67.710 96.000 67.990 100.000 ;
    END
  END pm_s2_i[6]
  PIN pm_s2_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 70.470 96.000 70.750 100.000 ;
    END
  END pm_s2_i[7]
  PIN pm_s2_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END pm_s2_o[0]
  PIN pm_s2_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END pm_s2_o[1]
  PIN pm_s2_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END pm_s2_o[2]
  PIN pm_s2_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END pm_s2_o[3]
  PIN pm_s2_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END pm_s2_o[4]
  PIN pm_s2_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END pm_s2_o[5]
  PIN pm_s2_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END pm_s2_o[6]
  PIN pm_s2_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END pm_s2_o[7]
  PIN pm_s3_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 73.230 96.000 73.510 100.000 ;
    END
  END pm_s3_i[0]
  PIN pm_s3_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 75.990 96.000 76.270 100.000 ;
    END
  END pm_s3_i[1]
  PIN pm_s3_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 78.750 96.000 79.030 100.000 ;
    END
  END pm_s3_i[2]
  PIN pm_s3_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 81.510 96.000 81.790 100.000 ;
    END
  END pm_s3_i[3]
  PIN pm_s3_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 84.270 96.000 84.550 100.000 ;
    END
  END pm_s3_i[4]
  PIN pm_s3_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 87.030 96.000 87.310 100.000 ;
    END
  END pm_s3_i[5]
  PIN pm_s3_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 89.790 96.000 90.070 100.000 ;
    END
  END pm_s3_i[6]
  PIN pm_s3_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 92.550 96.000 92.830 100.000 ;
    END
  END pm_s3_i[7]
  PIN pm_s3_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END pm_s3_o[0]
  PIN pm_s3_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END pm_s3_o[1]
  PIN pm_s3_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END pm_s3_o[2]
  PIN pm_s3_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END pm_s3_o[3]
  PIN pm_s3_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END pm_s3_o[4]
  PIN pm_s3_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END pm_s3_o[5]
  PIN pm_s3_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END pm_s3_o[6]
  PIN pm_s3_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END pm_s3_o[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 87.280 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 87.280 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 94.490 87.125 ;
      LAYER li1 ;
        RECT 5.520 10.795 94.300 87.125 ;
      LAYER met1 ;
        RECT 5.520 10.640 94.300 88.700 ;
      LAYER met2 ;
        RECT 5.610 95.720 6.710 96.000 ;
        RECT 7.550 95.720 9.470 96.000 ;
        RECT 10.310 95.720 12.230 96.000 ;
        RECT 13.070 95.720 14.990 96.000 ;
        RECT 15.830 95.720 17.750 96.000 ;
        RECT 18.590 95.720 20.510 96.000 ;
        RECT 21.350 95.720 23.270 96.000 ;
        RECT 24.110 95.720 26.030 96.000 ;
        RECT 26.870 95.720 28.790 96.000 ;
        RECT 29.630 95.720 31.550 96.000 ;
        RECT 32.390 95.720 34.310 96.000 ;
        RECT 35.150 95.720 37.070 96.000 ;
        RECT 37.910 95.720 39.830 96.000 ;
        RECT 40.670 95.720 42.590 96.000 ;
        RECT 43.430 95.720 45.350 96.000 ;
        RECT 46.190 95.720 48.110 96.000 ;
        RECT 48.950 95.720 50.870 96.000 ;
        RECT 51.710 95.720 53.630 96.000 ;
        RECT 54.470 95.720 56.390 96.000 ;
        RECT 57.230 95.720 59.150 96.000 ;
        RECT 59.990 95.720 61.910 96.000 ;
        RECT 62.750 95.720 64.670 96.000 ;
        RECT 65.510 95.720 67.430 96.000 ;
        RECT 68.270 95.720 70.190 96.000 ;
        RECT 71.030 95.720 72.950 96.000 ;
        RECT 73.790 95.720 75.710 96.000 ;
        RECT 76.550 95.720 78.470 96.000 ;
        RECT 79.310 95.720 81.230 96.000 ;
        RECT 82.070 95.720 83.990 96.000 ;
        RECT 84.830 95.720 86.750 96.000 ;
        RECT 87.590 95.720 89.510 96.000 ;
        RECT 90.350 95.720 92.270 96.000 ;
        RECT 5.610 4.280 92.820 95.720 ;
        RECT 5.610 4.000 6.710 4.280 ;
        RECT 7.550 4.000 9.470 4.280 ;
        RECT 10.310 4.000 12.230 4.280 ;
        RECT 13.070 4.000 14.990 4.280 ;
        RECT 15.830 4.000 17.750 4.280 ;
        RECT 18.590 4.000 20.510 4.280 ;
        RECT 21.350 4.000 23.270 4.280 ;
        RECT 24.110 4.000 26.030 4.280 ;
        RECT 26.870 4.000 28.790 4.280 ;
        RECT 29.630 4.000 31.550 4.280 ;
        RECT 32.390 4.000 34.310 4.280 ;
        RECT 35.150 4.000 37.070 4.280 ;
        RECT 37.910 4.000 39.830 4.280 ;
        RECT 40.670 4.000 42.590 4.280 ;
        RECT 43.430 4.000 45.350 4.280 ;
        RECT 46.190 4.000 48.110 4.280 ;
        RECT 48.950 4.000 50.870 4.280 ;
        RECT 51.710 4.000 53.630 4.280 ;
        RECT 54.470 4.000 56.390 4.280 ;
        RECT 57.230 4.000 59.150 4.280 ;
        RECT 59.990 4.000 61.910 4.280 ;
        RECT 62.750 4.000 64.670 4.280 ;
        RECT 65.510 4.000 67.430 4.280 ;
        RECT 68.270 4.000 70.190 4.280 ;
        RECT 71.030 4.000 72.950 4.280 ;
        RECT 73.790 4.000 75.710 4.280 ;
        RECT 76.550 4.000 78.470 4.280 ;
        RECT 79.310 4.000 81.230 4.280 ;
        RECT 82.070 4.000 83.990 4.280 ;
        RECT 84.830 4.000 86.750 4.280 ;
        RECT 87.590 4.000 89.510 4.280 ;
        RECT 90.350 4.000 92.270 4.280 ;
      LAYER met3 ;
        RECT 4.400 89.400 96.000 90.265 ;
        RECT 4.000 86.720 96.000 89.400 ;
        RECT 4.000 85.360 95.600 86.720 ;
        RECT 4.400 85.320 95.600 85.360 ;
        RECT 4.400 83.960 96.000 85.320 ;
        RECT 4.000 79.920 96.000 83.960 ;
        RECT 4.400 78.520 96.000 79.920 ;
        RECT 4.000 74.480 96.000 78.520 ;
        RECT 4.400 73.080 96.000 74.480 ;
        RECT 4.000 69.040 96.000 73.080 ;
        RECT 4.400 67.640 96.000 69.040 ;
        RECT 4.000 63.600 96.000 67.640 ;
        RECT 4.400 62.240 96.000 63.600 ;
        RECT 4.400 62.200 95.600 62.240 ;
        RECT 4.000 60.840 95.600 62.200 ;
        RECT 4.000 58.160 96.000 60.840 ;
        RECT 4.400 56.760 96.000 58.160 ;
        RECT 4.000 52.720 96.000 56.760 ;
        RECT 4.400 51.320 96.000 52.720 ;
        RECT 4.000 47.280 96.000 51.320 ;
        RECT 4.400 45.880 96.000 47.280 ;
        RECT 4.000 41.840 96.000 45.880 ;
        RECT 4.400 40.440 96.000 41.840 ;
        RECT 4.000 37.760 96.000 40.440 ;
        RECT 4.000 36.400 95.600 37.760 ;
        RECT 4.400 36.360 95.600 36.400 ;
        RECT 4.400 35.000 96.000 36.360 ;
        RECT 4.000 30.960 96.000 35.000 ;
        RECT 4.400 29.560 96.000 30.960 ;
        RECT 4.000 25.520 96.000 29.560 ;
        RECT 4.400 24.120 96.000 25.520 ;
        RECT 4.000 20.080 96.000 24.120 ;
        RECT 4.400 18.680 96.000 20.080 ;
        RECT 4.000 14.640 96.000 18.680 ;
        RECT 4.400 13.280 96.000 14.640 ;
        RECT 4.400 13.240 95.600 13.280 ;
        RECT 4.000 11.880 95.600 13.240 ;
        RECT 4.000 9.200 96.000 11.880 ;
        RECT 4.400 8.335 96.000 9.200 ;
      LAYER met4 ;
        RECT 44.455 12.415 45.705 76.665 ;
  END
END acsu
END LIBRARY

