module tbu (clk,
    decoded_bit_o,
    rst_n,
    valid_i,
    valid_o,
    dec_bits_i,
    pm_new_s0_i,
    pm_new_s1_i,
    pm_new_s2_i,
    pm_new_s3_i);
 input clk;
 output decoded_bit_o;
 input rst_n;
 input valid_i;
 output valid_o;
 input [3:0] dec_bits_i;
 input [7:0] pm_new_s0_i;
 input [7:0] pm_new_s1_i;
 input [7:0] pm_new_s2_i;
 input [7:0] pm_new_s3_i;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire \history_s0[10] ;
 wire \history_s0[11] ;
 wire \history_s0[12] ;
 wire \history_s0[13] ;
 wire \history_s0[14] ;
 wire \history_s0[2] ;
 wire \history_s0[3] ;
 wire \history_s0[4] ;
 wire \history_s0[5] ;
 wire \history_s0[6] ;
 wire \history_s0[7] ;
 wire \history_s0[8] ;
 wire \history_s0[9] ;
 wire \history_s1[10] ;
 wire \history_s1[11] ;
 wire \history_s1[12] ;
 wire \history_s1[13] ;
 wire \history_s1[14] ;
 wire \history_s1[1] ;
 wire \history_s1[2] ;
 wire \history_s1[3] ;
 wire \history_s1[4] ;
 wire \history_s1[5] ;
 wire \history_s1[6] ;
 wire \history_s1[7] ;
 wire \history_s1[8] ;
 wire \history_s1[9] ;
 wire \history_s2[0] ;
 wire \history_s2[10] ;
 wire \history_s2[11] ;
 wire \history_s2[12] ;
 wire \history_s2[13] ;
 wire \history_s2[14] ;
 wire \history_s2[2] ;
 wire \history_s2[3] ;
 wire \history_s2[4] ;
 wire \history_s2[5] ;
 wire \history_s2[6] ;
 wire \history_s2[7] ;
 wire \history_s2[8] ;
 wire \history_s2[9] ;
 wire \history_s3[10] ;
 wire \history_s3[11] ;
 wire \history_s3[12] ;
 wire \history_s3[13] ;
 wire \history_s3[14] ;
 wire \history_s3[2] ;
 wire \history_s3[3] ;
 wire \history_s3[4] ;
 wire \history_s3[5] ;
 wire \history_s3[6] ;
 wire \history_s3[7] ;
 wire \history_s3[8] ;
 wire \history_s3[9] ;
 wire \latency_counter[0] ;
 wire \latency_counter[1] ;
 wire \latency_counter[2] ;
 wire \latency_counter[3] ;
 wire pipeline_full;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sky130_fd_sc_hd__inv_2 _247_ (.A(net55),
    .Y(_061_));
 sky130_fd_sc_hd__inv_2 _248_ (.A(net5),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _249_ (.A(net21),
    .Y(_063_));
 sky130_fd_sc_hd__inv_2 _250_ (.A(net6),
    .Y(_064_));
 sky130_fd_sc_hd__inv_2 _251_ (.A(net8),
    .Y(_065_));
 sky130_fd_sc_hd__inv_2 _252_ (.A(net76),
    .Y(_066_));
 sky130_fd_sc_hd__inv_2 _253_ (.A(net7),
    .Y(_067_));
 sky130_fd_sc_hd__inv_2 _254_ (.A(net12),
    .Y(_068_));
 sky130_fd_sc_hd__inv_2 _255_ (.A(net28),
    .Y(_069_));
 sky130_fd_sc_hd__inv_2 _256_ (.A(net11),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _257_ (.A(net27),
    .Y(_071_));
 sky130_fd_sc_hd__inv_2 _258_ (.A(net10),
    .Y(_072_));
 sky130_fd_sc_hd__inv_2 _259_ (.A(net26),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _260_ (.A(net9),
    .Y(_074_));
 sky130_fd_sc_hd__inv_2 _261_ (.A(net25),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _262_ (.A(net13),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _263_ (.A(net20),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _264_ (.A(net19),
    .Y(_078_));
 sky130_fd_sc_hd__inv_2 _265_ (.A(net18),
    .Y(_079_));
 sky130_fd_sc_hd__inv_2 _266_ (.A(net17),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _267_ (.A(net35),
    .Y(_081_));
 sky130_fd_sc_hd__inv_2 _268_ (.A(net32),
    .Y(_082_));
 sky130_fd_sc_hd__inv_2 _269_ (.A(net31),
    .Y(_083_));
 sky130_fd_sc_hd__and2_1 _270_ (.A(net55),
    .B(pipeline_full),
    .X(_000_));
 sky130_fd_sc_hd__and3b_1 _271_ (.A_N(\latency_counter[0] ),
    .B(\latency_counter[3] ),
    .C(net55),
    .X(_084_));
 sky130_fd_sc_hd__a31o_1 _272_ (.A1(\latency_counter[1] ),
    .A2(\latency_counter[2] ),
    .A3(_084_),
    .B1(pipeline_full),
    .X(_001_));
 sky130_fd_sc_hd__nand2b_1 _273_ (.A_N(net28),
    .B(net20),
    .Y(_085_));
 sky130_fd_sc_hd__nand2b_1 _274_ (.A_N(net27),
    .B(net19),
    .Y(_086_));
 sky130_fd_sc_hd__nand2_1 _275_ (.A(_085_),
    .B(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__nand2b_1 _276_ (.A_N(net20),
    .B(net28),
    .Y(_088_));
 sky130_fd_sc_hd__nand2_1 _277_ (.A(net26),
    .B(_079_),
    .Y(_089_));
 sky130_fd_sc_hd__nand2b_1 _278_ (.A_N(net19),
    .B(net27),
    .Y(_090_));
 sky130_fd_sc_hd__and4_1 _279_ (.A(_085_),
    .B(_086_),
    .C(_088_),
    .D(_090_),
    .X(_091_));
 sky130_fd_sc_hd__o22a_1 _280_ (.A1(net26),
    .A2(_079_),
    .B1(_080_),
    .B2(net25),
    .X(_092_));
 sky130_fd_sc_hd__a22o_1 _281_ (.A1(_073_),
    .A2(net18),
    .B1(net17),
    .B2(_075_),
    .X(_093_));
 sky130_fd_sc_hd__o2111a_1 _282_ (.A1(_075_),
    .A2(net17),
    .B1(_089_),
    .C1(_091_),
    .D1(_092_),
    .X(_094_));
 sky130_fd_sc_hd__nand2b_1 _283_ (.A_N(net76),
    .B(net80),
    .Y(_095_));
 sky130_fd_sc_hd__nand2b_1 _284_ (.A_N(net80),
    .B(net76),
    .Y(_096_));
 sky130_fd_sc_hd__xnor2_1 _285_ (.A(net23),
    .B(net15),
    .Y(_097_));
 sky130_fd_sc_hd__and3_1 _286_ (.A(_095_),
    .B(_096_),
    .C(_097_),
    .X(_098_));
 sky130_fd_sc_hd__nand2b_1 _287_ (.A_N(net22),
    .B(net14),
    .Y(_099_));
 sky130_fd_sc_hd__nand2b_1 _288_ (.A_N(net14),
    .B(net22),
    .Y(_100_));
 sky130_fd_sc_hd__nand2b_1 _289_ (.A_N(net13),
    .B(net21),
    .Y(_101_));
 sky130_fd_sc_hd__and3_1 _290_ (.A(_099_),
    .B(_100_),
    .C(_101_),
    .X(_102_));
 sky130_fd_sc_hd__a21bo_1 _291_ (.A1(_100_),
    .A2(_101_),
    .B1_N(_099_),
    .X(_103_));
 sky130_fd_sc_hd__and3b_1 _292_ (.A_N(net23),
    .B(net15),
    .C(_096_),
    .X(_104_));
 sky130_fd_sc_hd__a221o_1 _293_ (.A1(_066_),
    .A2(net80),
    .B1(_098_),
    .B2(_103_),
    .C1(_104_),
    .X(_105_));
 sky130_fd_sc_hd__a32o_1 _294_ (.A1(_089_),
    .A2(_091_),
    .A3(_093_),
    .B1(_088_),
    .B2(_087_),
    .X(_106_));
 sky130_fd_sc_hd__a21oi_1 _295_ (.A1(_094_),
    .A2(_105_),
    .B1(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__o2111a_1 _296_ (.A1(net21),
    .A2(_076_),
    .B1(_094_),
    .C1(_098_),
    .D1(_102_),
    .X(_108_));
 sky130_fd_sc_hd__nand2b_1 _297_ (.A_N(net14),
    .B(net30),
    .Y(_109_));
 sky130_fd_sc_hd__nand2b_1 _298_ (.A_N(net13),
    .B(net29),
    .Y(_110_));
 sky130_fd_sc_hd__and2b_1 _299_ (.A_N(net30),
    .B(net14),
    .X(_111_));
 sky130_fd_sc_hd__a21o_1 _300_ (.A1(_109_),
    .A2(_110_),
    .B1(_111_),
    .X(_112_));
 sky130_fd_sc_hd__o22a_1 _301_ (.A1(_079_),
    .A2(net73),
    .B1(net33),
    .B2(_080_),
    .X(_113_));
 sky130_fd_sc_hd__and2b_1 _302_ (.A_N(net20),
    .B(net36),
    .X(_114_));
 sky130_fd_sc_hd__a21oi_1 _303_ (.A1(_080_),
    .A2(net33),
    .B1(_114_),
    .Y(_115_));
 sky130_fd_sc_hd__o22a_1 _304_ (.A1(_077_),
    .A2(net36),
    .B1(net35),
    .B2(_078_),
    .X(_116_));
 sky130_fd_sc_hd__o2bb2a_1 _305_ (.A1_N(net73),
    .A2_N(_079_),
    .B1(net19),
    .B2(_081_),
    .X(_117_));
 sky130_fd_sc_hd__a22o_1 _306_ (.A1(_078_),
    .A2(net35),
    .B1(net73),
    .B2(_079_),
    .X(_118_));
 sky130_fd_sc_hd__and4_1 _307_ (.A(_113_),
    .B(_115_),
    .C(_116_),
    .D(_117_),
    .X(_119_));
 sky130_fd_sc_hd__xnor2_1 _308_ (.A(net15),
    .B(net31),
    .Y(_120_));
 sky130_fd_sc_hd__nand2b_1 _309_ (.A_N(net80),
    .B(net32),
    .Y(_121_));
 sky130_fd_sc_hd__nand2b_1 _310_ (.A_N(net32),
    .B(net16),
    .Y(_122_));
 sky130_fd_sc_hd__and3_1 _311_ (.A(_120_),
    .B(_121_),
    .C(_122_),
    .X(_123_));
 sky130_fd_sc_hd__o21a_1 _312_ (.A1(_113_),
    .A2(_118_),
    .B1(_116_),
    .X(_124_));
 sky130_fd_sc_hd__and3_1 _313_ (.A(net15),
    .B(_083_),
    .C(_121_),
    .X(_125_));
 sky130_fd_sc_hd__a221o_1 _314_ (.A1(net16),
    .A2(_082_),
    .B1(_112_),
    .B2(_123_),
    .C1(_125_),
    .X(_126_));
 sky130_fd_sc_hd__o2bb2a_1 _315_ (.A1_N(_119_),
    .A2_N(_126_),
    .B1(_124_),
    .B2(_114_),
    .X(_127_));
 sky130_fd_sc_hd__o21ba_1 _316_ (.A1(_076_),
    .A2(net29),
    .B1_N(_111_),
    .X(_128_));
 sky130_fd_sc_hd__and3_1 _317_ (.A(_109_),
    .B(_110_),
    .C(_128_),
    .X(_129_));
 sky130_fd_sc_hd__and3_1 _318_ (.A(_119_),
    .B(_123_),
    .C(_129_),
    .X(_130_));
 sky130_fd_sc_hd__o22a_1 _319_ (.A1(_107_),
    .A2(_108_),
    .B1(_127_),
    .B2(_130_),
    .X(_131_));
 sky130_fd_sc_hd__and2b_1 _320_ (.A_N(net36),
    .B(net28),
    .X(_132_));
 sky130_fd_sc_hd__a22o_1 _321_ (.A1(_069_),
    .A2(net36),
    .B1(net35),
    .B2(_071_),
    .X(_133_));
 sky130_fd_sc_hd__a22o_1 _322_ (.A1(_073_),
    .A2(net73),
    .B1(net33),
    .B2(_075_),
    .X(_134_));
 sky130_fd_sc_hd__o22a_1 _323_ (.A1(_071_),
    .A2(net35),
    .B1(net34),
    .B2(_073_),
    .X(_135_));
 sky130_fd_sc_hd__a21oi_1 _324_ (.A1(_134_),
    .A2(_135_),
    .B1(_133_),
    .Y(_136_));
 sky130_fd_sc_hd__and2b_1 _325_ (.A_N(net30),
    .B(net22),
    .X(_137_));
 sky130_fd_sc_hd__and2b_1 _326_ (.A_N(net29),
    .B(net21),
    .X(_138_));
 sky130_fd_sc_hd__nand2b_1 _327_ (.A_N(net22),
    .B(net30),
    .Y(_139_));
 sky130_fd_sc_hd__o221a_1 _328_ (.A1(net23),
    .A2(_083_),
    .B1(_137_),
    .B2(_138_),
    .C1(_139_),
    .X(_140_));
 sky130_fd_sc_hd__a22o_1 _329_ (.A1(net76),
    .A2(_082_),
    .B1(_083_),
    .B2(net23),
    .X(_141_));
 sky130_fd_sc_hd__o22a_1 _330_ (.A1(net24),
    .A2(_082_),
    .B1(_140_),
    .B2(_141_),
    .X(_142_));
 sky130_fd_sc_hd__o21ba_1 _331_ (.A1(_075_),
    .A2(net33),
    .B1_N(_132_),
    .X(_143_));
 sky130_fd_sc_hd__or4bb_1 _332_ (.A(_133_),
    .B(_134_),
    .C_N(_135_),
    .D_N(_143_),
    .X(_144_));
 sky130_fd_sc_hd__o22a_1 _333_ (.A1(_132_),
    .A2(_136_),
    .B1(_142_),
    .B2(_144_),
    .X(_145_));
 sky130_fd_sc_hd__mux2_1 _334_ (.A0(\history_s2[14] ),
    .A1(\history_s3[14] ),
    .S(_145_),
    .X(_146_));
 sky130_fd_sc_hd__o22a_1 _335_ (.A1(_068_),
    .A2(net36),
    .B1(net35),
    .B2(_070_),
    .X(_147_));
 sky130_fd_sc_hd__o22a_1 _336_ (.A1(_072_),
    .A2(net73),
    .B1(net33),
    .B2(_074_),
    .X(_148_));
 sky130_fd_sc_hd__o22a_1 _337_ (.A1(_065_),
    .A2(net32),
    .B1(net31),
    .B2(_067_),
    .X(_149_));
 sky130_fd_sc_hd__nand2b_1 _338_ (.A_N(net30),
    .B(net6),
    .Y(_150_));
 sky130_fd_sc_hd__nand2b_1 _339_ (.A_N(net29),
    .B(net5),
    .Y(_151_));
 sky130_fd_sc_hd__and2b_1 _340_ (.A_N(net6),
    .B(net30),
    .X(_152_));
 sky130_fd_sc_hd__a221o_1 _341_ (.A1(_067_),
    .A2(net31),
    .B1(_150_),
    .B2(_151_),
    .C1(_152_),
    .X(_153_));
 sky130_fd_sc_hd__nor2_1 _342_ (.A(net8),
    .B(_082_),
    .Y(_154_));
 sky130_fd_sc_hd__a221o_1 _343_ (.A1(_074_),
    .A2(net33),
    .B1(_149_),
    .B2(_153_),
    .C1(_154_),
    .X(_155_));
 sky130_fd_sc_hd__nor2_1 _344_ (.A(net11),
    .B(_081_),
    .Y(_156_));
 sky130_fd_sc_hd__a221o_1 _345_ (.A1(_072_),
    .A2(net73),
    .B1(_148_),
    .B2(_155_),
    .C1(_156_),
    .X(_157_));
 sky130_fd_sc_hd__a22o_1 _346_ (.A1(_068_),
    .A2(net36),
    .B1(_147_),
    .B2(_157_),
    .X(_158_));
 sky130_fd_sc_hd__and2b_1 _347_ (.A_N(net10),
    .B(net26),
    .X(_159_));
 sky130_fd_sc_hd__and2b_1 _348_ (.A_N(net11),
    .B(net27),
    .X(_160_));
 sky130_fd_sc_hd__and2b_1 _349_ (.A_N(net12),
    .B(net28),
    .X(_161_));
 sky130_fd_sc_hd__a2111o_1 _350_ (.A1(_074_),
    .A2(net25),
    .B1(_159_),
    .C1(_160_),
    .D1(_161_),
    .X(_162_));
 sky130_fd_sc_hd__a22o_1 _351_ (.A1(net10),
    .A2(_073_),
    .B1(net9),
    .B2(_075_),
    .X(_163_));
 sky130_fd_sc_hd__a22o_1 _352_ (.A1(net12),
    .A2(_069_),
    .B1(net11),
    .B2(_071_),
    .X(_164_));
 sky130_fd_sc_hd__inv_2 _353_ (.A(_164_),
    .Y(_165_));
 sky130_fd_sc_hd__or3_1 _354_ (.A(_162_),
    .B(_163_),
    .C(_164_),
    .X(_166_));
 sky130_fd_sc_hd__nand2b_1 _355_ (.A_N(net76),
    .B(net8),
    .Y(_167_));
 sky130_fd_sc_hd__and2b_1 _356_ (.A_N(net8),
    .B(net76),
    .X(_168_));
 sky130_fd_sc_hd__xor2_1 _357_ (.A(net7),
    .B(net23),
    .X(_169_));
 sky130_fd_sc_hd__or3b_1 _358_ (.A(_169_),
    .B(_168_),
    .C_N(_167_),
    .X(_170_));
 sky130_fd_sc_hd__nand2b_1 _359_ (.A_N(net22),
    .B(net6),
    .Y(_171_));
 sky130_fd_sc_hd__nand2b_1 _360_ (.A_N(net6),
    .B(net22),
    .Y(_172_));
 sky130_fd_sc_hd__o211ai_1 _361_ (.A1(net5),
    .A2(_063_),
    .B1(_171_),
    .C1(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__a21o_1 _362_ (.A1(_171_),
    .A2(_173_),
    .B1(_170_),
    .X(_174_));
 sky130_fd_sc_hd__or3_1 _363_ (.A(_067_),
    .B(net23),
    .C(_168_),
    .X(_175_));
 sky130_fd_sc_hd__a31o_1 _364_ (.A1(_167_),
    .A2(_174_),
    .A3(_175_),
    .B1(_166_),
    .X(_176_));
 sky130_fd_sc_hd__or3b_1 _365_ (.A(_159_),
    .B(_160_),
    .C_N(_163_),
    .X(_177_));
 sky130_fd_sc_hd__a21o_1 _366_ (.A1(_165_),
    .A2(_177_),
    .B1(_161_),
    .X(_178_));
 sky130_fd_sc_hd__a211o_1 _367_ (.A1(net5),
    .A2(_063_),
    .B1(_170_),
    .C1(_173_),
    .X(_179_));
 sky130_fd_sc_hd__a2bb2o_1 _368_ (.A1_N(_166_),
    .A2_N(_179_),
    .B1(_178_),
    .B2(_176_),
    .X(_180_));
 sky130_fd_sc_hd__nand2_1 _369_ (.A(net12),
    .B(_077_),
    .Y(_181_));
 sky130_fd_sc_hd__o22a_1 _370_ (.A1(_070_),
    .A2(net19),
    .B1(net18),
    .B2(_072_),
    .X(_182_));
 sky130_fd_sc_hd__a22o_1 _371_ (.A1(_072_),
    .A2(net18),
    .B1(net17),
    .B2(_074_),
    .X(_183_));
 sky130_fd_sc_hd__a211o_1 _372_ (.A1(_064_),
    .A2(net14),
    .B1(net13),
    .C1(_062_),
    .X(_184_));
 sky130_fd_sc_hd__o22a_1 _373_ (.A1(_064_),
    .A2(net14),
    .B1(net15),
    .B2(_067_),
    .X(_185_));
 sky130_fd_sc_hd__a22o_1 _374_ (.A1(_065_),
    .A2(net80),
    .B1(net15),
    .B2(_067_),
    .X(_186_));
 sky130_fd_sc_hd__a21o_1 _375_ (.A1(_184_),
    .A2(_185_),
    .B1(_186_),
    .X(_187_));
 sky130_fd_sc_hd__o221a_1 _376_ (.A1(_065_),
    .A2(net80),
    .B1(net17),
    .B2(_074_),
    .C1(_187_),
    .X(_188_));
 sky130_fd_sc_hd__o21a_1 _377_ (.A1(_183_),
    .A2(_188_),
    .B1(_182_),
    .X(_189_));
 sky130_fd_sc_hd__a22o_1 _378_ (.A1(_068_),
    .A2(net20),
    .B1(net19),
    .B2(_070_),
    .X(_190_));
 sky130_fd_sc_hd__o2111a_1 _379_ (.A1(_189_),
    .A2(_190_),
    .B1(_158_),
    .C1(_180_),
    .D1(_181_),
    .X(_191_));
 sky130_fd_sc_hd__mux2_1 _380_ (.A0(_146_),
    .A1(\history_s1[14] ),
    .S(_131_),
    .X(_192_));
 sky130_fd_sc_hd__mux2_1 _381_ (.A0(_192_),
    .A1(\history_s0[14] ),
    .S(_191_),
    .X(_193_));
 sky130_fd_sc_hd__mux2_1 _382_ (.A0(net39),
    .A1(_193_),
    .S(_000_),
    .X(_002_));
 sky130_fd_sc_hd__and2_1 _383_ (.A(net53),
    .B(\history_s1[1] ),
    .X(_194_));
 sky130_fd_sc_hd__a22o_1 _384_ (.A1(_061_),
    .A2(\history_s2[2] ),
    .B1(net74),
    .B2(_194_),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _385_ (.A0(\history_s0[2] ),
    .A1(\history_s1[2] ),
    .S(net74),
    .X(_195_));
 sky130_fd_sc_hd__mux2_1 _386_ (.A0(\history_s2[3] ),
    .A1(_195_),
    .S(net55),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _387_ (.A0(\history_s0[3] ),
    .A1(\history_s1[3] ),
    .S(net74),
    .X(_196_));
 sky130_fd_sc_hd__mux2_1 _388_ (.A0(\history_s2[4] ),
    .A1(_196_),
    .S(net50),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _389_ (.A0(\history_s0[4] ),
    .A1(\history_s1[4] ),
    .S(net74),
    .X(_197_));
 sky130_fd_sc_hd__mux2_1 _390_ (.A0(\history_s2[5] ),
    .A1(_197_),
    .S(net50),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _391_ (.A0(\history_s0[5] ),
    .A1(\history_s1[5] ),
    .S(net74),
    .X(_198_));
 sky130_fd_sc_hd__mux2_1 _392_ (.A0(\history_s2[6] ),
    .A1(_198_),
    .S(net50),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _393_ (.A0(\history_s0[6] ),
    .A1(\history_s1[6] ),
    .S(net74),
    .X(_199_));
 sky130_fd_sc_hd__mux2_1 _394_ (.A0(\history_s2[7] ),
    .A1(_199_),
    .S(net48),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _395_ (.A0(\history_s0[7] ),
    .A1(\history_s1[7] ),
    .S(net75),
    .X(_200_));
 sky130_fd_sc_hd__mux2_1 _396_ (.A0(\history_s2[8] ),
    .A1(_200_),
    .S(net46),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _397_ (.A0(\history_s0[8] ),
    .A1(\history_s1[8] ),
    .S(net75),
    .X(_201_));
 sky130_fd_sc_hd__mux2_1 _398_ (.A0(\history_s2[9] ),
    .A1(_201_),
    .S(net44),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _399_ (.A0(\history_s0[9] ),
    .A1(\history_s1[9] ),
    .S(net75),
    .X(_202_));
 sky130_fd_sc_hd__mux2_1 _400_ (.A0(\history_s2[10] ),
    .A1(_202_),
    .S(net44),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _401_ (.A0(\history_s0[10] ),
    .A1(\history_s1[10] ),
    .S(net75),
    .X(_203_));
 sky130_fd_sc_hd__mux2_1 _402_ (.A0(\history_s2[11] ),
    .A1(_203_),
    .S(net45),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _403_ (.A0(\history_s0[11] ),
    .A1(\history_s1[11] ),
    .S(net75),
    .X(_204_));
 sky130_fd_sc_hd__mux2_1 _404_ (.A0(\history_s2[12] ),
    .A1(_204_),
    .S(net46),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _405_ (.A0(\history_s0[12] ),
    .A1(\history_s1[12] ),
    .S(net3),
    .X(_205_));
 sky130_fd_sc_hd__mux2_1 _406_ (.A0(\history_s2[13] ),
    .A1(_205_),
    .S(net53),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _407_ (.A0(\history_s0[13] ),
    .A1(\history_s1[13] ),
    .S(net3),
    .X(_206_));
 sky130_fd_sc_hd__mux2_1 _408_ (.A0(\history_s2[14] ),
    .A1(_206_),
    .S(net53),
    .X(_015_));
 sky130_fd_sc_hd__a22o_1 _409_ (.A1(_061_),
    .A2(\history_s0[2] ),
    .B1(net81),
    .B2(_194_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _410_ (.A0(\history_s0[2] ),
    .A1(\history_s1[2] ),
    .S(net81),
    .X(_207_));
 sky130_fd_sc_hd__mux2_1 _411_ (.A0(\history_s0[3] ),
    .A1(_207_),
    .S(net55),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _412_ (.A0(\history_s0[3] ),
    .A1(\history_s1[3] ),
    .S(net81),
    .X(_208_));
 sky130_fd_sc_hd__mux2_1 _413_ (.A0(\history_s0[4] ),
    .A1(_208_),
    .S(net51),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _414_ (.A0(\history_s0[4] ),
    .A1(\history_s1[4] ),
    .S(net81),
    .X(_209_));
 sky130_fd_sc_hd__mux2_1 _415_ (.A0(\history_s0[5] ),
    .A1(_209_),
    .S(net50),
    .X(_019_));
 sky130_fd_sc_hd__mux2_1 _416_ (.A0(\history_s0[5] ),
    .A1(\history_s1[5] ),
    .S(net81),
    .X(_210_));
 sky130_fd_sc_hd__mux2_1 _417_ (.A0(\history_s0[6] ),
    .A1(_210_),
    .S(net50),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _418_ (.A0(\history_s0[6] ),
    .A1(\history_s1[6] ),
    .S(net81),
    .X(_211_));
 sky130_fd_sc_hd__mux2_1 _419_ (.A0(\history_s0[7] ),
    .A1(_211_),
    .S(net48),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _420_ (.A0(\history_s0[7] ),
    .A1(\history_s1[7] ),
    .S(net82),
    .X(_212_));
 sky130_fd_sc_hd__mux2_1 _421_ (.A0(\history_s0[8] ),
    .A1(_212_),
    .S(net46),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _422_ (.A0(\history_s0[8] ),
    .A1(\history_s1[8] ),
    .S(net82),
    .X(_213_));
 sky130_fd_sc_hd__mux2_1 _423_ (.A0(\history_s0[9] ),
    .A1(_213_),
    .S(net44),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _424_ (.A0(\history_s0[9] ),
    .A1(\history_s1[9] ),
    .S(net82),
    .X(_214_));
 sky130_fd_sc_hd__mux2_1 _425_ (.A0(\history_s0[10] ),
    .A1(_214_),
    .S(net45),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _426_ (.A0(\history_s0[10] ),
    .A1(\history_s1[10] ),
    .S(net82),
    .X(_215_));
 sky130_fd_sc_hd__mux2_1 _427_ (.A0(\history_s0[11] ),
    .A1(_215_),
    .S(net46),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _428_ (.A0(\history_s0[11] ),
    .A1(\history_s1[11] ),
    .S(net82),
    .X(_216_));
 sky130_fd_sc_hd__mux2_1 _429_ (.A0(\history_s0[12] ),
    .A1(_216_),
    .S(net48),
    .X(_026_));
 sky130_fd_sc_hd__mux2_1 _430_ (.A0(\history_s0[12] ),
    .A1(\history_s1[12] ),
    .S(net1),
    .X(_217_));
 sky130_fd_sc_hd__mux2_1 _431_ (.A0(\history_s0[13] ),
    .A1(_217_),
    .S(net53),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _432_ (.A0(\history_s0[13] ),
    .A1(\history_s1[13] ),
    .S(net1),
    .X(_218_));
 sky130_fd_sc_hd__mux2_1 _433_ (.A0(\history_s0[14] ),
    .A1(_218_),
    .S(net54),
    .X(_028_));
 sky130_fd_sc_hd__or2_1 _434_ (.A(net54),
    .B(\history_s2[0] ),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _435_ (.A0(\history_s1[1] ),
    .A1(\history_s2[0] ),
    .S(net54),
    .X(_030_));
 sky130_fd_sc_hd__a22o_1 _436_ (.A1(_061_),
    .A2(\history_s3[2] ),
    .B1(_194_),
    .B2(net41),
    .X(_031_));
 sky130_fd_sc_hd__mux2_1 _437_ (.A0(\history_s2[2] ),
    .A1(\history_s3[2] ),
    .S(net41),
    .X(_219_));
 sky130_fd_sc_hd__mux2_1 _438_ (.A0(\history_s3[3] ),
    .A1(_219_),
    .S(net53),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _439_ (.A0(\history_s2[3] ),
    .A1(\history_s3[3] ),
    .S(net42),
    .X(_220_));
 sky130_fd_sc_hd__mux2_1 _440_ (.A0(\history_s3[4] ),
    .A1(_220_),
    .S(net51),
    .X(_033_));
 sky130_fd_sc_hd__mux2_1 _441_ (.A0(\history_s2[4] ),
    .A1(\history_s3[4] ),
    .S(net41),
    .X(_221_));
 sky130_fd_sc_hd__mux2_1 _442_ (.A0(\history_s3[5] ),
    .A1(_221_),
    .S(net49),
    .X(_034_));
 sky130_fd_sc_hd__mux2_1 _443_ (.A0(\history_s2[5] ),
    .A1(\history_s3[5] ),
    .S(net41),
    .X(_222_));
 sky130_fd_sc_hd__mux2_1 _444_ (.A0(\history_s3[6] ),
    .A1(_222_),
    .S(net49),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _445_ (.A0(\history_s2[6] ),
    .A1(\history_s3[6] ),
    .S(net41),
    .X(_223_));
 sky130_fd_sc_hd__mux2_1 _446_ (.A0(\history_s3[7] ),
    .A1(_223_),
    .S(net48),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _447_ (.A0(\history_s2[7] ),
    .A1(\history_s3[7] ),
    .S(net41),
    .X(_224_));
 sky130_fd_sc_hd__mux2_1 _448_ (.A0(\history_s3[8] ),
    .A1(_224_),
    .S(net47),
    .X(_037_));
 sky130_fd_sc_hd__mux2_1 _449_ (.A0(\history_s2[8] ),
    .A1(\history_s3[8] ),
    .S(net43),
    .X(_225_));
 sky130_fd_sc_hd__mux2_1 _450_ (.A0(\history_s3[9] ),
    .A1(_225_),
    .S(net47),
    .X(_038_));
 sky130_fd_sc_hd__mux2_1 _451_ (.A0(\history_s2[9] ),
    .A1(\history_s3[9] ),
    .S(net43),
    .X(_226_));
 sky130_fd_sc_hd__mux2_1 _452_ (.A0(\history_s3[10] ),
    .A1(_226_),
    .S(net44),
    .X(_039_));
 sky130_fd_sc_hd__mux2_1 _453_ (.A0(\history_s2[10] ),
    .A1(\history_s3[10] ),
    .S(net43),
    .X(_227_));
 sky130_fd_sc_hd__mux2_1 _454_ (.A0(\history_s3[11] ),
    .A1(_227_),
    .S(net45),
    .X(_040_));
 sky130_fd_sc_hd__mux2_1 _455_ (.A0(\history_s2[11] ),
    .A1(\history_s3[11] ),
    .S(net43),
    .X(_228_));
 sky130_fd_sc_hd__mux2_1 _456_ (.A0(\history_s3[12] ),
    .A1(_228_),
    .S(net47),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _457_ (.A0(\history_s2[12] ),
    .A1(\history_s3[12] ),
    .S(net42),
    .X(_229_));
 sky130_fd_sc_hd__mux2_1 _458_ (.A0(\history_s3[13] ),
    .A1(_229_),
    .S(net47),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _459_ (.A0(\history_s2[13] ),
    .A1(\history_s3[13] ),
    .S(net42),
    .X(_230_));
 sky130_fd_sc_hd__mux2_1 _460_ (.A0(\history_s3[14] ),
    .A1(_230_),
    .S(net47),
    .X(_043_));
 sky130_fd_sc_hd__a22o_1 _461_ (.A1(_061_),
    .A2(\history_s1[2] ),
    .B1(net77),
    .B2(_194_),
    .X(_044_));
 sky130_fd_sc_hd__mux2_1 _462_ (.A0(\history_s2[2] ),
    .A1(\history_s3[2] ),
    .S(net77),
    .X(_231_));
 sky130_fd_sc_hd__mux2_1 _463_ (.A0(\history_s1[3] ),
    .A1(_231_),
    .S(net55),
    .X(_045_));
 sky130_fd_sc_hd__mux2_1 _464_ (.A0(\history_s2[3] ),
    .A1(\history_s3[3] ),
    .S(net78),
    .X(_232_));
 sky130_fd_sc_hd__mux2_1 _465_ (.A0(\history_s1[4] ),
    .A1(_232_),
    .S(net51),
    .X(_046_));
 sky130_fd_sc_hd__mux2_1 _466_ (.A0(\history_s2[4] ),
    .A1(\history_s3[4] ),
    .S(net77),
    .X(_233_));
 sky130_fd_sc_hd__mux2_1 _467_ (.A0(\history_s1[5] ),
    .A1(_233_),
    .S(net50),
    .X(_047_));
 sky130_fd_sc_hd__mux2_1 _468_ (.A0(\history_s2[5] ),
    .A1(\history_s3[5] ),
    .S(net77),
    .X(_234_));
 sky130_fd_sc_hd__mux2_1 _469_ (.A0(\history_s1[6] ),
    .A1(_234_),
    .S(net48),
    .X(_048_));
 sky130_fd_sc_hd__mux2_1 _470_ (.A0(\history_s2[6] ),
    .A1(\history_s3[6] ),
    .S(net77),
    .X(_235_));
 sky130_fd_sc_hd__mux2_1 _471_ (.A0(\history_s1[7] ),
    .A1(_235_),
    .S(net48),
    .X(_049_));
 sky130_fd_sc_hd__mux2_1 _472_ (.A0(\history_s2[7] ),
    .A1(\history_s3[7] ),
    .S(net77),
    .X(_236_));
 sky130_fd_sc_hd__mux2_1 _473_ (.A0(\history_s1[8] ),
    .A1(_236_),
    .S(net44),
    .X(_050_));
 sky130_fd_sc_hd__mux2_1 _474_ (.A0(\history_s2[8] ),
    .A1(\history_s3[8] ),
    .S(net79),
    .X(_237_));
 sky130_fd_sc_hd__mux2_1 _475_ (.A0(\history_s1[9] ),
    .A1(_237_),
    .S(net44),
    .X(_051_));
 sky130_fd_sc_hd__mux2_1 _476_ (.A0(\history_s2[9] ),
    .A1(\history_s3[9] ),
    .S(net79),
    .X(_238_));
 sky130_fd_sc_hd__mux2_1 _477_ (.A0(\history_s1[10] ),
    .A1(_238_),
    .S(net45),
    .X(_052_));
 sky130_fd_sc_hd__mux2_1 _478_ (.A0(\history_s2[10] ),
    .A1(\history_s3[10] ),
    .S(net79),
    .X(_239_));
 sky130_fd_sc_hd__mux2_1 _479_ (.A0(\history_s1[11] ),
    .A1(_239_),
    .S(net45),
    .X(_053_));
 sky130_fd_sc_hd__mux2_1 _480_ (.A0(\history_s2[11] ),
    .A1(\history_s3[11] ),
    .S(net79),
    .X(_240_));
 sky130_fd_sc_hd__mux2_1 _481_ (.A0(\history_s1[12] ),
    .A1(_240_),
    .S(net49),
    .X(_054_));
 sky130_fd_sc_hd__mux2_1 _482_ (.A0(\history_s2[12] ),
    .A1(\history_s3[12] ),
    .S(net78),
    .X(_241_));
 sky130_fd_sc_hd__mux2_1 _483_ (.A0(\history_s1[13] ),
    .A1(_241_),
    .S(net53),
    .X(_055_));
 sky130_fd_sc_hd__mux2_1 _484_ (.A0(\history_s2[13] ),
    .A1(\history_s3[13] ),
    .S(net78),
    .X(_242_));
 sky130_fd_sc_hd__mux2_1 _485_ (.A0(\history_s1[14] ),
    .A1(_242_),
    .S(net57),
    .X(_056_));
 sky130_fd_sc_hd__and3b_1 _486_ (.A_N(pipeline_full),
    .B(\latency_counter[0] ),
    .C(net56),
    .X(_243_));
 sky130_fd_sc_hd__o21ba_1 _487_ (.A1(_061_),
    .A2(pipeline_full),
    .B1_N(\latency_counter[0] ),
    .X(_244_));
 sky130_fd_sc_hd__nor2_1 _488_ (.A(_243_),
    .B(_244_),
    .Y(_057_));
 sky130_fd_sc_hd__xor2_1 _489_ (.A(\latency_counter[1] ),
    .B(_243_),
    .X(_058_));
 sky130_fd_sc_hd__and3_1 _490_ (.A(\latency_counter[1] ),
    .B(\latency_counter[2] ),
    .C(_243_),
    .X(_245_));
 sky130_fd_sc_hd__a21oi_1 _491_ (.A1(\latency_counter[1] ),
    .A2(_243_),
    .B1(\latency_counter[2] ),
    .Y(_246_));
 sky130_fd_sc_hd__nor2_1 _492_ (.A(_245_),
    .B(_246_),
    .Y(_059_));
 sky130_fd_sc_hd__xor2_1 _493_ (.A(\latency_counter[3] ),
    .B(_245_),
    .X(_060_));
 sky130_fd_sc_hd__dfrtp_1 _494_ (.CLK(clknet_3_7__leaf_clk),
    .D(_001_),
    .RESET_B(net69),
    .Q(pipeline_full));
 sky130_fd_sc_hd__dfrtp_1 _495_ (.CLK(clknet_3_7__leaf_clk),
    .D(_000_),
    .RESET_B(net69),
    .Q(net40));
 sky130_fd_sc_hd__dfrtp_1 _496_ (.CLK(clknet_3_6__leaf_clk),
    .D(_002_),
    .RESET_B(net67),
    .Q(net39));
 sky130_fd_sc_hd__dfrtp_1 _497_ (.CLK(clknet_3_6__leaf_clk),
    .D(_003_),
    .RESET_B(net67),
    .Q(\history_s2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _498_ (.CLK(clknet_3_5__leaf_clk),
    .D(_004_),
    .RESET_B(net64),
    .Q(\history_s2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _499_ (.CLK(clknet_3_5__leaf_clk),
    .D(_005_),
    .RESET_B(net65),
    .Q(\history_s2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _500_ (.CLK(clknet_3_5__leaf_clk),
    .D(_006_),
    .RESET_B(net64),
    .Q(\history_s2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _501_ (.CLK(clknet_3_5__leaf_clk),
    .D(_007_),
    .RESET_B(net64),
    .Q(\history_s2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _502_ (.CLK(clknet_3_4__leaf_clk),
    .D(_008_),
    .RESET_B(net62),
    .Q(\history_s2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _503_ (.CLK(clknet_3_1__leaf_clk),
    .D(_009_),
    .RESET_B(net60),
    .Q(\history_s2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _504_ (.CLK(clknet_3_0__leaf_clk),
    .D(_010_),
    .RESET_B(net58),
    .Q(\history_s2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _505_ (.CLK(clknet_3_0__leaf_clk),
    .D(_011_),
    .RESET_B(net58),
    .Q(\history_s2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _506_ (.CLK(clknet_3_2__leaf_clk),
    .D(_012_),
    .RESET_B(net59),
    .Q(\history_s2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _507_ (.CLK(clknet_3_3__leaf_clk),
    .D(_013_),
    .RESET_B(net60),
    .Q(\history_s2[12] ));
 sky130_fd_sc_hd__dfrtp_1 _508_ (.CLK(clknet_3_6__leaf_clk),
    .D(_014_),
    .RESET_B(net67),
    .Q(\history_s2[13] ));
 sky130_fd_sc_hd__dfrtp_1 _509_ (.CLK(clknet_3_6__leaf_clk),
    .D(_015_),
    .RESET_B(net68),
    .Q(\history_s2[14] ));
 sky130_fd_sc_hd__dfrtp_1 _510_ (.CLK(clknet_3_7__leaf_clk),
    .D(_016_),
    .RESET_B(net69),
    .Q(\history_s0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _511_ (.CLK(clknet_3_7__leaf_clk),
    .D(_017_),
    .RESET_B(net69),
    .Q(\history_s0[3] ));
 sky130_fd_sc_hd__dfrtp_1 _512_ (.CLK(clknet_3_5__leaf_clk),
    .D(_018_),
    .RESET_B(net65),
    .Q(\history_s0[4] ));
 sky130_fd_sc_hd__dfrtp_1 _513_ (.CLK(clknet_3_5__leaf_clk),
    .D(_019_),
    .RESET_B(net64),
    .Q(\history_s0[5] ));
 sky130_fd_sc_hd__dfrtp_1 _514_ (.CLK(clknet_3_4__leaf_clk),
    .D(_020_),
    .RESET_B(net64),
    .Q(\history_s0[6] ));
 sky130_fd_sc_hd__dfrtp_1 _515_ (.CLK(clknet_3_4__leaf_clk),
    .D(_021_),
    .RESET_B(net62),
    .Q(\history_s0[7] ));
 sky130_fd_sc_hd__dfrtp_1 _516_ (.CLK(clknet_3_1__leaf_clk),
    .D(_022_),
    .RESET_B(net60),
    .Q(\history_s0[8] ));
 sky130_fd_sc_hd__dfrtp_1 _517_ (.CLK(clknet_3_0__leaf_clk),
    .D(_023_),
    .RESET_B(net58),
    .Q(\history_s0[9] ));
 sky130_fd_sc_hd__dfrtp_1 _518_ (.CLK(clknet_3_0__leaf_clk),
    .D(_024_),
    .RESET_B(net58),
    .Q(\history_s0[10] ));
 sky130_fd_sc_hd__dfrtp_1 _519_ (.CLK(clknet_3_2__leaf_clk),
    .D(_025_),
    .RESET_B(net60),
    .Q(\history_s0[11] ));
 sky130_fd_sc_hd__dfrtp_1 _520_ (.CLK(clknet_3_1__leaf_clk),
    .D(_026_),
    .RESET_B(net62),
    .Q(\history_s0[12] ));
 sky130_fd_sc_hd__dfrtp_1 _521_ (.CLK(clknet_3_6__leaf_clk),
    .D(_027_),
    .RESET_B(net67),
    .Q(\history_s0[13] ));
 sky130_fd_sc_hd__dfrtp_1 _522_ (.CLK(clknet_3_6__leaf_clk),
    .D(_028_),
    .RESET_B(net68),
    .Q(\history_s0[14] ));
 sky130_fd_sc_hd__dfrtp_1 _523_ (.CLK(clknet_3_6__leaf_clk),
    .D(_029_),
    .RESET_B(net68),
    .Q(\history_s2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _524_ (.CLK(clknet_3_6__leaf_clk),
    .D(_030_),
    .RESET_B(net68),
    .Q(\history_s1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _525_ (.CLK(clknet_3_6__leaf_clk),
    .D(_031_),
    .RESET_B(net67),
    .Q(\history_s3[2] ));
 sky130_fd_sc_hd__dfrtp_1 _526_ (.CLK(clknet_3_4__leaf_clk),
    .D(_032_),
    .RESET_B(net63),
    .Q(\history_s3[3] ));
 sky130_fd_sc_hd__dfrtp_1 _527_ (.CLK(clknet_3_4__leaf_clk),
    .D(_033_),
    .RESET_B(net63),
    .Q(\history_s3[4] ));
 sky130_fd_sc_hd__dfrtp_1 _528_ (.CLK(clknet_3_5__leaf_clk),
    .D(_034_),
    .RESET_B(net63),
    .Q(\history_s3[5] ));
 sky130_fd_sc_hd__dfrtp_1 _529_ (.CLK(clknet_3_4__leaf_clk),
    .D(_035_),
    .RESET_B(net63),
    .Q(\history_s3[6] ));
 sky130_fd_sc_hd__dfrtp_1 _530_ (.CLK(clknet_3_1__leaf_clk),
    .D(_036_),
    .RESET_B(net62),
    .Q(\history_s3[7] ));
 sky130_fd_sc_hd__dfrtp_1 _531_ (.CLK(clknet_3_1__leaf_clk),
    .D(_037_),
    .RESET_B(net60),
    .Q(\history_s3[8] ));
 sky130_fd_sc_hd__dfrtp_1 _532_ (.CLK(clknet_3_1__leaf_clk),
    .D(_038_),
    .RESET_B(net61),
    .Q(\history_s3[9] ));
 sky130_fd_sc_hd__dfrtp_1 _533_ (.CLK(clknet_3_0__leaf_clk),
    .D(_039_),
    .RESET_B(net58),
    .Q(\history_s3[10] ));
 sky130_fd_sc_hd__dfrtp_1 _534_ (.CLK(clknet_3_2__leaf_clk),
    .D(_040_),
    .RESET_B(net59),
    .Q(\history_s3[11] ));
 sky130_fd_sc_hd__dfrtp_1 _535_ (.CLK(clknet_3_2__leaf_clk),
    .D(_041_),
    .RESET_B(net61),
    .Q(\history_s3[12] ));
 sky130_fd_sc_hd__dfrtp_1 _536_ (.CLK(clknet_3_3__leaf_clk),
    .D(_042_),
    .RESET_B(net61),
    .Q(\history_s3[13] ));
 sky130_fd_sc_hd__dfrtp_1 _537_ (.CLK(clknet_3_3__leaf_clk),
    .D(_043_),
    .RESET_B(net61),
    .Q(\history_s3[14] ));
 sky130_fd_sc_hd__dfrtp_1 _538_ (.CLK(clknet_3_7__leaf_clk),
    .D(_044_),
    .RESET_B(net69),
    .Q(\history_s1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _539_ (.CLK(clknet_3_5__leaf_clk),
    .D(_045_),
    .RESET_B(net69),
    .Q(\history_s1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _540_ (.CLK(clknet_3_5__leaf_clk),
    .D(_046_),
    .RESET_B(net65),
    .Q(\history_s1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _541_ (.CLK(clknet_3_5__leaf_clk),
    .D(_047_),
    .RESET_B(net64),
    .Q(\history_s1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _542_ (.CLK(clknet_3_4__leaf_clk),
    .D(_048_),
    .RESET_B(net62),
    .Q(\history_s1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _543_ (.CLK(clknet_3_1__leaf_clk),
    .D(_049_),
    .RESET_B(net62),
    .Q(\history_s1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _544_ (.CLK(clknet_3_0__leaf_clk),
    .D(_050_),
    .RESET_B(net59),
    .Q(\history_s1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _545_ (.CLK(clknet_3_0__leaf_clk),
    .D(_051_),
    .RESET_B(net58),
    .Q(\history_s1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _546_ (.CLK(clknet_3_0__leaf_clk),
    .D(_052_),
    .RESET_B(net59),
    .Q(\history_s1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _547_ (.CLK(clknet_3_0__leaf_clk),
    .D(_053_),
    .RESET_B(net59),
    .Q(\history_s1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _548_ (.CLK(clknet_3_3__leaf_clk),
    .D(_054_),
    .RESET_B(net63),
    .Q(\history_s1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _549_ (.CLK(clknet_3_6__leaf_clk),
    .D(_055_),
    .RESET_B(net67),
    .Q(\history_s1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _550_ (.CLK(clknet_3_3__leaf_clk),
    .D(_056_),
    .RESET_B(net61),
    .Q(\history_s1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _551_ (.CLK(clknet_3_7__leaf_clk),
    .D(_057_),
    .RESET_B(net70),
    .Q(\latency_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _552_ (.CLK(clknet_3_7__leaf_clk),
    .D(_058_),
    .RESET_B(net70),
    .Q(\latency_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _553_ (.CLK(clknet_3_7__leaf_clk),
    .D(_059_),
    .RESET_B(net70),
    .Q(\latency_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _554_ (.CLK(clknet_3_7__leaf_clk),
    .D(_060_),
    .RESET_B(net70),
    .Q(\latency_counter[3] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_338 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(dec_bits_i[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(dec_bits_i[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(dec_bits_i[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(dec_bits_i[3]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(pm_new_s0_i[0]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(pm_new_s0_i[1]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(pm_new_s0_i[2]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(pm_new_s0_i[3]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(pm_new_s0_i[4]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(pm_new_s0_i[5]),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(pm_new_s0_i[6]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(pm_new_s0_i[7]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(pm_new_s1_i[0]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(pm_new_s1_i[1]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(pm_new_s1_i[2]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(pm_new_s1_i[3]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(pm_new_s1_i[4]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(pm_new_s1_i[5]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(pm_new_s1_i[6]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(pm_new_s1_i[7]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(pm_new_s2_i[0]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(pm_new_s2_i[1]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(pm_new_s2_i[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(pm_new_s2_i[3]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(pm_new_s2_i[4]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(pm_new_s2_i[5]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(pm_new_s2_i[6]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(pm_new_s2_i[7]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(pm_new_s3_i[0]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(pm_new_s3_i[1]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(pm_new_s3_i[2]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(pm_new_s3_i[3]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(pm_new_s3_i[4]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(pm_new_s3_i[5]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(pm_new_s3_i[6]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(pm_new_s3_i[7]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(rst_n),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(valid_i),
    .X(net38));
 sky130_fd_sc_hd__buf_4 output39 (.A(net39),
    .X(decoded_bit_o));
 sky130_fd_sc_hd__buf_4 output40 (.A(net40),
    .X(valid_o));
 sky130_fd_sc_hd__clkbuf_2 fanout41 (.A(net43),
    .X(net41));
 sky130_fd_sc_hd__buf_1 fanout42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(net4),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 fanout44 (.A(net46),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__buf_2 fanout46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__buf_2 fanout47 (.A(net57),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 fanout48 (.A(net52),
    .X(net48));
 sky130_fd_sc_hd__buf_1 fanout49 (.A(net52),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 fanout50 (.A(net52),
    .X(net50));
 sky130_fd_sc_hd__buf_1 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__buf_1 fanout52 (.A(net57),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 fanout53 (.A(net56),
    .X(net53));
 sky130_fd_sc_hd__buf_1 fanout54 (.A(net56),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout56 (.A(net57),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 fanout57 (.A(net38),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 fanout58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__buf_2 fanout59 (.A(net60),
    .X(net59));
 sky130_fd_sc_hd__buf_2 fanout60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__buf_2 fanout61 (.A(net72),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 fanout62 (.A(net66),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 fanout63 (.A(net66),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 fanout64 (.A(net66),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 fanout65 (.A(net66),
    .X(net65));
 sky130_fd_sc_hd__buf_1 fanout66 (.A(net72),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 fanout67 (.A(net71),
    .X(net67));
 sky130_fd_sc_hd__buf_1 fanout68 (.A(net71),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 fanout69 (.A(net71),
    .X(net69));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout71 (.A(net72),
    .X(net71));
 sky130_fd_sc_hd__buf_1 fanout72 (.A(net37),
    .X(net72));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout73 (.A(net34),
    .X(net73));
 sky130_fd_sc_hd__buf_2 fanout74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__buf_2 fanout75 (.A(net3),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 fanout76 (.A(net24),
    .X(net76));
 sky130_fd_sc_hd__buf_2 fanout77 (.A(net79),
    .X(net77));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__buf_2 fanout79 (.A(net2),
    .X(net79));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout80 (.A(net16),
    .X(net80));
 sky130_fd_sc_hd__buf_2 fanout81 (.A(net82),
    .X(net81));
 sky130_fd_sc_hd__buf_2 fanout82 (.A(net1),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload0 (.A(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload1 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload2 (.A(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload3 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload4 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload5 (.A(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(dec_bits_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(dec_bits_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(dec_bits_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(dec_bits_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(pm_new_s0_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(pm_new_s0_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(pm_new_s0_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(pm_new_s0_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(pm_new_s0_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(pm_new_s0_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(pm_new_s0_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(pm_new_s0_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(pm_new_s1_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(pm_new_s1_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(pm_new_s1_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(pm_new_s1_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(pm_new_s1_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(pm_new_s1_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(pm_new_s1_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(pm_new_s1_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(pm_new_s2_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(pm_new_s2_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(pm_new_s2_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(pm_new_s2_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(pm_new_s2_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(pm_new_s2_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(pm_new_s2_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(pm_new_s2_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(pm_new_s3_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(pm_new_s3_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(pm_new_s3_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(pm_new_s3_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(pm_new_s3_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(pm_new_s3_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(pm_new_s3_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(pm_new_s3_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(rst_n));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(valid_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__432__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__430__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_X (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__407__S (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__405__S (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__496__Q (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__382__A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_X (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__460__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__458__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__456__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__448__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__450__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout46_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_X (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__485__S (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_X (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__550__RESET_B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__537__RESET_B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__536__RESET_B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__535__RESET_B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__532__RESET_B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_X (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_X (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__403__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__401__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__399__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__397__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__395__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__480__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__478__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__476__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__474__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__428__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__426__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__424__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__422__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__420__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_293 ();
endmodule
