* NGSPICE file created from piso.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

.subckt piso clk data_serial_o[0] data_serial_o[1] fifo_data_i[0] fifo_data_i[10]
+ fifo_data_i[11] fifo_data_i[12] fifo_data_i[13] fifo_data_i[14] fifo_data_i[15]
+ fifo_data_i[1] fifo_data_i[2] fifo_data_i[3] fifo_data_i[4] fifo_data_i[5] fifo_data_i[6]
+ fifo_data_i[7] fifo_data_i[8] fifo_data_i[9] fifo_empty_i fifo_rd_en_o rst_n valid_serial_o
+ vccd1 vssd1
X_062_ _023_ net25 count\[3\] vssd1 vssd1 vccd1 vccd1 _042_ sky130_fd_sc_hd__and3b_1
XFILLER_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_114_ clknet_1_1__leaf_clk _038_ net41 vssd1 vssd1 vccd1 vccd1 state\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_6_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_45 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input18_A rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 data_serial_o[1] sky130_fd_sc_hd__buf_4
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_55 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_061_ count\[3\] _023_ net25 _027_ net32 vssd1 vssd1 vccd1 vccd1 _041_ sky130_fd_sc_hd__a311o_1
X_113_ clknet_1_0__leaf_clk _042_ net40 vssd1 vssd1 vccd1 vccd1 count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 fifo_rd_en_o sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_56 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_060_ _022_ net25 count\[2\] vssd1 vssd1 vccd1 vccd1 _027_ sky130_fd_sc_hd__and3b_1
X_112_ clknet_1_0__leaf_clk _041_ net40 vssd1 vssd1 vccd1 vccd1 count\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_6_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 valid_serial_o sky130_fd_sc_hd__buf_4
XFILLER_15_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_111_ clknet_1_1__leaf_clk _040_ net40 vssd1 vssd1 vccd1 vccd1 count\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input16_A fifo_data_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input8_A fifo_data_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_110_ clknet_1_0__leaf_clk _039_ net40 vssd1 vssd1 vccd1 vccd1 count\[0\] sky130_fd_sc_hd__dfrtp_1
Xclkload0 clknet_1_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload0/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_49 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_099_ clknet_1_1__leaf_clk _007_ net39 vssd1 vssd1 vccd1 vccd1 shift_reg\[9\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_3_Left_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input6_A fifo_data_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_A fifo_data_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_098_ clknet_1_0__leaf_clk _006_ net39 vssd1 vssd1 vccd1 vccd1 shift_reg\[8\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_7_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_51 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_097_ clknet_1_0__leaf_clk _005_ net38 vssd1 vssd1 vccd1 vccd1 shift_reg\[7\] sky130_fd_sc_hd__dfrtp_1
Xfanout40 net42 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_2
XFILLER_16_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_61 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_42 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout41 net42 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout30 net31 vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_1
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_52 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Left_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_096_ clknet_1_0__leaf_clk _004_ net38 vssd1 vssd1 vccd1 vccd1 shift_reg\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_1_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_62 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_079_ shift_reg\[8\] net27 net23 net15 net37 vssd1 vssd1 vccd1 vccd1 _034_ sky130_fd_sc_hd__a32o_1
XFILLER_7_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input12_A fifo_data_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input4_A fifo_data_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout31 _024_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_1
Xfanout42 net18 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_2
X_095_ clknet_1_0__leaf_clk _003_ net38 vssd1 vssd1 vccd1 vccd1 shift_reg\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_53 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_078_ shift_reg\[9\] _033_ net34 vssd1 vssd1 vccd1 vccd1 _007_ sky130_fd_sc_hd__mux2_1
Xoutput19 net19 vssd1 vssd1 vccd1 vccd1 data_serial_o[0] sky130_fd_sc_hd__buf_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout32 _021_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_2
X_094_ clknet_1_0__leaf_clk _002_ net38 vssd1 vssd1 vccd1 vccd1 shift_reg\[4\] sky130_fd_sc_hd__dfrtp_1
X_077_ shift_reg\[7\] net27 net23 net14 net36 vssd1 vssd1 vccd1 vccd1 _033_ sky130_fd_sc_hd__a32o_1
XFILLER_4_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout33 _021_ vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_1
XFILLER_13_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_093_ clknet_1_0__leaf_clk _001_ net38 vssd1 vssd1 vccd1 vccd1 shift_reg\[3\] sky130_fd_sc_hd__dfrtp_1
X_076_ shift_reg\[8\] _032_ net35 vssd1 vssd1 vccd1 vccd1 _006_ sky130_fd_sc_hd__mux2_1
XFILLER_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput1 fifo_data_i[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_059_ net32 _022_ _026_ _038_ vssd1 vssd1 vccd1 vccd1 _040_ sky130_fd_sc_hd__o31a_1
XFILLER_7_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout34 net35 vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout23 net24 vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_0_36 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input10_A fifo_data_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput2 fifo_data_i[10] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input2_A fifo_data_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_092_ clknet_1_0__leaf_clk _000_ net38 vssd1 vssd1 vccd1 vccd1 shift_reg\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_075_ shift_reg\[6\] net28 net24 net13 net36 vssd1 vssd1 vccd1 vccd1 _032_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_6_46 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_058_ count\[0\] count\[1\] vssd1 vssd1 vccd1 vccd1 _026_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_14_Left_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout35 _020_ vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout24 net26 vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_0_37 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_091_ net30 net25 net33 vssd1 vssd1 vccd1 vccd1 _045_ sky130_fd_sc_hd__a21o_1
Xinput3 fifo_data_i[11] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_47 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_074_ shift_reg\[7\] _031_ net35 vssd1 vssd1 vccd1 vccd1 _005_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_2_Left_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_057_ _018_ net28 net25 net32 vssd1 vssd1 vccd1 vccd1 _039_ sky130_fd_sc_hd__a31o_1
X_109_ clknet_1_1__leaf_clk _045_ net41 vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__dfrtp_1
Xfanout25 net26 vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_13_57 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout36 _017_ vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_0_38 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_090_ shift_reg\[15\] _016_ net34 vssd1 vssd1 vccd1 vccd1 _013_ sky130_fd_sc_hd__mux2_1
Xinput4 fifo_data_i[12] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_056_ net30 net26 net33 vssd1 vssd1 vccd1 vccd1 _038_ sky130_fd_sc_hd__a21o_1
XFILLER_10_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_073_ shift_reg\[5\] net27 net23 net12 net36 vssd1 vssd1 vccd1 vccd1 _031_ sky130_fd_sc_hd__a32o_1
X_108_ clknet_1_1__leaf_clk _044_ net41 vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__dfrtp_1
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout37 _017_ vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_2
Xfanout26 _025_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_1
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 fifo_data_i[13] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_072_ shift_reg\[6\] _030_ net35 vssd1 vssd1 vccd1 vccd1 _004_ sky130_fd_sc_hd__mux2_1
X_055_ net21 state\[1\] vssd1 vssd1 vccd1 vccd1 _025_ sky130_fd_sc_hd__and2b_1
X_107_ clknet_1_0__leaf_clk _043_ net40 vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__dfrtp_1
Xfanout38 net39 vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_2
Xfanout27 net28 vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput6 fifo_data_i[14] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_071_ shift_reg\[4\] net27 net23 net11 net36 vssd1 vssd1 vccd1 vccd1 _030_ sky130_fd_sc_hd__a32o_1
XFILLER_2_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_106_ clknet_1_1__leaf_clk _037_ net42 vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__dfrtp_1
XFILLER_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_054_ count\[2\] count\[3\] count\[0\] count\[1\] vssd1 vssd1 vccd1 vccd1 _024_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout39 net42 vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout28 net31 vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_1
Xinput7 fifo_data_i[15] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
X_070_ shift_reg\[5\] _029_ net35 vssd1 vssd1 vccd1 vccd1 _003_ sky130_fd_sc_hd__mux2_1
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_053_ count\[2\] _022_ vssd1 vssd1 vccd1 vccd1 _023_ sky130_fd_sc_hd__and2b_1
XFILLER_2_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput10 fifo_data_i[3] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_105_ clknet_1_1__leaf_clk _013_ net42 vssd1 vssd1 vccd1 vccd1 shift_reg\[15\] sky130_fd_sc_hd__dfrtp_1
Xfanout29 net31 vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput8 fifo_data_i[1] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
X_104_ clknet_1_1__leaf_clk _012_ net41 vssd1 vssd1 vccd1 vccd1 shift_reg\[14\] sky130_fd_sc_hd__dfrtp_1
X_052_ count\[0\] count\[1\] vssd1 vssd1 vccd1 vccd1 _022_ sky130_fd_sc_hd__nor2_1
Xinput11 fifo_data_i[4] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_input17_A fifo_empty_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input9_A fifo_data_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput9 fifo_data_i[2] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
X_051_ state\[1\] net21 vssd1 vssd1 vccd1 vccd1 _021_ sky130_fd_sc_hd__and2b_1
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput12 fifo_data_i[5] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_103_ clknet_1_1__leaf_clk _011_ net39 vssd1 vssd1 vccd1 vccd1 shift_reg\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_050_ net17 net34 vssd1 vssd1 vccd1 vccd1 _037_ sky130_fd_sc_hd__nor2_1
X_102_ clknet_1_1__leaf_clk _010_ net40 vssd1 vssd1 vccd1 vccd1 shift_reg\[12\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Left_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput13 fifo_data_i[6] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_13_Left_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_43 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput14 fifo_data_i[7] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_17_63 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_101_ clknet_1_1__leaf_clk _009_ net39 vssd1 vssd1 vccd1 vccd1 shift_reg\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input15_A fifo_data_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_44 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input7_A fifo_data_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_54 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_100_ clknet_1_1__leaf_clk _008_ net39 vssd1 vssd1 vccd1 vccd1 shift_reg\[10\] sky130_fd_sc_hd__dfrtp_1
Xinput15 fifo_data_i[8] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_17_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_64 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_65 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput16 fifo_data_i[9] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput17 fifo_empty_i vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_089_ shift_reg\[13\] net29 net26 net5 net37 vssd1 vssd1 vccd1 vccd1 _016_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_5_Left_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_input13_A fifo_data_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input5_A fifo_data_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_088_ shift_reg\[14\] _015_ _020_ vssd1 vssd1 vccd1 vccd1 _012_ sky130_fd_sc_hd__mux2_1
XFILLER_8_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput18 rst_n vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_48 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_087_ shift_reg\[12\] net29 net26 net4 net37 vssd1 vssd1 vccd1 vccd1 _015_ sky130_fd_sc_hd__a32o_1
XFILLER_11_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_58 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_39 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_086_ shift_reg\[13\] _014_ net34 vssd1 vssd1 vccd1 vccd1 _011_ sky130_fd_sc_hd__mux2_1
XFILLER_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Left_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_069_ shift_reg\[3\] net27 net23 net10 net36 vssd1 vssd1 vccd1 vccd1 _029_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_14_59 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input3_A fifo_data_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A fifo_data_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_085_ shift_reg\[11\] net29 net24 net3 net37 vssd1 vssd1 vccd1 vccd1 _014_ sky130_fd_sc_hd__a32o_1
X_068_ shift_reg\[4\] _028_ net35 vssd1 vssd1 vccd1 vccd1 _002_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_12_Left_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_40 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_084_ shift_reg\[12\] _036_ _020_ vssd1 vssd1 vccd1 vccd1 _010_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_50 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_067_ shift_reg\[2\] net27 net23 net9 net36 vssd1 vssd1 vccd1 vccd1 _028_ sky130_fd_sc_hd__a32o_1
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_60 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_41 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_083_ shift_reg\[10\] net29 net24 net2 net37 vssd1 vssd1 vccd1 vccd1 _036_ sky130_fd_sc_hd__a32o_1
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_049_ net21 state\[1\] vssd1 vssd1 vccd1 vccd1 _020_ sky130_fd_sc_hd__or2_1
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_066_ shift_reg\[3\] _019_ net32 net8 vssd1 vssd1 vccd1 vccd1 _001_ sky130_fd_sc_hd__a22o_1
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_082_ shift_reg\[11\] _035_ net34 vssd1 vssd1 vccd1 vccd1 _009_ sky130_fd_sc_hd__mux2_1
XANTENNA_input1_A fifo_data_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_065_ shift_reg\[2\] _019_ net32 net1 vssd1 vssd1 vccd1 vccd1 _000_ sky130_fd_sc_hd__a22o_1
X_048_ net21 state\[1\] vssd1 vssd1 vccd1 vccd1 _019_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_16_Left_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Left_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_081_ shift_reg\[9\] net29 net24 net16 net37 vssd1 vssd1 vccd1 vccd1 _035_ sky130_fd_sc_hd__a32o_1
XFILLER_6_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_064_ shift_reg\[15\] net30 net24 net7 net33 vssd1 vssd1 vccd1 vccd1 _044_ sky130_fd_sc_hd__a32o_1
XFILLER_9_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Left_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_047_ count\[0\] vssd1 vssd1 vccd1 vccd1 _018_ sky130_fd_sc_hd__inv_2
X_063_ shift_reg\[14\] net29 net25 net6 net32 vssd1 vssd1 vccd1 vccd1 _043_ sky130_fd_sc_hd__a32o_1
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_080_ shift_reg\[10\] _034_ net34 vssd1 vssd1 vccd1 vccd1 _008_ sky130_fd_sc_hd__mux2_1
X_046_ state\[1\] vssd1 vssd1 vccd1 vccd1 _017_ sky130_fd_sc_hd__inv_2
XFILLER_9_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
.ends

