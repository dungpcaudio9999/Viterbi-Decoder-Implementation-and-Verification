// bmu.v - Block Metric Unit
// T�nh to�n Chi ph� Hamming (Branch Metric)
module bmu (
    input  [1:0] piso_data_i,    // D? li?u nh?n ???c (2 bits)
    
    // ??u ra Chi ph� Hamming (2 bits)
    output [1:0] bm_s0_s0_o,
    output [1:0] bm_s0_s2_o,
    output [1:0] bm_s1_s0_o,
    output [1:0] bm_s1_s2_o,
    output [1:0] bm_s2_s1_o,
    output [1:0] bm_s2_s3_o,
    output [1:0] bm_s3_s1_o,
    output [1:0] bm_s3_s3_o
);

// --- Khai b�o Codeword D? ki?n (Expected Codewords) ---
parameter C00 = 2'b00; // Expected Codeword cho S0 -> S0
parameter C02 = 2'b11; // Expected Codeword cho S0 -> S2
parameter C10 = 2'b11; // Expected Codeword cho S1 -> S0
parameter C12 = 2'b00; // Expected Codeword cho S1 -> S2
parameter C21 = 2'b10; // Expected Codeword cho S2 -> S1
parameter C23 = 2'b01; // Expected Codeword cho S2 -> S3
parameter C31 = 2'b01; // Expected Codeword cho S3 -> S1
parameter C33 = 2'b10; // Expected Codeword cho S3 -> S3

// --- Khai b�o wire trung gian cho k?t qu? XOR (Hamming Distance) ---
// M?i wire c� ?? r?ng 2 bit
wire [1:0] diff_s0_s0 = piso_data_i ^ C00;
wire [1:0] diff_s0_s2 = piso_data_i ^ C02;
wire [1:0] diff_s1_s0 = piso_data_i ^ C10;
wire [1:0] diff_s1_s2 = piso_data_i ^ C12;
wire [1:0] diff_s2_s1 = piso_data_i ^ C21;
wire [1:0] diff_s2_s3 = piso_data_i ^ C23;
wire [1:0] diff_s3_s1 = piso_data_i ^ C31;
wire [1:0] diff_s3_s3 = piso_data_i ^ C33;

// --- H�m t�nh to�n Chi ph� Hamming (Hamming Weight) ---
// S? d?ng ph�p c?ng c�c bit ??n, nh?ng v?i bi?n trung gian, gi�p tr�nh bi�n d?ch x? l� d? h?n.

assign bm_s0_s0_o = diff_s0_s0[1] + diff_s0_s0[0];
assign bm_s0_s2_o = diff_s0_s2[1] + diff_s0_s2[0];

assign bm_s1_s0_o = diff_s1_s0[1] + diff_s1_s0[0];
assign bm_s1_s2_o = diff_s1_s2[1] + diff_s1_s2[0];

assign bm_s2_s1_o = diff_s2_s1[1] + diff_s2_s1[0];
assign bm_s2_s3_o = diff_s2_s3[1] + diff_s2_s3[0];

assign bm_s3_s1_o = diff_s3_s1[1] + diff_s3_s1[0];
assign bm_s3_s3_o = diff_s3_s3[1] + diff_s3_s3[0];

endmodule