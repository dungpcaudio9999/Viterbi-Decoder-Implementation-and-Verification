module sync_fifo (clk,
    empty_o,
    full_o,
    rd_en_i,
    rst_n,
    wr_en_i,
    rd_data_o,
    wr_data_i);
 input clk;
 output empty_o;
 output full_o;
 input rd_en_i;
 input rst_n;
 input wr_en_i;
 output [15:0] rd_data_o;
 input [15:0] wr_data_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire \count[0] ;
 wire \count[1] ;
 wire \count[2] ;
 wire \count[3] ;
 wire \count[4] ;
 wire \mem[0][0] ;
 wire \mem[0][10] ;
 wire \mem[0][11] ;
 wire \mem[0][12] ;
 wire \mem[0][13] ;
 wire \mem[0][14] ;
 wire \mem[0][15] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[0][8] ;
 wire \mem[0][9] ;
 wire \mem[10][0] ;
 wire \mem[10][10] ;
 wire \mem[10][11] ;
 wire \mem[10][12] ;
 wire \mem[10][13] ;
 wire \mem[10][14] ;
 wire \mem[10][15] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[10][8] ;
 wire \mem[10][9] ;
 wire \mem[11][0] ;
 wire \mem[11][10] ;
 wire \mem[11][11] ;
 wire \mem[11][12] ;
 wire \mem[11][13] ;
 wire \mem[11][14] ;
 wire \mem[11][15] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[11][8] ;
 wire \mem[11][9] ;
 wire \mem[12][0] ;
 wire \mem[12][10] ;
 wire \mem[12][11] ;
 wire \mem[12][12] ;
 wire \mem[12][13] ;
 wire \mem[12][14] ;
 wire \mem[12][15] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[12][8] ;
 wire \mem[12][9] ;
 wire \mem[13][0] ;
 wire \mem[13][10] ;
 wire \mem[13][11] ;
 wire \mem[13][12] ;
 wire \mem[13][13] ;
 wire \mem[13][14] ;
 wire \mem[13][15] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[13][8] ;
 wire \mem[13][9] ;
 wire \mem[14][0] ;
 wire \mem[14][10] ;
 wire \mem[14][11] ;
 wire \mem[14][12] ;
 wire \mem[14][13] ;
 wire \mem[14][14] ;
 wire \mem[14][15] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[14][8] ;
 wire \mem[14][9] ;
 wire \mem[15][0] ;
 wire \mem[15][10] ;
 wire \mem[15][11] ;
 wire \mem[15][12] ;
 wire \mem[15][13] ;
 wire \mem[15][14] ;
 wire \mem[15][15] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[15][8] ;
 wire \mem[15][9] ;
 wire \mem[1][0] ;
 wire \mem[1][10] ;
 wire \mem[1][11] ;
 wire \mem[1][12] ;
 wire \mem[1][13] ;
 wire \mem[1][14] ;
 wire \mem[1][15] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[1][8] ;
 wire \mem[1][9] ;
 wire \mem[2][0] ;
 wire \mem[2][10] ;
 wire \mem[2][11] ;
 wire \mem[2][12] ;
 wire \mem[2][13] ;
 wire \mem[2][14] ;
 wire \mem[2][15] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[2][8] ;
 wire \mem[2][9] ;
 wire \mem[3][0] ;
 wire \mem[3][10] ;
 wire \mem[3][11] ;
 wire \mem[3][12] ;
 wire \mem[3][13] ;
 wire \mem[3][14] ;
 wire \mem[3][15] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[3][8] ;
 wire \mem[3][9] ;
 wire \mem[4][0] ;
 wire \mem[4][10] ;
 wire \mem[4][11] ;
 wire \mem[4][12] ;
 wire \mem[4][13] ;
 wire \mem[4][14] ;
 wire \mem[4][15] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[4][8] ;
 wire \mem[4][9] ;
 wire \mem[5][0] ;
 wire \mem[5][10] ;
 wire \mem[5][11] ;
 wire \mem[5][12] ;
 wire \mem[5][13] ;
 wire \mem[5][14] ;
 wire \mem[5][15] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[5][8] ;
 wire \mem[5][9] ;
 wire \mem[6][0] ;
 wire \mem[6][10] ;
 wire \mem[6][11] ;
 wire \mem[6][12] ;
 wire \mem[6][13] ;
 wire \mem[6][14] ;
 wire \mem[6][15] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[6][8] ;
 wire \mem[6][9] ;
 wire \mem[7][0] ;
 wire \mem[7][10] ;
 wire \mem[7][11] ;
 wire \mem[7][12] ;
 wire \mem[7][13] ;
 wire \mem[7][14] ;
 wire \mem[7][15] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[7][8] ;
 wire \mem[7][9] ;
 wire \mem[8][0] ;
 wire \mem[8][10] ;
 wire \mem[8][11] ;
 wire \mem[8][12] ;
 wire \mem[8][13] ;
 wire \mem[8][14] ;
 wire \mem[8][15] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[8][8] ;
 wire \mem[8][9] ;
 wire \mem[9][0] ;
 wire \mem[9][10] ;
 wire \mem[9][11] ;
 wire \mem[9][12] ;
 wire \mem[9][13] ;
 wire \mem[9][14] ;
 wire \mem[9][15] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \mem[9][8] ;
 wire \mem[9][9] ;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sky130_fd_sc_hd__inv_2 _0519_ (.A(\count[4] ),
    .Y(_0292_));
 sky130_fd_sc_hd__inv_2 _0520_ (.A(\wr_ptr[3] ),
    .Y(_0293_));
 sky130_fd_sc_hd__inv_2 _0521_ (.A(net166),
    .Y(_0294_));
 sky130_fd_sc_hd__or4_2 _0522_ (.A(\count[1] ),
    .B(\count[0] ),
    .C(\count[3] ),
    .D(\count[2] ),
    .X(_0295_));
 sky130_fd_sc_hd__nor2_1 _0523_ (.A(\count[4] ),
    .B(_0295_),
    .Y(net20));
 sky130_fd_sc_hd__nor2_1 _0524_ (.A(_0292_),
    .B(_0295_),
    .Y(net21));
 sky130_fd_sc_hd__o21a_1 _0525_ (.A1(\count[4] ),
    .A2(_0295_),
    .B1(net1),
    .X(_0296_));
 sky130_fd_sc_hd__o21ai_1 _0526_ (.A1(\count[4] ),
    .A2(_0295_),
    .B1(net1),
    .Y(_0297_));
 sky130_fd_sc_hd__o21a_2 _0527_ (.A1(_0292_),
    .A2(_0295_),
    .B1(net19),
    .X(_0298_));
 sky130_fd_sc_hd__o21ai_1 _0528_ (.A1(_0292_),
    .A2(_0295_),
    .B1(net19),
    .Y(_0299_));
 sky130_fd_sc_hd__nor2_2 _0529_ (.A(net121),
    .B(_0298_),
    .Y(_0300_));
 sky130_fd_sc_hd__nor2_1 _0530_ (.A(net126),
    .B(net120),
    .Y(_0301_));
 sky130_fd_sc_hd__or2_2 _0531_ (.A(_0300_),
    .B(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__xor2_1 _0532_ (.A(\count[0] ),
    .B(_0302_),
    .X(_0000_));
 sky130_fd_sc_hd__a21o_1 _0533_ (.A1(net126),
    .A2(net120),
    .B1(\count[1] ),
    .X(_0303_));
 sky130_fd_sc_hd__and3_1 _0534_ (.A(\count[1] ),
    .B(net126),
    .C(net120),
    .X(_0304_));
 sky130_fd_sc_hd__nand2_1 _0535_ (.A(\count[1] ),
    .B(_0300_),
    .Y(_0305_));
 sky130_fd_sc_hd__nand2_1 _0536_ (.A(_0303_),
    .B(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__xnor2_1 _0537_ (.A(\count[0] ),
    .B(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__mux2_1 _0538_ (.A0(\count[1] ),
    .A1(_0307_),
    .S(_0302_),
    .X(_0001_));
 sky130_fd_sc_hd__xor2_1 _0539_ (.A(\count[2] ),
    .B(_0300_),
    .X(_0308_));
 sky130_fd_sc_hd__a21o_1 _0540_ (.A1(\count[0] ),
    .A2(_0303_),
    .B1(_0304_),
    .X(_0309_));
 sky130_fd_sc_hd__xor2_1 _0541_ (.A(_0308_),
    .B(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _0542_ (.A0(\count[2] ),
    .A1(_0310_),
    .S(_0302_),
    .X(_0002_));
 sky130_fd_sc_hd__xor2_1 _0543_ (.A(\count[3] ),
    .B(_0300_),
    .X(_0311_));
 sky130_fd_sc_hd__a32o_1 _0544_ (.A1(\count[2] ),
    .A2(net1),
    .A3(_0299_),
    .B1(_0308_),
    .B2(_0309_),
    .X(_0312_));
 sky130_fd_sc_hd__xor2_1 _0545_ (.A(_0311_),
    .B(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _0546_ (.A0(\count[3] ),
    .A1(_0313_),
    .S(_0302_),
    .X(_0003_));
 sky130_fd_sc_hd__o21a_1 _0547_ (.A1(\count[3] ),
    .A2(\count[2] ),
    .B1(_0300_),
    .X(_0314_));
 sky130_fd_sc_hd__a31o_1 _0548_ (.A1(_0308_),
    .A2(_0309_),
    .A3(_0311_),
    .B1(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__xnor2_1 _0549_ (.A(\count[4] ),
    .B(_0300_),
    .Y(_0316_));
 sky130_fd_sc_hd__xnor2_1 _0550_ (.A(_0315_),
    .B(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__mux2_1 _0551_ (.A0(\count[4] ),
    .A1(_0317_),
    .S(_0302_),
    .X(_0004_));
 sky130_fd_sc_hd__and4b_1 _0552_ (.A_N(net167),
    .B(net160),
    .C(net172),
    .D(net176),
    .X(_0318_));
 sky130_fd_sc_hd__nor4b_1 _0553_ (.A(net168),
    .B(net166),
    .C(net172),
    .D_N(net178),
    .Y(_0319_));
 sky130_fd_sc_hd__nor4_1 _0554_ (.A(net175),
    .B(net167),
    .C(net165),
    .D(net171),
    .Y(_0320_));
 sky130_fd_sc_hd__or4_1 _0555_ (.A(net177),
    .B(net169),
    .C(net166),
    .D(net173),
    .X(_0321_));
 sky130_fd_sc_hd__and4b_1 _0556_ (.A_N(net176),
    .B(net168),
    .C(net166),
    .D(net172),
    .X(_0322_));
 sky130_fd_sc_hd__and4bb_1 _0557_ (.A_N(net167),
    .B_N(net171),
    .C(net165),
    .D(net175),
    .X(_0323_));
 sky130_fd_sc_hd__and4b_1 _0558_ (.A_N(net167),
    .B(net165),
    .C(net171),
    .D(net175),
    .X(_0324_));
 sky130_fd_sc_hd__and4bb_2 _0559_ (.A_N(net177),
    .B_N(net170),
    .C(net166),
    .D(net174),
    .X(_0325_));
 sky130_fd_sc_hd__and4b_1 _0560_ (.A_N(net177),
    .B(net169),
    .C(net160),
    .D(net173),
    .X(_0326_));
 sky130_fd_sc_hd__or3b_1 _0561_ (.A(net176),
    .B(net172),
    .C_N(net168),
    .X(_0327_));
 sky130_fd_sc_hd__nor2_1 _0562_ (.A(net165),
    .B(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__nor4_1 _0563_ (.A(net175),
    .B(net168),
    .C(net160),
    .D(net171),
    .Y(_0329_));
 sky130_fd_sc_hd__nor2_1 _0564_ (.A(net160),
    .B(_0327_),
    .Y(_0330_));
 sky130_fd_sc_hd__and4_1 _0565_ (.A(net175),
    .B(net167),
    .C(net165),
    .D(net171),
    .X(_0331_));
 sky130_fd_sc_hd__and4b_1 _0566_ (.A_N(net173),
    .B(net169),
    .C(net177),
    .D(net160),
    .X(_0332_));
 sky130_fd_sc_hd__and4_1 _0567_ (.A(net176),
    .B(net169),
    .C(_0294_),
    .D(net173),
    .X(_0333_));
 sky130_fd_sc_hd__and4bb_1 _0568_ (.A_N(net175),
    .B_N(net167),
    .C(net160),
    .D(net172),
    .X(_0334_));
 sky130_fd_sc_hd__and4b_1 _0569_ (.A_N(net171),
    .B(net165),
    .C(net168),
    .D(net176),
    .X(_0335_));
 sky130_fd_sc_hd__a22o_1 _0570_ (.A1(\mem[10][0] ),
    .A2(net137),
    .B1(net131),
    .B2(\mem[13][0] ),
    .X(_0336_));
 sky130_fd_sc_hd__a221o_1 _0571_ (.A1(\mem[9][0] ),
    .A2(net143),
    .B1(net110),
    .B2(\mem[4][0] ),
    .C1(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__a22o_1 _0572_ (.A1(\mem[14][0] ),
    .A2(net147),
    .B1(net140),
    .B2(\mem[11][0] ),
    .X(_0338_));
 sky130_fd_sc_hd__a22o_1 _0573_ (.A1(\mem[1][0] ),
    .A2(net157),
    .B1(net99),
    .B2(\mem[5][0] ),
    .X(_0339_));
 sky130_fd_sc_hd__a221o_1 _0574_ (.A1(\mem[3][0] ),
    .A2(net117),
    .B1(net91),
    .B2(\mem[2][0] ),
    .C1(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__a22o_1 _0575_ (.A1(\mem[12][0] ),
    .A2(net103),
    .B1(net95),
    .B2(\mem[7][0] ),
    .X(_0341_));
 sky130_fd_sc_hd__a221o_1 _0576_ (.A1(\mem[6][0] ),
    .A2(net114),
    .B1(net106),
    .B2(\mem[8][0] ),
    .C1(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__a211o_1 _0577_ (.A1(\mem[15][0] ),
    .A2(net134),
    .B1(_0338_),
    .C1(net154),
    .X(_0343_));
 sky130_fd_sc_hd__or3_1 _0578_ (.A(_0337_),
    .B(_0342_),
    .C(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__o221a_1 _0579_ (.A1(\mem[0][0] ),
    .A2(net151),
    .B1(_0340_),
    .B2(_0344_),
    .C1(net127),
    .X(_0345_));
 sky130_fd_sc_hd__a21o_1 _0580_ (.A1(net22),
    .A2(net121),
    .B1(_0345_),
    .X(_0005_));
 sky130_fd_sc_hd__a22o_1 _0581_ (.A1(\mem[14][1] ),
    .A2(net149),
    .B1(net100),
    .B2(\mem[5][1] ),
    .X(_0346_));
 sky130_fd_sc_hd__a22o_1 _0582_ (.A1(\mem[10][1] ),
    .A2(net137),
    .B1(net131),
    .B2(\mem[13][1] ),
    .X(_0347_));
 sky130_fd_sc_hd__a22o_1 _0583_ (.A1(\mem[11][1] ),
    .A2(net140),
    .B1(net134),
    .B2(\mem[15][1] ),
    .X(_0348_));
 sky130_fd_sc_hd__a221o_1 _0584_ (.A1(\mem[7][1] ),
    .A2(net95),
    .B1(net91),
    .B2(\mem[2][1] ),
    .C1(_0346_),
    .X(_0349_));
 sky130_fd_sc_hd__a221o_1 _0585_ (.A1(\mem[6][1] ),
    .A2(net114),
    .B1(net106),
    .B2(\mem[8][1] ),
    .C1(_0347_),
    .X(_0350_));
 sky130_fd_sc_hd__a22o_1 _0586_ (.A1(\mem[1][1] ),
    .A2(net157),
    .B1(net103),
    .B2(\mem[12][1] ),
    .X(_0351_));
 sky130_fd_sc_hd__a221o_1 _0587_ (.A1(\mem[3][1] ),
    .A2(net117),
    .B1(net143),
    .B2(\mem[9][1] ),
    .C1(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__a211o_1 _0588_ (.A1(\mem[4][1] ),
    .A2(net110),
    .B1(_0348_),
    .C1(net154),
    .X(_0353_));
 sky130_fd_sc_hd__or3_1 _0589_ (.A(_0350_),
    .B(_0352_),
    .C(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__o221a_1 _0590_ (.A1(\mem[0][1] ),
    .A2(net151),
    .B1(_0349_),
    .B2(_0354_),
    .C1(net127),
    .X(_0355_));
 sky130_fd_sc_hd__a21o_1 _0591_ (.A1(net29),
    .A2(net121),
    .B1(_0355_),
    .X(_0006_));
 sky130_fd_sc_hd__a22o_1 _0592_ (.A1(\mem[10][2] ),
    .A2(net137),
    .B1(net91),
    .B2(\mem[2][2] ),
    .X(_0356_));
 sky130_fd_sc_hd__a22o_1 _0593_ (.A1(\mem[12][2] ),
    .A2(net103),
    .B1(net134),
    .B2(\mem[15][2] ),
    .X(_0357_));
 sky130_fd_sc_hd__a22o_1 _0594_ (.A1(\mem[9][2] ),
    .A2(net143),
    .B1(net140),
    .B2(\mem[11][2] ),
    .X(_0358_));
 sky130_fd_sc_hd__a221o_1 _0595_ (.A1(\mem[8][2] ),
    .A2(net108),
    .B1(net132),
    .B2(\mem[13][2] ),
    .C1(_0357_),
    .X(_0359_));
 sky130_fd_sc_hd__a221o_1 _0596_ (.A1(\mem[3][2] ),
    .A2(net117),
    .B1(net95),
    .B2(\mem[7][2] ),
    .C1(_0358_),
    .X(_0360_));
 sky130_fd_sc_hd__a22o_1 _0597_ (.A1(\mem[14][2] ),
    .A2(net147),
    .B1(net99),
    .B2(\mem[5][2] ),
    .X(_0361_));
 sky130_fd_sc_hd__a221o_1 _0598_ (.A1(\mem[1][2] ),
    .A2(net157),
    .B1(net114),
    .B2(\mem[6][2] ),
    .C1(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__a211o_1 _0599_ (.A1(\mem[4][2] ),
    .A2(net110),
    .B1(_0356_),
    .C1(net154),
    .X(_0363_));
 sky130_fd_sc_hd__or3_1 _0600_ (.A(_0360_),
    .B(_0362_),
    .C(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__o221a_1 _0601_ (.A1(\mem[0][2] ),
    .A2(net151),
    .B1(_0359_),
    .B2(_0364_),
    .C1(net127),
    .X(_0365_));
 sky130_fd_sc_hd__a21o_1 _0602_ (.A1(net30),
    .A2(net121),
    .B1(_0365_),
    .X(_0007_));
 sky130_fd_sc_hd__a22o_1 _0603_ (.A1(\mem[11][3] ),
    .A2(net142),
    .B1(net91),
    .B2(\mem[2][3] ),
    .X(_0366_));
 sky130_fd_sc_hd__a22o_1 _0604_ (.A1(\mem[15][3] ),
    .A2(net134),
    .B1(net132),
    .B2(\mem[13][3] ),
    .X(_0367_));
 sky130_fd_sc_hd__a221o_1 _0605_ (.A1(\mem[4][3] ),
    .A2(net110),
    .B1(net95),
    .B2(\mem[7][3] ),
    .C1(_0366_),
    .X(_0368_));
 sky130_fd_sc_hd__a221o_1 _0606_ (.A1(\mem[6][3] ),
    .A2(net115),
    .B1(net108),
    .B2(\mem[8][3] ),
    .C1(_0367_),
    .X(_0369_));
 sky130_fd_sc_hd__a22o_1 _0607_ (.A1(\mem[1][3] ),
    .A2(net157),
    .B1(net143),
    .B2(\mem[9][3] ),
    .X(_0370_));
 sky130_fd_sc_hd__a221o_1 _0608_ (.A1(\mem[10][3] ),
    .A2(net139),
    .B1(net100),
    .B2(\mem[5][3] ),
    .C1(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__a22o_1 _0609_ (.A1(\mem[3][3] ),
    .A2(net119),
    .B1(net149),
    .B2(\mem[14][3] ),
    .X(_0372_));
 sky130_fd_sc_hd__a2111o_1 _0610_ (.A1(\mem[12][3] ),
    .A2(net105),
    .B1(_0371_),
    .C1(_0372_),
    .D1(net154),
    .X(_0373_));
 sky130_fd_sc_hd__or3_1 _0611_ (.A(_0368_),
    .B(_0369_),
    .C(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__o21a_1 _0612_ (.A1(\mem[0][3] ),
    .A2(net153),
    .B1(net126),
    .X(_0375_));
 sky130_fd_sc_hd__a22o_1 _0613_ (.A1(net31),
    .A2(net121),
    .B1(_0374_),
    .B2(_0375_),
    .X(_0008_));
 sky130_fd_sc_hd__and2_1 _0614_ (.A(\mem[5][4] ),
    .B(net99),
    .X(_0376_));
 sky130_fd_sc_hd__a22o_1 _0615_ (.A1(\mem[2][4] ),
    .A2(net91),
    .B1(net131),
    .B2(\mem[13][4] ),
    .X(_0377_));
 sky130_fd_sc_hd__a22o_1 _0616_ (.A1(\mem[14][4] ),
    .A2(net147),
    .B1(net143),
    .B2(\mem[9][4] ),
    .X(_0378_));
 sky130_fd_sc_hd__a221o_1 _0617_ (.A1(\mem[6][4] ),
    .A2(net114),
    .B1(net103),
    .B2(\mem[12][4] ),
    .C1(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__a221o_1 _0618_ (.A1(\mem[3][4] ),
    .A2(net117),
    .B1(net140),
    .B2(\mem[11][4] ),
    .C1(_0377_),
    .X(_0380_));
 sky130_fd_sc_hd__a22o_1 _0619_ (.A1(\mem[10][4] ),
    .A2(net137),
    .B1(net134),
    .B2(\mem[15][4] ),
    .X(_0381_));
 sky130_fd_sc_hd__a221o_1 _0620_ (.A1(\mem[1][4] ),
    .A2(net157),
    .B1(net106),
    .B2(\mem[8][4] ),
    .C1(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__a221o_1 _0621_ (.A1(\mem[4][4] ),
    .A2(net110),
    .B1(net95),
    .B2(\mem[7][4] ),
    .C1(_0376_),
    .X(_0383_));
 sky130_fd_sc_hd__or4_1 _0622_ (.A(net154),
    .B(_0380_),
    .C(_0382_),
    .D(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__o221a_1 _0623_ (.A1(\mem[0][4] ),
    .A2(net151),
    .B1(_0379_),
    .B2(_0384_),
    .C1(net127),
    .X(_0385_));
 sky130_fd_sc_hd__a21o_1 _0624_ (.A1(net32),
    .A2(net121),
    .B1(_0385_),
    .X(_0009_));
 sky130_fd_sc_hd__a22o_1 _0625_ (.A1(\mem[3][5] ),
    .A2(net117),
    .B1(net159),
    .B2(\mem[1][5] ),
    .X(_0386_));
 sky130_fd_sc_hd__a221o_1 _0626_ (.A1(\mem[11][5] ),
    .A2(net140),
    .B1(net96),
    .B2(\mem[7][5] ),
    .C1(net156),
    .X(_0387_));
 sky130_fd_sc_hd__a221o_1 _0627_ (.A1(\mem[10][5] ),
    .A2(_0325_),
    .B1(net132),
    .B2(\mem[13][5] ),
    .C1(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__a211o_1 _0628_ (.A1(\mem[9][5] ),
    .A2(net146),
    .B1(_0386_),
    .C1(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__a22o_1 _0629_ (.A1(\mem[14][5] ),
    .A2(net149),
    .B1(net103),
    .B2(\mem[12][5] ),
    .X(_0390_));
 sky130_fd_sc_hd__a221o_1 _0630_ (.A1(\mem[6][5] ),
    .A2(net115),
    .B1(net100),
    .B2(\mem[5][5] ),
    .C1(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__a22o_1 _0631_ (.A1(\mem[15][5] ),
    .A2(net136),
    .B1(net94),
    .B2(\mem[2][5] ),
    .X(_0392_));
 sky130_fd_sc_hd__a221o_1 _0632_ (.A1(\mem[4][5] ),
    .A2(net113),
    .B1(net108),
    .B2(\mem[8][5] ),
    .C1(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__or3_1 _0633_ (.A(_0389_),
    .B(_0391_),
    .C(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__o21a_1 _0634_ (.A1(\mem[0][5] ),
    .A2(net153),
    .B1(net130),
    .X(_0395_));
 sky130_fd_sc_hd__a22o_1 _0635_ (.A1(net33),
    .A2(net122),
    .B1(_0394_),
    .B2(_0395_),
    .X(_0010_));
 sky130_fd_sc_hd__a22o_1 _0636_ (.A1(\mem[3][6] ),
    .A2(net117),
    .B1(net147),
    .B2(\mem[14][6] ),
    .X(_0396_));
 sky130_fd_sc_hd__a221o_1 _0637_ (.A1(\mem[4][6] ),
    .A2(net110),
    .B1(net99),
    .B2(\mem[5][6] ),
    .C1(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__a22o_1 _0638_ (.A1(\mem[12][6] ),
    .A2(net103),
    .B1(net131),
    .B2(\mem[13][6] ),
    .X(_0398_));
 sky130_fd_sc_hd__a22o_1 _0639_ (.A1(\mem[9][6] ),
    .A2(net143),
    .B1(net134),
    .B2(\mem[15][6] ),
    .X(_0399_));
 sky130_fd_sc_hd__a22o_1 _0640_ (.A1(\mem[10][6] ),
    .A2(net137),
    .B1(net91),
    .B2(\mem[2][6] ),
    .X(_0400_));
 sky130_fd_sc_hd__a221o_1 _0641_ (.A1(\mem[11][6] ),
    .A2(net140),
    .B1(net106),
    .B2(\mem[8][6] ),
    .C1(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__a22o_1 _0642_ (.A1(\mem[1][6] ),
    .A2(net157),
    .B1(net95),
    .B2(\mem[7][6] ),
    .X(_0402_));
 sky130_fd_sc_hd__a211o_1 _0643_ (.A1(\mem[6][6] ),
    .A2(net114),
    .B1(_0402_),
    .C1(net154),
    .X(_0403_));
 sky130_fd_sc_hd__or4_1 _0644_ (.A(_0398_),
    .B(_0399_),
    .C(_0401_),
    .D(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__o221a_1 _0645_ (.A1(\mem[0][6] ),
    .A2(net151),
    .B1(_0397_),
    .B2(_0404_),
    .C1(net127),
    .X(_0405_));
 sky130_fd_sc_hd__a21o_1 _0646_ (.A1(net34),
    .A2(net122),
    .B1(_0405_),
    .X(_0011_));
 sky130_fd_sc_hd__a22o_1 _0647_ (.A1(\mem[10][7] ),
    .A2(net139),
    .B1(net112),
    .B2(\mem[4][7] ),
    .X(_0406_));
 sky130_fd_sc_hd__a22o_1 _0648_ (.A1(\mem[5][7] ),
    .A2(net99),
    .B1(net92),
    .B2(\mem[2][7] ),
    .X(_0407_));
 sky130_fd_sc_hd__a221o_1 _0649_ (.A1(\mem[8][7] ),
    .A2(net108),
    .B1(net96),
    .B2(\mem[7][7] ),
    .C1(_0406_),
    .X(_0408_));
 sky130_fd_sc_hd__a221o_1 _0650_ (.A1(\mem[14][7] ),
    .A2(net149),
    .B1(net142),
    .B2(\mem[11][7] ),
    .C1(_0407_),
    .X(_0409_));
 sky130_fd_sc_hd__a22o_1 _0651_ (.A1(\mem[6][7] ),
    .A2(net115),
    .B1(net132),
    .B2(\mem[13][7] ),
    .X(_0410_));
 sky130_fd_sc_hd__a22o_1 _0652_ (.A1(\mem[1][7] ),
    .A2(net159),
    .B1(net105),
    .B2(\mem[12][7] ),
    .X(_0411_));
 sky130_fd_sc_hd__a22o_1 _0653_ (.A1(\mem[9][7] ),
    .A2(net144),
    .B1(net136),
    .B2(\mem[15][7] ),
    .X(_0412_));
 sky130_fd_sc_hd__a211o_1 _0654_ (.A1(\mem[3][7] ),
    .A2(net119),
    .B1(net156),
    .C1(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__or4_1 _0655_ (.A(_0409_),
    .B(_0410_),
    .C(_0411_),
    .D(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__o221a_1 _0656_ (.A1(\mem[0][7] ),
    .A2(net151),
    .B1(_0408_),
    .B2(_0414_),
    .C1(net128),
    .X(_0415_));
 sky130_fd_sc_hd__a21o_1 _0657_ (.A1(net35),
    .A2(net123),
    .B1(_0415_),
    .X(_0012_));
 sky130_fd_sc_hd__a22o_1 _0658_ (.A1(\mem[3][8] ),
    .A2(net118),
    .B1(net97),
    .B2(\mem[7][8] ),
    .X(_0416_));
 sky130_fd_sc_hd__a221o_1 _0659_ (.A1(\mem[8][8] ),
    .A2(net107),
    .B1(net104),
    .B2(\mem[12][8] ),
    .C1(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__a22o_1 _0660_ (.A1(\mem[9][8] ),
    .A2(net144),
    .B1(net99),
    .B2(\mem[5][8] ),
    .X(_0418_));
 sky130_fd_sc_hd__a221o_1 _0661_ (.A1(\mem[11][8] ),
    .A2(net141),
    .B1(net135),
    .B2(\mem[15][8] ),
    .C1(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__a22o_1 _0662_ (.A1(\mem[6][8] ),
    .A2(net116),
    .B1(net92),
    .B2(\mem[2][8] ),
    .X(_0420_));
 sky130_fd_sc_hd__a22o_1 _0663_ (.A1(\mem[14][8] ),
    .A2(net147),
    .B1(net137),
    .B2(\mem[10][8] ),
    .X(_0421_));
 sky130_fd_sc_hd__a22o_1 _0664_ (.A1(\mem[1][8] ),
    .A2(net158),
    .B1(net133),
    .B2(\mem[13][8] ),
    .X(_0422_));
 sky130_fd_sc_hd__a211o_1 _0665_ (.A1(\mem[4][8] ),
    .A2(net111),
    .B1(_0422_),
    .C1(net155),
    .X(_0423_));
 sky130_fd_sc_hd__or4_1 _0666_ (.A(_0419_),
    .B(_0420_),
    .C(_0421_),
    .D(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__o221a_1 _0667_ (.A1(\mem[0][8] ),
    .A2(net152),
    .B1(_0417_),
    .B2(_0424_),
    .C1(net128),
    .X(_0425_));
 sky130_fd_sc_hd__a21o_1 _0668_ (.A1(net36),
    .A2(net123),
    .B1(_0425_),
    .X(_0013_));
 sky130_fd_sc_hd__and2_1 _0669_ (.A(\mem[10][9] ),
    .B(net139),
    .X(_0426_));
 sky130_fd_sc_hd__a221o_1 _0670_ (.A1(\mem[6][9] ),
    .A2(net115),
    .B1(net101),
    .B2(\mem[5][9] ),
    .C1(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__a221o_1 _0671_ (.A1(\mem[3][9] ),
    .A2(net118),
    .B1(net159),
    .B2(\mem[1][9] ),
    .C1(net155),
    .X(_0428_));
 sky130_fd_sc_hd__a221o_1 _0672_ (.A1(\mem[12][9] ),
    .A2(net105),
    .B1(net98),
    .B2(\mem[7][9] ),
    .C1(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__a22o_1 _0673_ (.A1(\mem[14][9] ),
    .A2(net150),
    .B1(net92),
    .B2(\mem[2][9] ),
    .X(_0430_));
 sky130_fd_sc_hd__a221o_1 _0674_ (.A1(\mem[9][9] ),
    .A2(net144),
    .B1(net108),
    .B2(\mem[8][9] ),
    .C1(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__a22o_1 _0675_ (.A1(\mem[11][9] ),
    .A2(net142),
    .B1(net111),
    .B2(\mem[4][9] ),
    .X(_0432_));
 sky130_fd_sc_hd__a221o_1 _0676_ (.A1(\mem[15][9] ),
    .A2(net135),
    .B1(net133),
    .B2(\mem[13][9] ),
    .C1(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__or3_1 _0677_ (.A(_0429_),
    .B(_0431_),
    .C(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__o221a_1 _0678_ (.A1(\mem[0][9] ),
    .A2(net153),
    .B1(_0427_),
    .B2(_0434_),
    .C1(net128),
    .X(_0435_));
 sky130_fd_sc_hd__a21o_1 _0679_ (.A1(net37),
    .A2(net123),
    .B1(_0435_),
    .X(_0014_));
 sky130_fd_sc_hd__a22o_1 _0680_ (.A1(\mem[4][10] ),
    .A2(net111),
    .B1(net106),
    .B2(\mem[8][10] ),
    .X(_0436_));
 sky130_fd_sc_hd__a22o_1 _0681_ (.A1(\mem[10][10] ),
    .A2(net138),
    .B1(net101),
    .B2(\mem[5][10] ),
    .X(_0437_));
 sky130_fd_sc_hd__a22o_1 _0682_ (.A1(\mem[15][10] ),
    .A2(net135),
    .B1(net93),
    .B2(\mem[2][10] ),
    .X(_0438_));
 sky130_fd_sc_hd__a221o_1 _0683_ (.A1(\mem[9][10] ),
    .A2(net145),
    .B1(net115),
    .B2(\mem[6][10] ),
    .C1(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__a221o_1 _0684_ (.A1(\mem[3][10] ),
    .A2(net118),
    .B1(net158),
    .B2(\mem[1][10] ),
    .C1(_0436_),
    .X(_0440_));
 sky130_fd_sc_hd__a22o_1 _0685_ (.A1(\mem[14][10] ),
    .A2(net147),
    .B1(net141),
    .B2(\mem[11][10] ),
    .X(_0441_));
 sky130_fd_sc_hd__a221o_1 _0686_ (.A1(\mem[12][10] ),
    .A2(net104),
    .B1(net133),
    .B2(\mem[13][10] ),
    .C1(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__a211o_1 _0687_ (.A1(\mem[7][10] ),
    .A2(net97),
    .B1(_0437_),
    .C1(net155),
    .X(_0443_));
 sky130_fd_sc_hd__or3_1 _0688_ (.A(_0440_),
    .B(_0442_),
    .C(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__o221a_1 _0689_ (.A1(\mem[0][10] ),
    .A2(net152),
    .B1(_0439_),
    .B2(_0444_),
    .C1(net128),
    .X(_0445_));
 sky130_fd_sc_hd__a21o_1 _0690_ (.A1(net23),
    .A2(net123),
    .B1(_0445_),
    .X(_0015_));
 sky130_fd_sc_hd__a22o_1 _0691_ (.A1(\mem[6][11] ),
    .A2(net115),
    .B1(net105),
    .B2(\mem[12][11] ),
    .X(_0446_));
 sky130_fd_sc_hd__a21o_1 _0692_ (.A1(\mem[9][11] ),
    .A2(net145),
    .B1(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__a22o_1 _0693_ (.A1(\mem[11][11] ),
    .A2(net141),
    .B1(net135),
    .B2(\mem[15][11] ),
    .X(_0448_));
 sky130_fd_sc_hd__a221o_1 _0694_ (.A1(\mem[3][11] ),
    .A2(net118),
    .B1(net158),
    .B2(\mem[1][11] ),
    .C1(net155),
    .X(_0449_));
 sky130_fd_sc_hd__a22o_1 _0695_ (.A1(\mem[2][11] ),
    .A2(net92),
    .B1(net131),
    .B2(\mem[13][11] ),
    .X(_0450_));
 sky130_fd_sc_hd__a221o_1 _0696_ (.A1(\mem[14][11] ),
    .A2(net148),
    .B1(net107),
    .B2(\mem[8][11] ),
    .C1(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__a22o_1 _0697_ (.A1(\mem[10][11] ),
    .A2(net138),
    .B1(net97),
    .B2(\mem[7][11] ),
    .X(_0452_));
 sky130_fd_sc_hd__a221o_1 _0698_ (.A1(\mem[4][11] ),
    .A2(net111),
    .B1(net101),
    .B2(\mem[5][11] ),
    .C1(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__or4_1 _0699_ (.A(_0448_),
    .B(_0449_),
    .C(_0451_),
    .D(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__o221a_1 _0700_ (.A1(\mem[0][11] ),
    .A2(net153),
    .B1(_0447_),
    .B2(_0454_),
    .C1(net129),
    .X(_0455_));
 sky130_fd_sc_hd__a21o_1 _0701_ (.A1(net24),
    .A2(net123),
    .B1(_0455_),
    .X(_0016_));
 sky130_fd_sc_hd__a22o_1 _0702_ (.A1(\mem[10][12] ),
    .A2(_0325_),
    .B1(net102),
    .B2(\mem[5][12] ),
    .X(_0456_));
 sky130_fd_sc_hd__a221o_1 _0703_ (.A1(\mem[1][12] ),
    .A2(net158),
    .B1(net132),
    .B2(\mem[13][12] ),
    .C1(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__a22o_1 _0704_ (.A1(\mem[9][12] ),
    .A2(net145),
    .B1(net93),
    .B2(\mem[2][12] ),
    .X(_0458_));
 sky130_fd_sc_hd__a221o_1 _0705_ (.A1(\mem[8][12] ),
    .A2(net108),
    .B1(net136),
    .B2(\mem[15][12] ),
    .C1(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__a22o_1 _0706_ (.A1(\mem[3][12] ),
    .A2(net119),
    .B1(net97),
    .B2(\mem[7][12] ),
    .X(_0460_));
 sky130_fd_sc_hd__a221o_1 _0707_ (.A1(\mem[4][12] ),
    .A2(net112),
    .B1(net104),
    .B2(\mem[12][12] ),
    .C1(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__a22o_1 _0708_ (.A1(\mem[11][12] ),
    .A2(net142),
    .B1(net116),
    .B2(\mem[6][12] ),
    .X(_0462_));
 sky130_fd_sc_hd__a211o_1 _0709_ (.A1(\mem[14][12] ),
    .A2(net149),
    .B1(_0462_),
    .C1(net156),
    .X(_0463_));
 sky130_fd_sc_hd__or3_1 _0710_ (.A(_0459_),
    .B(_0461_),
    .C(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__o221a_1 _0711_ (.A1(\mem[0][12] ),
    .A2(net152),
    .B1(_0457_),
    .B2(_0464_),
    .C1(net129),
    .X(_0465_));
 sky130_fd_sc_hd__a21o_1 _0712_ (.A1(net25),
    .A2(net123),
    .B1(_0465_),
    .X(_0017_));
 sky130_fd_sc_hd__and2_1 _0713_ (.A(\mem[9][13] ),
    .B(net144),
    .X(_0466_));
 sky130_fd_sc_hd__a221o_1 _0714_ (.A1(\mem[4][13] ),
    .A2(net111),
    .B1(net104),
    .B2(\mem[12][13] ),
    .C1(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__a22o_1 _0715_ (.A1(\mem[15][13] ),
    .A2(net135),
    .B1(net92),
    .B2(\mem[2][13] ),
    .X(_0468_));
 sky130_fd_sc_hd__a221o_1 _0716_ (.A1(\mem[3][13] ),
    .A2(net118),
    .B1(net158),
    .B2(\mem[1][13] ),
    .C1(net155),
    .X(_0469_));
 sky130_fd_sc_hd__a22o_1 _0717_ (.A1(\mem[5][13] ),
    .A2(net101),
    .B1(net97),
    .B2(\mem[7][13] ),
    .X(_0470_));
 sky130_fd_sc_hd__a221o_1 _0718_ (.A1(\mem[11][13] ),
    .A2(net141),
    .B1(net116),
    .B2(\mem[6][13] ),
    .C1(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__a22o_1 _0719_ (.A1(\mem[14][13] ),
    .A2(net148),
    .B1(net131),
    .B2(\mem[13][13] ),
    .X(_0472_));
 sky130_fd_sc_hd__a221o_1 _0720_ (.A1(\mem[10][13] ),
    .A2(net138),
    .B1(net107),
    .B2(\mem[8][13] ),
    .C1(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__or4_1 _0721_ (.A(_0468_),
    .B(_0469_),
    .C(_0471_),
    .D(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__o221a_1 _0722_ (.A1(\mem[0][13] ),
    .A2(net152),
    .B1(_0467_),
    .B2(_0474_),
    .C1(net128),
    .X(_0475_));
 sky130_fd_sc_hd__a21o_1 _0723_ (.A1(net26),
    .A2(net124),
    .B1(_0475_),
    .X(_0018_));
 sky130_fd_sc_hd__a22o_1 _0724_ (.A1(\mem[6][14] ),
    .A2(net116),
    .B1(net104),
    .B2(\mem[12][14] ),
    .X(_0476_));
 sky130_fd_sc_hd__a22o_1 _0725_ (.A1(\mem[14][14] ),
    .A2(net149),
    .B1(net139),
    .B2(\mem[10][14] ),
    .X(_0477_));
 sky130_fd_sc_hd__a221o_1 _0726_ (.A1(\mem[4][14] ),
    .A2(net112),
    .B1(net98),
    .B2(\mem[7][14] ),
    .C1(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__a22o_1 _0727_ (.A1(\mem[1][14] ),
    .A2(net159),
    .B1(net136),
    .B2(\mem[15][14] ),
    .X(_0479_));
 sky130_fd_sc_hd__a22o_1 _0728_ (.A1(\mem[5][14] ),
    .A2(net101),
    .B1(net132),
    .B2(\mem[13][14] ),
    .X(_0480_));
 sky130_fd_sc_hd__a221o_1 _0729_ (.A1(\mem[3][14] ),
    .A2(net119),
    .B1(net141),
    .B2(\mem[11][14] ),
    .C1(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__a22o_1 _0730_ (.A1(\mem[9][14] ),
    .A2(net144),
    .B1(net93),
    .B2(\mem[2][14] ),
    .X(_0482_));
 sky130_fd_sc_hd__a211o_1 _0731_ (.A1(\mem[8][14] ),
    .A2(net109),
    .B1(_0482_),
    .C1(net156),
    .X(_0483_));
 sky130_fd_sc_hd__or4_1 _0732_ (.A(_0476_),
    .B(_0479_),
    .C(_0481_),
    .D(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__o221a_1 _0733_ (.A1(\mem[0][14] ),
    .A2(net152),
    .B1(_0478_),
    .B2(_0484_),
    .C1(net129),
    .X(_0485_));
 sky130_fd_sc_hd__a21o_1 _0734_ (.A1(net27),
    .A2(net124),
    .B1(_0485_),
    .X(_0019_));
 sky130_fd_sc_hd__a22o_1 _0735_ (.A1(\mem[11][15] ),
    .A2(net141),
    .B1(net101),
    .B2(\mem[5][15] ),
    .X(_0486_));
 sky130_fd_sc_hd__a221o_1 _0736_ (.A1(\mem[3][15] ),
    .A2(net118),
    .B1(net106),
    .B2(\mem[8][15] ),
    .C1(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__a22o_1 _0737_ (.A1(\mem[10][15] ),
    .A2(net138),
    .B1(net135),
    .B2(\mem[15][15] ),
    .X(_0488_));
 sky130_fd_sc_hd__a221o_1 _0738_ (.A1(\mem[6][15] ),
    .A2(net114),
    .B1(net111),
    .B2(\mem[4][15] ),
    .C1(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__a22o_1 _0739_ (.A1(\mem[9][15] ),
    .A2(net144),
    .B1(net133),
    .B2(\mem[13][15] ),
    .X(_0490_));
 sky130_fd_sc_hd__a221o_1 _0740_ (.A1(\mem[14][15] ),
    .A2(net148),
    .B1(net97),
    .B2(\mem[7][15] ),
    .C1(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__a22o_1 _0741_ (.A1(\mem[1][15] ),
    .A2(net158),
    .B1(net92),
    .B2(\mem[2][15] ),
    .X(_0492_));
 sky130_fd_sc_hd__a211o_1 _0742_ (.A1(\mem[12][15] ),
    .A2(net104),
    .B1(_0492_),
    .C1(net155),
    .X(_0493_));
 sky130_fd_sc_hd__or3_1 _0743_ (.A(_0489_),
    .B(_0491_),
    .C(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__o221a_1 _0744_ (.A1(\mem[0][15] ),
    .A2(net152),
    .B1(_0487_),
    .B2(_0494_),
    .C1(net128),
    .X(_0495_));
 sky130_fd_sc_hd__a21o_1 _0745_ (.A1(net28),
    .A2(net124),
    .B1(_0495_),
    .X(_0020_));
 sky130_fd_sc_hd__xnor2_1 _0746_ (.A(net177),
    .B(net122),
    .Y(_0021_));
 sky130_fd_sc_hd__and3_1 _0747_ (.A(net177),
    .B(net173),
    .C(net126),
    .X(_0496_));
 sky130_fd_sc_hd__a21oi_1 _0748_ (.A1(net178),
    .A2(net126),
    .B1(net173),
    .Y(_0497_));
 sky130_fd_sc_hd__nor2_1 _0749_ (.A(_0496_),
    .B(_0497_),
    .Y(_0022_));
 sky130_fd_sc_hd__xor2_1 _0750_ (.A(net169),
    .B(_0496_),
    .X(_0023_));
 sky130_fd_sc_hd__a21oi_1 _0751_ (.A1(net169),
    .A2(_0496_),
    .B1(_0294_),
    .Y(_0498_));
 sky130_fd_sc_hd__a21o_1 _0752_ (.A1(net130),
    .A2(net96),
    .B1(_0498_),
    .X(_0024_));
 sky130_fd_sc_hd__xnor2_1 _0753_ (.A(net163),
    .B(net120),
    .Y(_0025_));
 sky130_fd_sc_hd__nand2_1 _0754_ (.A(net163),
    .B(net161),
    .Y(_0499_));
 sky130_fd_sc_hd__or2_1 _0755_ (.A(net120),
    .B(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__a21o_1 _0756_ (.A1(net163),
    .A2(_0298_),
    .B1(net161),
    .X(_0501_));
 sky130_fd_sc_hd__and2_1 _0757_ (.A(_0500_),
    .B(_0501_),
    .X(_0026_));
 sky130_fd_sc_hd__and4_1 _0758_ (.A(net163),
    .B(net161),
    .C(\wr_ptr[2] ),
    .D(_0298_),
    .X(_0502_));
 sky130_fd_sc_hd__xnor2_1 _0759_ (.A(\wr_ptr[2] ),
    .B(_0500_),
    .Y(_0027_));
 sky130_fd_sc_hd__xnor2_1 _0760_ (.A(_0293_),
    .B(_0502_),
    .Y(_0028_));
 sky130_fd_sc_hd__and4b_1 _0761_ (.A_N(\wr_ptr[2] ),
    .B(_0293_),
    .C(_0298_),
    .D(net203),
    .X(_0503_));
 sky130_fd_sc_hd__or2_1 _0762_ (.A(net164),
    .B(net161),
    .X(_0504_));
 sky130_fd_sc_hd__or3b_1 _0763_ (.A(net163),
    .B(net162),
    .C_N(_0503_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _0764_ (.A0(net202),
    .A1(\mem[0][0] ),
    .S(net87),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _0765_ (.A0(net242),
    .A1(\mem[0][1] ),
    .S(net87),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _0766_ (.A0(net238),
    .A1(\mem[0][2] ),
    .S(net87),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _0767_ (.A0(net235),
    .A1(\mem[0][3] ),
    .S(net87),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _0768_ (.A0(net231),
    .A1(\mem[0][4] ),
    .S(net87),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _0769_ (.A0(net228),
    .A1(\mem[0][5] ),
    .S(net90),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _0770_ (.A0(net223),
    .A1(\mem[0][6] ),
    .S(net87),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _0771_ (.A0(net221),
    .A1(\mem[0][7] ),
    .S(net88),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _0772_ (.A0(net217),
    .A1(\mem[0][8] ),
    .S(net88),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _0773_ (.A0(net214),
    .A1(\mem[0][9] ),
    .S(net88),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _0774_ (.A0(net196),
    .A1(\mem[0][10] ),
    .S(net88),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _0775_ (.A0(net195),
    .A1(\mem[0][11] ),
    .S(net89),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _0776_ (.A0(net192),
    .A1(\mem[0][12] ),
    .S(net89),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _0777_ (.A0(net187),
    .A1(\mem[0][13] ),
    .S(net88),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _0778_ (.A0(net185),
    .A1(\mem[0][14] ),
    .S(net89),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _0779_ (.A0(net180),
    .A1(\mem[0][15] ),
    .S(net88),
    .X(_0044_));
 sky130_fd_sc_hd__nand2b_1 _0780_ (.A_N(net161),
    .B(net164),
    .Y(_0506_));
 sky130_fd_sc_hd__nand3b_1 _0781_ (.A_N(net162),
    .B(_0503_),
    .C(net164),
    .Y(_0507_));
 sky130_fd_sc_hd__mux2_1 _0782_ (.A0(net202),
    .A1(\mem[1][0] ),
    .S(net84),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _0783_ (.A0(net241),
    .A1(\mem[1][1] ),
    .S(net84),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _0784_ (.A0(net238),
    .A1(\mem[1][2] ),
    .S(net84),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _0785_ (.A0(net235),
    .A1(\mem[1][3] ),
    .S(net86),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _0786_ (.A0(net231),
    .A1(\mem[1][4] ),
    .S(net84),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _0787_ (.A0(net226),
    .A1(\mem[1][5] ),
    .S(net86),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _0788_ (.A0(net223),
    .A1(\mem[1][6] ),
    .S(net84),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _0789_ (.A0(net219),
    .A1(\mem[1][7] ),
    .S(net84),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _0790_ (.A0(net217),
    .A1(\mem[1][8] ),
    .S(net85),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _0791_ (.A0(net213),
    .A1(\mem[1][9] ),
    .S(net85),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _0792_ (.A0(net197),
    .A1(\mem[1][10] ),
    .S(net85),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _0793_ (.A0(net194),
    .A1(\mem[1][11] ),
    .S(net85),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _0794_ (.A0(net192),
    .A1(\mem[1][12] ),
    .S(net86),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _0795_ (.A0(net187),
    .A1(\mem[1][13] ),
    .S(net85),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _0796_ (.A0(net184),
    .A1(\mem[1][14] ),
    .S(net86),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _0797_ (.A0(net180),
    .A1(\mem[1][15] ),
    .S(net85),
    .X(_0060_));
 sky130_fd_sc_hd__nand2b_1 _0798_ (.A_N(net164),
    .B(net161),
    .Y(_0508_));
 sky130_fd_sc_hd__nand3b_2 _0799_ (.A_N(net163),
    .B(net162),
    .C(_0503_),
    .Y(_0509_));
 sky130_fd_sc_hd__mux2_1 _0800_ (.A0(net202),
    .A1(\mem[2][0] ),
    .S(net83),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _0801_ (.A0(net242),
    .A1(\mem[2][1] ),
    .S(net83),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _0802_ (.A0(net240),
    .A1(\mem[2][2] ),
    .S(net83),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _0803_ (.A0(net234),
    .A1(\mem[2][3] ),
    .S(net83),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _0804_ (.A0(net230),
    .A1(\mem[2][4] ),
    .S(net83),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _0805_ (.A0(net226),
    .A1(\mem[2][5] ),
    .S(net83),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _0806_ (.A0(net222),
    .A1(\mem[2][6] ),
    .S(net81),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _0807_ (.A0(net219),
    .A1(\mem[2][7] ),
    .S(net81),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _0808_ (.A0(net215),
    .A1(\mem[2][8] ),
    .S(net81),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _0809_ (.A0(net212),
    .A1(\mem[2][9] ),
    .S(net82),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _0810_ (.A0(net196),
    .A1(\mem[2][10] ),
    .S(net82),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _0811_ (.A0(net193),
    .A1(\mem[2][11] ),
    .S(net81),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _0812_ (.A0(net190),
    .A1(\mem[2][12] ),
    .S(net82),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _0813_ (.A0(net186),
    .A1(\mem[2][13] ),
    .S(net81),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _0814_ (.A0(net182),
    .A1(\mem[2][14] ),
    .S(net82),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _0815_ (.A0(net180),
    .A1(\mem[2][15] ),
    .S(net81),
    .X(_0076_));
 sky130_fd_sc_hd__nand2b_1 _0816_ (.A_N(_0499_),
    .B(_0503_),
    .Y(_0510_));
 sky130_fd_sc_hd__mux2_1 _0817_ (.A0(net202),
    .A1(\mem[3][0] ),
    .S(net78),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _0818_ (.A0(net241),
    .A1(\mem[3][1] ),
    .S(net78),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _0819_ (.A0(net238),
    .A1(\mem[3][2] ),
    .S(net78),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _0820_ (.A0(net234),
    .A1(\mem[3][3] ),
    .S(net78),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _0821_ (.A0(net231),
    .A1(\mem[3][4] ),
    .S(net78),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _0822_ (.A0(net227),
    .A1(\mem[3][5] ),
    .S(net80),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _0823_ (.A0(net223),
    .A1(\mem[3][6] ),
    .S(net78),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _0824_ (.A0(net219),
    .A1(\mem[3][7] ),
    .S(net80),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _0825_ (.A0(net217),
    .A1(\mem[3][8] ),
    .S(net79),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _0826_ (.A0(net213),
    .A1(\mem[3][9] ),
    .S(net79),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _0827_ (.A0(net196),
    .A1(\mem[3][10] ),
    .S(net79),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _0828_ (.A0(net194),
    .A1(\mem[3][11] ),
    .S(net79),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _0829_ (.A0(net190),
    .A1(\mem[3][12] ),
    .S(net80),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _0830_ (.A0(net187),
    .A1(\mem[3][13] ),
    .S(net79),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _0831_ (.A0(net182),
    .A1(\mem[3][14] ),
    .S(net80),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _0832_ (.A0(net180),
    .A1(\mem[3][15] ),
    .S(net79),
    .X(_0092_));
 sky130_fd_sc_hd__nand4_2 _0833_ (.A(net204),
    .B(\wr_ptr[2] ),
    .C(_0293_),
    .D(_0298_),
    .Y(_0511_));
 sky130_fd_sc_hd__nor2_1 _0834_ (.A(_0504_),
    .B(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__mux2_1 _0835_ (.A0(\mem[4][0] ),
    .A1(net200),
    .S(net74),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _0836_ (.A0(\mem[4][1] ),
    .A1(net241),
    .S(net74),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _0837_ (.A0(\mem[4][2] ),
    .A1(net240),
    .S(net74),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _0838_ (.A0(\mem[4][3] ),
    .A1(net234),
    .S(net74),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _0839_ (.A0(\mem[4][4] ),
    .A1(net230),
    .S(net74),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _0840_ (.A0(\mem[4][5] ),
    .A1(net228),
    .S(net77),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _0841_ (.A0(\mem[4][6] ),
    .A1(net224),
    .S(net74),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _0842_ (.A0(\mem[4][7] ),
    .A1(net221),
    .S(net76),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _0843_ (.A0(\mem[4][8] ),
    .A1(net216),
    .S(net75),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _0844_ (.A0(\mem[4][9] ),
    .A1(net212),
    .S(net75),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _0845_ (.A0(\mem[4][10] ),
    .A1(net198),
    .S(net75),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _0846_ (.A0(\mem[4][11] ),
    .A1(net194),
    .S(net75),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _0847_ (.A0(\mem[4][12] ),
    .A1(net192),
    .S(net76),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _0848_ (.A0(\mem[4][13] ),
    .A1(net188),
    .S(net75),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _0849_ (.A0(\mem[4][14] ),
    .A1(net185),
    .S(net76),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _0850_ (.A0(\mem[4][15] ),
    .A1(net181),
    .S(net75),
    .X(_0108_));
 sky130_fd_sc_hd__nor2_1 _0851_ (.A(_0506_),
    .B(_0511_),
    .Y(_0513_));
 sky130_fd_sc_hd__mux2_1 _0852_ (.A0(\mem[5][0] ),
    .A1(net3),
    .S(net70),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _0853_ (.A0(\mem[5][1] ),
    .A1(net242),
    .S(net71),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _0854_ (.A0(\mem[5][2] ),
    .A1(net240),
    .S(net70),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _0855_ (.A0(\mem[5][3] ),
    .A1(net235),
    .S(net71),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _0856_ (.A0(\mem[5][4] ),
    .A1(net230),
    .S(net70),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _0857_ (.A0(\mem[5][5] ),
    .A1(net228),
    .S(net71),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _0858_ (.A0(\mem[5][6] ),
    .A1(net224),
    .S(net70),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _0859_ (.A0(\mem[5][7] ),
    .A1(net219),
    .S(net70),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _0860_ (.A0(\mem[5][8] ),
    .A1(net215),
    .S(net70),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _0861_ (.A0(\mem[5][9] ),
    .A1(net214),
    .S(net73),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _0862_ (.A0(\mem[5][10] ),
    .A1(net199),
    .S(net72),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _0863_ (.A0(\mem[5][11] ),
    .A1(net193),
    .S(net72),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _0864_ (.A0(\mem[5][12] ),
    .A1(net192),
    .S(net72),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _0865_ (.A0(\mem[5][13] ),
    .A1(net186),
    .S(net72),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _0866_ (.A0(\mem[5][14] ),
    .A1(net182),
    .S(net72),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _0867_ (.A0(\mem[5][15] ),
    .A1(net180),
    .S(net72),
    .X(_0124_));
 sky130_fd_sc_hd__nor2_1 _0868_ (.A(_0508_),
    .B(_0511_),
    .Y(_0514_));
 sky130_fd_sc_hd__mux2_1 _0869_ (.A0(\mem[6][0] ),
    .A1(net201),
    .S(net67),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _0870_ (.A0(\mem[6][1] ),
    .A1(net243),
    .S(net67),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _0871_ (.A0(\mem[6][2] ),
    .A1(net240),
    .S(net67),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _0872_ (.A0(\mem[6][3] ),
    .A1(net236),
    .S(net68),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _0873_ (.A0(\mem[6][4] ),
    .A1(net231),
    .S(net67),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _0874_ (.A0(\mem[6][5] ),
    .A1(net228),
    .S(net68),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _0875_ (.A0(\mem[6][6] ),
    .A1(net223),
    .S(net67),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _0876_ (.A0(\mem[6][7] ),
    .A1(net221),
    .S(net68),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _0877_ (.A0(\mem[6][8] ),
    .A1(net215),
    .S(net69),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _0878_ (.A0(\mem[6][9] ),
    .A1(net214),
    .S(net68),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _0879_ (.A0(\mem[6][10] ),
    .A1(net196),
    .S(net69),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _0880_ (.A0(\mem[6][11] ),
    .A1(net195),
    .S(net68),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _0881_ (.A0(\mem[6][12] ),
    .A1(net191),
    .S(net68),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _0882_ (.A0(\mem[6][13] ),
    .A1(net187),
    .S(net69),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _0883_ (.A0(\mem[6][14] ),
    .A1(net183),
    .S(net69),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _0884_ (.A0(\mem[6][15] ),
    .A1(net181),
    .S(net67),
    .X(_0140_));
 sky130_fd_sc_hd__nor2_1 _0885_ (.A(_0499_),
    .B(_0511_),
    .Y(_0515_));
 sky130_fd_sc_hd__mux2_1 _0886_ (.A0(\mem[7][0] ),
    .A1(net201),
    .S(net64),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _0887_ (.A0(\mem[7][1] ),
    .A1(net242),
    .S(net64),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _0888_ (.A0(\mem[7][2] ),
    .A1(net238),
    .S(net64),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _0889_ (.A0(\mem[7][3] ),
    .A1(net234),
    .S(net66),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _0890_ (.A0(\mem[7][4] ),
    .A1(net233),
    .S(net64),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _0891_ (.A0(\mem[7][5] ),
    .A1(net226),
    .S(net66),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _0892_ (.A0(\mem[7][6] ),
    .A1(net223),
    .S(net64),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _0893_ (.A0(\mem[7][7] ),
    .A1(net221),
    .S(net64),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _0894_ (.A0(\mem[7][8] ),
    .A1(net217),
    .S(net65),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _0895_ (.A0(\mem[7][9] ),
    .A1(net214),
    .S(net66),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _0896_ (.A0(\mem[7][10] ),
    .A1(net199),
    .S(net65),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _0897_ (.A0(\mem[7][11] ),
    .A1(net193),
    .S(net65),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _0898_ (.A0(\mem[7][12] ),
    .A1(net191),
    .S(net65),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _0899_ (.A0(\mem[7][13] ),
    .A1(net189),
    .S(net65),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _0900_ (.A0(\mem[7][14] ),
    .A1(net185),
    .S(net66),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _0901_ (.A0(\mem[7][15] ),
    .A1(net179),
    .S(net65),
    .X(_0156_));
 sky130_fd_sc_hd__or4b_2 _0902_ (.A(\wr_ptr[2] ),
    .B(_0293_),
    .C(net120),
    .D_N(net203),
    .X(_0516_));
 sky130_fd_sc_hd__nor2_1 _0903_ (.A(_0504_),
    .B(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__mux2_1 _0904_ (.A0(\mem[8][0] ),
    .A1(net201),
    .S(net61),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _0905_ (.A0(\mem[8][1] ),
    .A1(net243),
    .S(net61),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _0906_ (.A0(\mem[8][2] ),
    .A1(net239),
    .S(net61),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _0907_ (.A0(\mem[8][3] ),
    .A1(net236),
    .S(net63),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _0908_ (.A0(\mem[8][4] ),
    .A1(net231),
    .S(net61),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _0909_ (.A0(\mem[8][5] ),
    .A1(net228),
    .S(net63),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _0910_ (.A0(\mem[8][6] ),
    .A1(net222),
    .S(net61),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _0911_ (.A0(\mem[8][7] ),
    .A1(net16),
    .S(net61),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _0912_ (.A0(\mem[8][8] ),
    .A1(net217),
    .S(net62),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _0913_ (.A0(\mem[8][9] ),
    .A1(net213),
    .S(net63),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _0914_ (.A0(\mem[8][10] ),
    .A1(net198),
    .S(net62),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _0915_ (.A0(\mem[8][11] ),
    .A1(net193),
    .S(net62),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _0916_ (.A0(\mem[8][12] ),
    .A1(net191),
    .S(net62),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _0917_ (.A0(\mem[8][13] ),
    .A1(net186),
    .S(net62),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _0918_ (.A0(\mem[8][14] ),
    .A1(net184),
    .S(net63),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _0919_ (.A0(\mem[8][15] ),
    .A1(net180),
    .S(net62),
    .X(_0172_));
 sky130_fd_sc_hd__nor2_2 _0920_ (.A(_0506_),
    .B(_0516_),
    .Y(_0518_));
 sky130_fd_sc_hd__mux2_1 _0921_ (.A0(\mem[9][0] ),
    .A1(net200),
    .S(net60),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _0922_ (.A0(\mem[9][1] ),
    .A1(net241),
    .S(net60),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _0923_ (.A0(\mem[9][2] ),
    .A1(net238),
    .S(net60),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _0924_ (.A0(\mem[9][3] ),
    .A1(net235),
    .S(net60),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _0925_ (.A0(\mem[9][4] ),
    .A1(net232),
    .S(net60),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _0926_ (.A0(\mem[9][5] ),
    .A1(net227),
    .S(net60),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _0927_ (.A0(\mem[9][6] ),
    .A1(net222),
    .S(net58),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _0928_ (.A0(\mem[9][7] ),
    .A1(net219),
    .S(net58),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _0929_ (.A0(\mem[9][8] ),
    .A1(net216),
    .S(net58),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _0930_ (.A0(\mem[9][9] ),
    .A1(net213),
    .S(net58),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _0931_ (.A0(\mem[9][10] ),
    .A1(net196),
    .S(net59),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _0932_ (.A0(\mem[9][11] ),
    .A1(net195),
    .S(net59),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _0933_ (.A0(\mem[9][12] ),
    .A1(net190),
    .S(net59),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _0934_ (.A0(\mem[9][13] ),
    .A1(net188),
    .S(net58),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _0935_ (.A0(\mem[9][14] ),
    .A1(net182),
    .S(net59),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _0936_ (.A0(\mem[9][15] ),
    .A1(net179),
    .S(net58),
    .X(_0188_));
 sky130_fd_sc_hd__nor2_2 _0937_ (.A(_0508_),
    .B(_0516_),
    .Y(_0285_));
 sky130_fd_sc_hd__mux2_1 _0938_ (.A0(\mem[10][0] ),
    .A1(net200),
    .S(net55),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _0939_ (.A0(\mem[10][1] ),
    .A1(net243),
    .S(net55),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _0940_ (.A0(\mem[10][2] ),
    .A1(net240),
    .S(net55),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _0941_ (.A0(\mem[10][3] ),
    .A1(net235),
    .S(net57),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _0942_ (.A0(\mem[10][4] ),
    .A1(net230),
    .S(net55),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _0943_ (.A0(\mem[10][5] ),
    .A1(net226),
    .S(_0285_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _0944_ (.A0(\mem[10][6] ),
    .A1(net222),
    .S(net55),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _0945_ (.A0(\mem[10][7] ),
    .A1(net16),
    .S(net57),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _0946_ (.A0(\mem[10][8] ),
    .A1(net215),
    .S(net55),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _0947_ (.A0(\mem[10][9] ),
    .A1(net18),
    .S(net57),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _0948_ (.A0(\mem[10][10] ),
    .A1(net199),
    .S(net56),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _0949_ (.A0(\mem[10][11] ),
    .A1(net194),
    .S(net56),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _0950_ (.A0(\mem[10][12] ),
    .A1(net6),
    .S(_0285_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _0951_ (.A0(\mem[10][13] ),
    .A1(net186),
    .S(net56),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _0952_ (.A0(\mem[10][14] ),
    .A1(net185),
    .S(net57),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _0953_ (.A0(\mem[10][15] ),
    .A1(net179),
    .S(net56),
    .X(_0204_));
 sky130_fd_sc_hd__nor2_1 _0954_ (.A(_0499_),
    .B(_0516_),
    .Y(_0286_));
 sky130_fd_sc_hd__mux2_1 _0955_ (.A0(\mem[11][0] ),
    .A1(net200),
    .S(net52),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _0956_ (.A0(\mem[11][1] ),
    .A1(net241),
    .S(net52),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _0957_ (.A0(\mem[11][2] ),
    .A1(net238),
    .S(net52),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _0958_ (.A0(\mem[11][3] ),
    .A1(net234),
    .S(net54),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _0959_ (.A0(\mem[11][4] ),
    .A1(net231),
    .S(net52),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _0960_ (.A0(\mem[11][5] ),
    .A1(net226),
    .S(net52),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _0961_ (.A0(\mem[11][6] ),
    .A1(net222),
    .S(net52),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _0962_ (.A0(\mem[11][7] ),
    .A1(net220),
    .S(net54),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _0963_ (.A0(\mem[11][8] ),
    .A1(net216),
    .S(net53),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _0964_ (.A0(\mem[11][9] ),
    .A1(net212),
    .S(net53),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _0965_ (.A0(\mem[11][10] ),
    .A1(net198),
    .S(net53),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _0966_ (.A0(\mem[11][11] ),
    .A1(net194),
    .S(net53),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _0967_ (.A0(\mem[11][12] ),
    .A1(net191),
    .S(net54),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _0968_ (.A0(\mem[11][13] ),
    .A1(net187),
    .S(net53),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _0969_ (.A0(\mem[11][14] ),
    .A1(net183),
    .S(net54),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _0970_ (.A0(\mem[11][15] ),
    .A1(net181),
    .S(net53),
    .X(_0220_));
 sky130_fd_sc_hd__nand4_2 _0971_ (.A(net203),
    .B(\wr_ptr[2] ),
    .C(\wr_ptr[3] ),
    .D(_0298_),
    .Y(_0287_));
 sky130_fd_sc_hd__nor2_1 _0972_ (.A(_0504_),
    .B(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__mux2_1 _0973_ (.A0(\mem[12][0] ),
    .A1(net201),
    .S(net48),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _0974_ (.A0(\mem[12][1] ),
    .A1(net243),
    .S(net48),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _0975_ (.A0(\mem[12][2] ),
    .A1(net239),
    .S(net48),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _0976_ (.A0(\mem[12][3] ),
    .A1(net235),
    .S(net48),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _0977_ (.A0(\mem[12][4] ),
    .A1(net232),
    .S(net48),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _0978_ (.A0(\mem[12][5] ),
    .A1(net228),
    .S(net51),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _0979_ (.A0(\mem[12][6] ),
    .A1(net223),
    .S(net49),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _0980_ (.A0(\mem[12][7] ),
    .A1(net220),
    .S(net48),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _0981_ (.A0(\mem[12][8] ),
    .A1(net218),
    .S(net49),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _0982_ (.A0(\mem[12][9] ),
    .A1(net18),
    .S(net50),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _0983_ (.A0(\mem[12][10] ),
    .A1(net197),
    .S(net49),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _0984_ (.A0(\mem[12][11] ),
    .A1(net195),
    .S(net50),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _0985_ (.A0(\mem[12][12] ),
    .A1(net191),
    .S(net50),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _0986_ (.A0(\mem[12][13] ),
    .A1(net188),
    .S(net49),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _0987_ (.A0(\mem[12][14] ),
    .A1(net183),
    .S(net49),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _0988_ (.A0(\mem[12][15] ),
    .A1(net181),
    .S(net49),
    .X(_0236_));
 sky130_fd_sc_hd__nor2_1 _0989_ (.A(_0506_),
    .B(_0287_),
    .Y(_0289_));
 sky130_fd_sc_hd__mux2_1 _0990_ (.A0(\mem[13][0] ),
    .A1(net200),
    .S(net45),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _0991_ (.A0(\mem[13][1] ),
    .A1(net243),
    .S(net45),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _0992_ (.A0(\mem[13][2] ),
    .A1(net239),
    .S(net46),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _0993_ (.A0(\mem[13][3] ),
    .A1(net234),
    .S(net46),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _0994_ (.A0(\mem[13][4] ),
    .A1(net230),
    .S(net45),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _0995_ (.A0(\mem[13][5] ),
    .A1(net226),
    .S(net46),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _0996_ (.A0(\mem[13][6] ),
    .A1(net222),
    .S(net47),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _0997_ (.A0(\mem[13][7] ),
    .A1(net220),
    .S(net46),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _0998_ (.A0(\mem[13][8] ),
    .A1(net217),
    .S(net47),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _0999_ (.A0(\mem[13][9] ),
    .A1(net212),
    .S(net47),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _1000_ (.A0(\mem[13][10] ),
    .A1(net197),
    .S(net47),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _1001_ (.A0(\mem[13][11] ),
    .A1(net193),
    .S(net45),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _1002_ (.A0(\mem[13][12] ),
    .A1(net190),
    .S(net46),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _1003_ (.A0(\mem[13][13] ),
    .A1(net186),
    .S(net45),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _1004_ (.A0(\mem[13][14] ),
    .A1(net182),
    .S(net46),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _1005_ (.A0(\mem[13][15] ),
    .A1(net179),
    .S(net45),
    .X(_0252_));
 sky130_fd_sc_hd__nor2_1 _1006_ (.A(_0508_),
    .B(_0287_),
    .Y(_0290_));
 sky130_fd_sc_hd__mux2_1 _1007_ (.A0(\mem[14][0] ),
    .A1(net200),
    .S(net41),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _1008_ (.A0(\mem[14][1] ),
    .A1(net242),
    .S(net43),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _1009_ (.A0(\mem[14][2] ),
    .A1(net240),
    .S(net41),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _1010_ (.A0(\mem[14][3] ),
    .A1(net236),
    .S(net43),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _1011_ (.A0(\mem[14][4] ),
    .A1(net232),
    .S(net41),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _1012_ (.A0(\mem[14][5] ),
    .A1(net229),
    .S(net43),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _1013_ (.A0(\mem[14][6] ),
    .A1(net224),
    .S(net41),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _1014_ (.A0(\mem[14][7] ),
    .A1(net220),
    .S(net43),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _1015_ (.A0(\mem[14][8] ),
    .A1(net215),
    .S(net41),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _1016_ (.A0(\mem[14][9] ),
    .A1(net212),
    .S(net44),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _1017_ (.A0(\mem[14][10] ),
    .A1(net198),
    .S(net41),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _1018_ (.A0(\mem[14][11] ),
    .A1(net193),
    .S(net42),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _1019_ (.A0(\mem[14][12] ),
    .A1(net190),
    .S(net43),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _1020_ (.A0(\mem[14][13] ),
    .A1(net186),
    .S(net42),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _1021_ (.A0(\mem[14][14] ),
    .A1(net185),
    .S(net43),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _1022_ (.A0(\mem[14][15] ),
    .A1(net179),
    .S(net42),
    .X(_0268_));
 sky130_fd_sc_hd__nor2_1 _1023_ (.A(_0499_),
    .B(_0287_),
    .Y(_0291_));
 sky130_fd_sc_hd__mux2_1 _1024_ (.A0(\mem[15][0] ),
    .A1(net201),
    .S(net38),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _1025_ (.A0(\mem[15][1] ),
    .A1(net241),
    .S(net38),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _1026_ (.A0(\mem[15][2] ),
    .A1(net239),
    .S(net38),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _1027_ (.A0(\mem[15][3] ),
    .A1(net237),
    .S(net40),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _1028_ (.A0(\mem[15][4] ),
    .A1(net230),
    .S(net38),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _1029_ (.A0(\mem[15][5] ),
    .A1(net227),
    .S(net38),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _1030_ (.A0(\mem[15][6] ),
    .A1(net225),
    .S(net38),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _1031_ (.A0(\mem[15][7] ),
    .A1(net219),
    .S(net40),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _1032_ (.A0(\mem[15][8] ),
    .A1(net215),
    .S(net39),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _1033_ (.A0(\mem[15][9] ),
    .A1(net212),
    .S(net39),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _1034_ (.A0(\mem[15][10] ),
    .A1(net196),
    .S(net39),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _1035_ (.A0(\mem[15][11] ),
    .A1(net195),
    .S(net39),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _1036_ (.A0(\mem[15][12] ),
    .A1(net190),
    .S(net40),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _1037_ (.A0(\mem[15][13] ),
    .A1(net187),
    .S(net39),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _1038_ (.A0(\mem[15][14] ),
    .A1(net182),
    .S(net40),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _1039_ (.A0(\mem[15][15] ),
    .A1(net179),
    .S(net39),
    .X(_0284_));
 sky130_fd_sc_hd__dfrtp_1 _1040_ (.CLK(clknet_leaf_21_clk),
    .D(_0000_),
    .RESET_B(net205),
    .Q(\count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1041_ (.CLK(clknet_leaf_20_clk),
    .D(_0001_),
    .RESET_B(net205),
    .Q(\count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1042_ (.CLK(clknet_leaf_21_clk),
    .D(_0002_),
    .RESET_B(net203),
    .Q(\count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1043_ (.CLK(clknet_leaf_21_clk),
    .D(_0003_),
    .RESET_B(net205),
    .Q(\count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _1044_ (.CLK(clknet_leaf_21_clk),
    .D(_0004_),
    .RESET_B(net205),
    .Q(\count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1045_ (.CLK(clknet_leaf_20_clk),
    .D(_0005_),
    .RESET_B(net205),
    .Q(net22));
 sky130_fd_sc_hd__dfrtp_1 _1046_ (.CLK(clknet_leaf_20_clk),
    .D(_0006_),
    .RESET_B(net205),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_1 _1047_ (.CLK(clknet_leaf_20_clk),
    .D(_0007_),
    .RESET_B(net206),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_1 _1048_ (.CLK(clknet_leaf_19_clk),
    .D(_0008_),
    .RESET_B(net207),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_1 _1049_ (.CLK(clknet_leaf_19_clk),
    .D(_0009_),
    .RESET_B(net207),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_1 _1050_ (.CLK(clknet_leaf_19_clk),
    .D(_0010_),
    .RESET_B(net207),
    .Q(net33));
 sky130_fd_sc_hd__dfrtp_1 _1051_ (.CLK(clknet_leaf_19_clk),
    .D(_0011_),
    .RESET_B(net207),
    .Q(net34));
 sky130_fd_sc_hd__dfrtp_1 _1052_ (.CLK(clknet_leaf_15_clk),
    .D(_0012_),
    .RESET_B(net209),
    .Q(net35));
 sky130_fd_sc_hd__dfrtp_1 _1053_ (.CLK(clknet_leaf_15_clk),
    .D(_0013_),
    .RESET_B(net209),
    .Q(net36));
 sky130_fd_sc_hd__dfrtp_1 _1054_ (.CLK(clknet_leaf_14_clk),
    .D(_0014_),
    .RESET_B(net209),
    .Q(net37));
 sky130_fd_sc_hd__dfrtp_1 _1055_ (.CLK(clknet_leaf_14_clk),
    .D(_0015_),
    .RESET_B(net209),
    .Q(net23));
 sky130_fd_sc_hd__dfrtp_1 _1056_ (.CLK(clknet_leaf_14_clk),
    .D(_0016_),
    .RESET_B(net209),
    .Q(net24));
 sky130_fd_sc_hd__dfrtp_1 _1057_ (.CLK(clknet_leaf_14_clk),
    .D(_0017_),
    .RESET_B(net210),
    .Q(net25));
 sky130_fd_sc_hd__dfrtp_1 _1058_ (.CLK(clknet_leaf_13_clk),
    .D(_0018_),
    .RESET_B(net210),
    .Q(net26));
 sky130_fd_sc_hd__dfrtp_1 _1059_ (.CLK(clknet_leaf_13_clk),
    .D(_0019_),
    .RESET_B(net210),
    .Q(net27));
 sky130_fd_sc_hd__dfrtp_1 _1060_ (.CLK(clknet_leaf_13_clk),
    .D(_0020_),
    .RESET_B(net210),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_1 _1061_ (.CLK(clknet_leaf_19_clk),
    .D(_0021_),
    .RESET_B(net207),
    .Q(\rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1062_ (.CLK(clknet_leaf_18_clk),
    .D(_0022_),
    .RESET_B(net207),
    .Q(\rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1063_ (.CLK(clknet_leaf_18_clk),
    .D(_0023_),
    .RESET_B(net209),
    .Q(\rd_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1064_ (.CLK(clknet_leaf_18_clk),
    .D(_0024_),
    .RESET_B(net208),
    .Q(\rd_ptr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1065_ (.CLK(clknet_leaf_22_clk),
    .D(_0025_),
    .RESET_B(net203),
    .Q(\wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1066_ (.CLK(clknet_leaf_22_clk),
    .D(_0026_),
    .RESET_B(net203),
    .Q(\wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_2 _1067_ (.CLK(clknet_leaf_22_clk),
    .D(_0027_),
    .RESET_B(net204),
    .Q(\wr_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1068_ (.CLK(clknet_leaf_21_clk),
    .D(_0028_),
    .RESET_B(net204),
    .Q(\wr_ptr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1069_ (.CLK(clknet_leaf_26_clk),
    .D(_0029_),
    .Q(\mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1070_ (.CLK(clknet_leaf_22_clk),
    .D(_0030_),
    .Q(\mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1071_ (.CLK(clknet_leaf_24_clk),
    .D(_0031_),
    .Q(\mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1072_ (.CLK(clknet_leaf_19_clk),
    .D(_0032_),
    .Q(\mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1073_ (.CLK(clknet_leaf_24_clk),
    .D(_0033_),
    .Q(\mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1074_ (.CLK(clknet_leaf_18_clk),
    .D(_0034_),
    .Q(\mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1075_ (.CLK(clknet_leaf_2_clk),
    .D(_0035_),
    .Q(\mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1076_ (.CLK(clknet_leaf_15_clk),
    .D(_0036_),
    .Q(\mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1077_ (.CLK(clknet_leaf_10_clk),
    .D(_0037_),
    .Q(\mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1078_ (.CLK(clknet_leaf_14_clk),
    .D(_0038_),
    .Q(\mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1079_ (.CLK(clknet_leaf_11_clk),
    .D(_0039_),
    .Q(\mem[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1080_ (.CLK(clknet_leaf_14_clk),
    .D(_0040_),
    .Q(\mem[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1081_ (.CLK(clknet_leaf_13_clk),
    .D(_0041_),
    .Q(\mem[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1082_ (.CLK(clknet_leaf_8_clk),
    .D(_0042_),
    .Q(\mem[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1083_ (.CLK(clknet_leaf_13_clk),
    .D(_0043_),
    .Q(\mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1084_ (.CLK(clknet_leaf_8_clk),
    .D(_0044_),
    .Q(\mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1085_ (.CLK(clknet_leaf_25_clk),
    .D(_0045_),
    .Q(\mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1086_ (.CLK(clknet_leaf_26_clk),
    .D(_0046_),
    .Q(\mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1087_ (.CLK(clknet_leaf_1_clk),
    .D(_0047_),
    .Q(\mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1088_ (.CLK(clknet_leaf_21_clk),
    .D(_0048_),
    .Q(\mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1089_ (.CLK(clknet_leaf_1_clk),
    .D(_0049_),
    .Q(\mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1090_ (.CLK(clknet_leaf_24_clk),
    .D(_0050_),
    .Q(\mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1091_ (.CLK(clknet_leaf_1_clk),
    .D(_0051_),
    .Q(\mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1092_ (.CLK(clknet_leaf_17_clk),
    .D(_0052_),
    .Q(\mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1093_ (.CLK(clknet_leaf_3_clk),
    .D(_0053_),
    .Q(\mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1094_ (.CLK(clknet_leaf_16_clk),
    .D(_0054_),
    .Q(\mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1095_ (.CLK(clknet_leaf_9_clk),
    .D(_0055_),
    .Q(\mem[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1096_ (.CLK(clknet_leaf_3_clk),
    .D(_0056_),
    .Q(\mem[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1097_ (.CLK(clknet_leaf_13_clk),
    .D(_0057_),
    .Q(\mem[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1098_ (.CLK(clknet_leaf_7_clk),
    .D(_0058_),
    .Q(\mem[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1099_ (.CLK(clknet_leaf_11_clk),
    .D(_0059_),
    .Q(\mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1100_ (.CLK(clknet_leaf_7_clk),
    .D(_0060_),
    .Q(\mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1101_ (.CLK(clknet_leaf_25_clk),
    .D(_0061_),
    .Q(\mem[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1102_ (.CLK(clknet_leaf_22_clk),
    .D(_0062_),
    .Q(\mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1103_ (.CLK(clknet_leaf_0_clk),
    .D(_0063_),
    .Q(\mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1104_ (.CLK(clknet_leaf_23_clk),
    .D(_0064_),
    .Q(\mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1105_ (.CLK(clknet_leaf_0_clk),
    .D(_0065_),
    .Q(\mem[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1106_ (.CLK(clknet_leaf_17_clk),
    .D(_0066_),
    .Q(\mem[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1107_ (.CLK(clknet_leaf_0_clk),
    .D(_0067_),
    .Q(\mem[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1108_ (.CLK(clknet_leaf_10_clk),
    .D(_0068_),
    .Q(\mem[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1109_ (.CLK(clknet_leaf_4_clk),
    .D(_0069_),
    .Q(\mem[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1110_ (.CLK(clknet_leaf_11_clk),
    .D(_0070_),
    .Q(\mem[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1111_ (.CLK(clknet_leaf_10_clk),
    .D(_0071_),
    .Q(\mem[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1112_ (.CLK(clknet_leaf_4_clk),
    .D(_0072_),
    .Q(\mem[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1113_ (.CLK(clknet_leaf_11_clk),
    .D(_0073_),
    .Q(\mem[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1114_ (.CLK(clknet_leaf_7_clk),
    .D(_0074_),
    .Q(\mem[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1115_ (.CLK(clknet_leaf_11_clk),
    .D(_0075_),
    .Q(\mem[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1116_ (.CLK(clknet_leaf_7_clk),
    .D(_0076_),
    .Q(\mem[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1117_ (.CLK(clknet_leaf_26_clk),
    .D(_0077_),
    .Q(\mem[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1118_ (.CLK(clknet_leaf_26_clk),
    .D(_0078_),
    .Q(\mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1119_ (.CLK(clknet_leaf_25_clk),
    .D(_0079_),
    .Q(\mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1120_ (.CLK(clknet_leaf_23_clk),
    .D(_0080_),
    .Q(\mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1121_ (.CLK(clknet_leaf_1_clk),
    .D(_0081_),
    .Q(\mem[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1122_ (.CLK(clknet_leaf_17_clk),
    .D(_0082_),
    .Q(\mem[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1123_ (.CLK(clknet_leaf_2_clk),
    .D(_0083_),
    .Q(\mem[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1124_ (.CLK(clknet_leaf_17_clk),
    .D(_0084_),
    .Q(\mem[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1125_ (.CLK(clknet_leaf_2_clk),
    .D(_0085_),
    .Q(\mem[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1126_ (.CLK(clknet_leaf_16_clk),
    .D(_0086_),
    .Q(\mem[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1127_ (.CLK(clknet_leaf_10_clk),
    .D(_0087_),
    .Q(\mem[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1128_ (.CLK(clknet_leaf_9_clk),
    .D(_0088_),
    .Q(\mem[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1129_ (.CLK(clknet_leaf_13_clk),
    .D(_0089_),
    .Q(\mem[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1130_ (.CLK(clknet_leaf_7_clk),
    .D(_0090_),
    .Q(\mem[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1131_ (.CLK(clknet_leaf_8_clk),
    .D(_0091_),
    .Q(\mem[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1132_ (.CLK(clknet_leaf_8_clk),
    .D(_0092_),
    .Q(\mem[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1133_ (.CLK(clknet_leaf_28_clk),
    .D(_0093_),
    .Q(\mem[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1134_ (.CLK(clknet_leaf_25_clk),
    .D(_0094_),
    .Q(\mem[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1135_ (.CLK(clknet_leaf_28_clk),
    .D(_0095_),
    .Q(\mem[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1136_ (.CLK(clknet_leaf_23_clk),
    .D(_0096_),
    .Q(\mem[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1137_ (.CLK(clknet_leaf_1_clk),
    .D(_0097_),
    .Q(\mem[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1138_ (.CLK(clknet_leaf_17_clk),
    .D(_0098_),
    .Q(\mem[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1139_ (.CLK(clknet_leaf_2_clk),
    .D(_0099_),
    .Q(\mem[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1140_ (.CLK(clknet_leaf_15_clk),
    .D(_0100_),
    .Q(\mem[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1141_ (.CLK(clknet_leaf_3_clk),
    .D(_0101_),
    .Q(\mem[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1142_ (.CLK(clknet_leaf_10_clk),
    .D(_0102_),
    .Q(\mem[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1143_ (.CLK(clknet_leaf_9_clk),
    .D(_0103_),
    .Q(\mem[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1144_ (.CLK(clknet_leaf_3_clk),
    .D(_0104_),
    .Q(\mem[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1145_ (.CLK(clknet_leaf_13_clk),
    .D(_0105_),
    .Q(\mem[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1146_ (.CLK(clknet_leaf_9_clk),
    .D(_0106_),
    .Q(\mem[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1147_ (.CLK(clknet_leaf_13_clk),
    .D(_0107_),
    .Q(\mem[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1148_ (.CLK(clknet_leaf_6_clk),
    .D(_0108_),
    .Q(\mem[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1149_ (.CLK(clknet_leaf_25_clk),
    .D(_0109_),
    .Q(\mem[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1150_ (.CLK(clknet_leaf_23_clk),
    .D(_0110_),
    .Q(\mem[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1151_ (.CLK(clknet_leaf_28_clk),
    .D(_0111_),
    .Q(\mem[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1152_ (.CLK(clknet_leaf_20_clk),
    .D(_0112_),
    .Q(\mem[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1153_ (.CLK(clknet_leaf_0_clk),
    .D(_0113_),
    .Q(\mem[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1154_ (.CLK(clknet_leaf_18_clk),
    .D(_0114_),
    .Q(\mem[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1155_ (.CLK(clknet_leaf_2_clk),
    .D(_0115_),
    .Q(\mem[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1156_ (.CLK(clknet_leaf_10_clk),
    .D(_0116_),
    .Q(\mem[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1157_ (.CLK(clknet_leaf_4_clk),
    .D(_0117_),
    .Q(\mem[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1158_ (.CLK(clknet_leaf_15_clk),
    .D(_0118_),
    .Q(\mem[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1159_ (.CLK(clknet_leaf_5_clk),
    .D(_0119_),
    .Q(\mem[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1160_ (.CLK(clknet_leaf_3_clk),
    .D(_0120_),
    .Q(\mem[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1161_ (.CLK(clknet_leaf_13_clk),
    .D(_0121_),
    .Q(\mem[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1162_ (.CLK(clknet_leaf_6_clk),
    .D(_0122_),
    .Q(\mem[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1163_ (.CLK(clknet_leaf_8_clk),
    .D(_0123_),
    .Q(\mem[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1164_ (.CLK(clknet_leaf_7_clk),
    .D(_0124_),
    .Q(\mem[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1165_ (.CLK(clknet_leaf_26_clk),
    .D(_0125_),
    .Q(\mem[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1166_ (.CLK(clknet_leaf_28_clk),
    .D(_0126_),
    .Q(\mem[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1167_ (.CLK(clknet_leaf_1_clk),
    .D(_0127_),
    .Q(\mem[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1168_ (.CLK(clknet_leaf_18_clk),
    .D(_0128_),
    .Q(\mem[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1169_ (.CLK(clknet_leaf_1_clk),
    .D(_0129_),
    .Q(\mem[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1170_ (.CLK(clknet_leaf_19_clk),
    .D(_0130_),
    .Q(\mem[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1171_ (.CLK(clknet_leaf_1_clk),
    .D(_0131_),
    .Q(\mem[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1172_ (.CLK(clknet_leaf_16_clk),
    .D(_0132_),
    .Q(\mem[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1173_ (.CLK(clknet_leaf_4_clk),
    .D(_0133_),
    .Q(\mem[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1174_ (.CLK(clknet_leaf_14_clk),
    .D(_0134_),
    .Q(\mem[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1175_ (.CLK(clknet_leaf_9_clk),
    .D(_0135_),
    .Q(\mem[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1176_ (.CLK(clknet_leaf_13_clk),
    .D(_0136_),
    .Q(\mem[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1177_ (.CLK(clknet_leaf_12_clk),
    .D(_0137_),
    .Q(\mem[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1178_ (.CLK(clknet_leaf_7_clk),
    .D(_0138_),
    .Q(\mem[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1179_ (.CLK(clknet_leaf_12_clk),
    .D(_0139_),
    .Q(\mem[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1180_ (.CLK(clknet_leaf_6_clk),
    .D(_0140_),
    .Q(\mem[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1181_ (.CLK(clknet_leaf_27_clk),
    .D(_0141_),
    .Q(\mem[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1182_ (.CLK(clknet_leaf_22_clk),
    .D(_0142_),
    .Q(\mem[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1183_ (.CLK(clknet_leaf_25_clk),
    .D(_0143_),
    .Q(\mem[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1184_ (.CLK(clknet_leaf_23_clk),
    .D(_0144_),
    .Q(\mem[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1185_ (.CLK(clknet_leaf_1_clk),
    .D(_0145_),
    .Q(\mem[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1186_ (.CLK(clknet_leaf_24_clk),
    .D(_0146_),
    .Q(\mem[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1187_ (.CLK(clknet_leaf_2_clk),
    .D(_0147_),
    .Q(\mem[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1188_ (.CLK(clknet_leaf_15_clk),
    .D(_0148_),
    .Q(\mem[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1189_ (.CLK(clknet_leaf_2_clk),
    .D(_0149_),
    .Q(\mem[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1190_ (.CLK(clknet_leaf_16_clk),
    .D(_0150_),
    .Q(\mem[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1191_ (.CLK(clknet_leaf_5_clk),
    .D(_0151_),
    .Q(\mem[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1192_ (.CLK(clknet_leaf_4_clk),
    .D(_0152_),
    .Q(\mem[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1193_ (.CLK(clknet_leaf_12_clk),
    .D(_0153_),
    .Q(\mem[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1194_ (.CLK(clknet_leaf_6_clk),
    .D(_0154_),
    .Q(\mem[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1195_ (.CLK(clknet_leaf_13_clk),
    .D(_0155_),
    .Q(\mem[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1196_ (.CLK(clknet_leaf_7_clk),
    .D(_0156_),
    .Q(\mem[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1197_ (.CLK(clknet_leaf_27_clk),
    .D(_0157_),
    .Q(\mem[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1198_ (.CLK(clknet_leaf_28_clk),
    .D(_0158_),
    .Q(\mem[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1199_ (.CLK(clknet_leaf_25_clk),
    .D(_0159_),
    .Q(\mem[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1200_ (.CLK(clknet_leaf_23_clk),
    .D(_0160_),
    .Q(\mem[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1201_ (.CLK(clknet_leaf_1_clk),
    .D(_0161_),
    .Q(\mem[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1202_ (.CLK(clknet_leaf_17_clk),
    .D(_0162_),
    .Q(\mem[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1203_ (.CLK(clknet_leaf_4_clk),
    .D(_0163_),
    .Q(\mem[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1204_ (.CLK(clknet_leaf_16_clk),
    .D(_0164_),
    .Q(\mem[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1205_ (.CLK(clknet_leaf_2_clk),
    .D(_0165_),
    .Q(\mem[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1206_ (.CLK(clknet_leaf_11_clk),
    .D(_0166_),
    .Q(\mem[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1207_ (.CLK(clknet_leaf_9_clk),
    .D(_0167_),
    .Q(\mem[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1208_ (.CLK(clknet_leaf_4_clk),
    .D(_0168_),
    .Q(\mem[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1209_ (.CLK(clknet_leaf_12_clk),
    .D(_0169_),
    .Q(\mem[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1210_ (.CLK(clknet_leaf_6_clk),
    .D(_0170_),
    .Q(\mem[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1211_ (.CLK(clknet_leaf_12_clk),
    .D(_0171_),
    .Q(\mem[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1212_ (.CLK(clknet_leaf_8_clk),
    .D(_0172_),
    .Q(\mem[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1213_ (.CLK(clknet_leaf_27_clk),
    .D(_0173_),
    .Q(\mem[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1214_ (.CLK(clknet_leaf_26_clk),
    .D(_0174_),
    .Q(\mem[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1215_ (.CLK(clknet_leaf_25_clk),
    .D(_0175_),
    .Q(\mem[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1216_ (.CLK(clknet_leaf_22_clk),
    .D(_0176_),
    .Q(\mem[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1217_ (.CLK(clknet_leaf_1_clk),
    .D(_0177_),
    .Q(\mem[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1218_ (.CLK(clknet_leaf_23_clk),
    .D(_0178_),
    .Q(\mem[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1219_ (.CLK(clknet_leaf_1_clk),
    .D(_0179_),
    .Q(\mem[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1220_ (.CLK(clknet_leaf_17_clk),
    .D(_0180_),
    .Q(\mem[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1221_ (.CLK(clknet_leaf_3_clk),
    .D(_0181_),
    .Q(\mem[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1222_ (.CLK(clknet_leaf_11_clk),
    .D(_0182_),
    .Q(\mem[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1223_ (.CLK(clknet_leaf_10_clk),
    .D(_0183_),
    .Q(\mem[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1224_ (.CLK(clknet_leaf_14_clk),
    .D(_0184_),
    .Q(\mem[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1225_ (.CLK(clknet_leaf_11_clk),
    .D(_0185_),
    .Q(\mem[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1226_ (.CLK(clknet_leaf_9_clk),
    .D(_0186_),
    .Q(\mem[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1227_ (.CLK(clknet_leaf_11_clk),
    .D(_0187_),
    .Q(\mem[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1228_ (.CLK(clknet_leaf_5_clk),
    .D(_0188_),
    .Q(\mem[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1229_ (.CLK(clknet_leaf_28_clk),
    .D(_0189_),
    .Q(\mem[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1230_ (.CLK(clknet_leaf_28_clk),
    .D(_0190_),
    .Q(\mem[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1231_ (.CLK(clknet_leaf_0_clk),
    .D(_0191_),
    .Q(\mem[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1232_ (.CLK(clknet_leaf_20_clk),
    .D(_0192_),
    .Q(\mem[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1233_ (.CLK(clknet_leaf_0_clk),
    .D(_0193_),
    .Q(\mem[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1234_ (.CLK(clknet_leaf_23_clk),
    .D(_0194_),
    .Q(\mem[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1235_ (.CLK(clknet_leaf_0_clk),
    .D(_0195_),
    .Q(\mem[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1236_ (.CLK(clknet_leaf_15_clk),
    .D(_0196_),
    .Q(\mem[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1237_ (.CLK(clknet_leaf_4_clk),
    .D(_0197_),
    .Q(\mem[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1238_ (.CLK(clknet_leaf_15_clk),
    .D(_0198_),
    .Q(\mem[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1239_ (.CLK(clknet_leaf_5_clk),
    .D(_0199_),
    .Q(\mem[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1240_ (.CLK(clknet_leaf_4_clk),
    .D(_0200_),
    .Q(\mem[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1241_ (.CLK(clknet_leaf_14_clk),
    .D(_0201_),
    .Q(\mem[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1242_ (.CLK(clknet_leaf_6_clk),
    .D(_0202_),
    .Q(\mem[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1243_ (.CLK(clknet_leaf_13_clk),
    .D(_0203_),
    .Q(\mem[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1244_ (.CLK(clknet_leaf_5_clk),
    .D(_0204_),
    .Q(\mem[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1245_ (.CLK(clknet_leaf_28_clk),
    .D(_0205_),
    .Q(\mem[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1246_ (.CLK(clknet_leaf_25_clk),
    .D(_0206_),
    .Q(\mem[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1247_ (.CLK(clknet_leaf_28_clk),
    .D(_0207_),
    .Q(\mem[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1248_ (.CLK(clknet_leaf_23_clk),
    .D(_0208_),
    .Q(\mem[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1249_ (.CLK(clknet_leaf_1_clk),
    .D(_0209_),
    .Q(\mem[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1250_ (.CLK(clknet_leaf_24_clk),
    .D(_0210_),
    .Q(\mem[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1251_ (.CLK(clknet_leaf_0_clk),
    .D(_0211_),
    .Q(\mem[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1252_ (.CLK(clknet_leaf_10_clk),
    .D(_0212_),
    .Q(\mem[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1253_ (.CLK(clknet_leaf_3_clk),
    .D(_0213_),
    .Q(\mem[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1254_ (.CLK(clknet_leaf_11_clk),
    .D(_0214_),
    .Q(\mem[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1255_ (.CLK(clknet_leaf_9_clk),
    .D(_0215_),
    .Q(\mem[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1256_ (.CLK(clknet_leaf_9_clk),
    .D(_0216_),
    .Q(\mem[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1257_ (.CLK(clknet_leaf_12_clk),
    .D(_0217_),
    .Q(\mem[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1258_ (.CLK(clknet_leaf_7_clk),
    .D(_0218_),
    .Q(\mem[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1259_ (.CLK(clknet_leaf_8_clk),
    .D(_0219_),
    .Q(\mem[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1260_ (.CLK(clknet_leaf_8_clk),
    .D(_0220_),
    .Q(\mem[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1261_ (.CLK(clknet_leaf_27_clk),
    .D(_0221_),
    .Q(\mem[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1262_ (.CLK(clknet_leaf_26_clk),
    .D(_0222_),
    .Q(\mem[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1263_ (.CLK(clknet_leaf_25_clk),
    .D(_0223_),
    .Q(\mem[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1264_ (.CLK(clknet_leaf_20_clk),
    .D(_0224_),
    .Q(\mem[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1265_ (.CLK(clknet_leaf_24_clk),
    .D(_0225_),
    .Q(\mem[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1266_ (.CLK(clknet_leaf_18_clk),
    .D(_0226_),
    .Q(\mem[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1267_ (.CLK(clknet_leaf_3_clk),
    .D(_0227_),
    .Q(\mem[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1268_ (.CLK(clknet_leaf_17_clk),
    .D(_0228_),
    .Q(\mem[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1269_ (.CLK(clknet_leaf_2_clk),
    .D(_0229_),
    .Q(\mem[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1270_ (.CLK(clknet_leaf_15_clk),
    .D(_0230_),
    .Q(\mem[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1271_ (.CLK(clknet_leaf_11_clk),
    .D(_0231_),
    .Q(\mem[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1272_ (.CLK(clknet_leaf_11_clk),
    .D(_0232_),
    .Q(\mem[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1273_ (.CLK(clknet_leaf_12_clk),
    .D(_0233_),
    .Q(\mem[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1274_ (.CLK(clknet_leaf_9_clk),
    .D(_0234_),
    .Q(\mem[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1275_ (.CLK(clknet_leaf_12_clk),
    .D(_0235_),
    .Q(\mem[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1276_ (.CLK(clknet_leaf_7_clk),
    .D(_0236_),
    .Q(\mem[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1277_ (.CLK(clknet_leaf_27_clk),
    .D(_0237_),
    .Q(\mem[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1278_ (.CLK(clknet_leaf_27_clk),
    .D(_0238_),
    .Q(\mem[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1279_ (.CLK(clknet_leaf_24_clk),
    .D(_0239_),
    .Q(\mem[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1280_ (.CLK(clknet_leaf_23_clk),
    .D(_0240_),
    .Q(\mem[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1281_ (.CLK(clknet_leaf_0_clk),
    .D(_0241_),
    .Q(\mem[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1282_ (.CLK(clknet_leaf_23_clk),
    .D(_0242_),
    .Q(\mem[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1283_ (.CLK(clknet_leaf_3_clk),
    .D(_0243_),
    .Q(\mem[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1284_ (.CLK(clknet_leaf_16_clk),
    .D(_0244_),
    .Q(\mem[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1285_ (.CLK(clknet_leaf_3_clk),
    .D(_0245_),
    .Q(\mem[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1286_ (.CLK(clknet_leaf_11_clk),
    .D(_0246_),
    .Q(\mem[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1287_ (.CLK(clknet_leaf_8_clk),
    .D(_0247_),
    .Q(\mem[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1288_ (.CLK(clknet_leaf_5_clk),
    .D(_0248_),
    .Q(\mem[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1289_ (.CLK(clknet_leaf_12_clk),
    .D(_0249_),
    .Q(\mem[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1290_ (.CLK(clknet_leaf_5_clk),
    .D(_0250_),
    .Q(\mem[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1291_ (.CLK(clknet_leaf_8_clk),
    .D(_0251_),
    .Q(\mem[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1292_ (.CLK(clknet_leaf_5_clk),
    .D(_0252_),
    .Q(\mem[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1293_ (.CLK(clknet_leaf_28_clk),
    .D(_0253_),
    .Q(\mem[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1294_ (.CLK(clknet_leaf_23_clk),
    .D(_0254_),
    .Q(\mem[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1295_ (.CLK(clknet_leaf_28_clk),
    .D(_0255_),
    .Q(\mem[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1296_ (.CLK(clknet_leaf_20_clk),
    .D(_0256_),
    .Q(\mem[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1297_ (.CLK(clknet_leaf_2_clk),
    .D(_0257_),
    .Q(\mem[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1298_ (.CLK(clknet_leaf_18_clk),
    .D(_0258_),
    .Q(\mem[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1299_ (.CLK(clknet_leaf_1_clk),
    .D(_0259_),
    .Q(\mem[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1300_ (.CLK(clknet_leaf_16_clk),
    .D(_0260_),
    .Q(\mem[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1301_ (.CLK(clknet_leaf_4_clk),
    .D(_0261_),
    .Q(\mem[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1302_ (.CLK(clknet_leaf_11_clk),
    .D(_0262_),
    .Q(\mem[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1303_ (.CLK(clknet_leaf_9_clk),
    .D(_0263_),
    .Q(\mem[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1304_ (.CLK(clknet_leaf_4_clk),
    .D(_0264_),
    .Q(\mem[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1305_ (.CLK(clknet_leaf_12_clk),
    .D(_0265_),
    .Q(\mem[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1306_ (.CLK(clknet_leaf_5_clk),
    .D(_0266_),
    .Q(\mem[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1307_ (.CLK(clknet_leaf_13_clk),
    .D(_0267_),
    .Q(\mem[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1308_ (.CLK(clknet_leaf_7_clk),
    .D(_0268_),
    .Q(\mem[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _1309_ (.CLK(clknet_leaf_28_clk),
    .D(_0269_),
    .Q(\mem[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1310_ (.CLK(clknet_leaf_26_clk),
    .D(_0270_),
    .Q(\mem[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1311_ (.CLK(clknet_leaf_24_clk),
    .D(_0271_),
    .Q(\mem[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1312_ (.CLK(clknet_leaf_23_clk),
    .D(_0272_),
    .Q(\mem[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1313_ (.CLK(clknet_leaf_0_clk),
    .D(_0273_),
    .Q(\mem[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1314_ (.CLK(clknet_leaf_17_clk),
    .D(_0274_),
    .Q(\mem[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1315_ (.CLK(clknet_leaf_1_clk),
    .D(_0275_),
    .Q(\mem[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1316_ (.CLK(clknet_leaf_2_clk),
    .D(_0276_),
    .Q(\mem[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1317_ (.CLK(clknet_leaf_4_clk),
    .D(_0277_),
    .Q(\mem[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _1318_ (.CLK(clknet_leaf_11_clk),
    .D(_0278_),
    .Q(\mem[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _1319_ (.CLK(clknet_leaf_10_clk),
    .D(_0279_),
    .Q(\mem[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _1320_ (.CLK(clknet_leaf_5_clk),
    .D(_0280_),
    .Q(\mem[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _1321_ (.CLK(clknet_leaf_11_clk),
    .D(_0281_),
    .Q(\mem[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _1322_ (.CLK(clknet_leaf_7_clk),
    .D(_0282_),
    .Q(\mem[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _1323_ (.CLK(clknet_leaf_12_clk),
    .D(_0283_),
    .Q(\mem[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _1324_ (.CLK(clknet_leaf_7_clk),
    .D(_0284_),
    .Q(\mem[15][15] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_539 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(rd_en_i),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(rst_n),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(wr_data_i[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(wr_data_i[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(wr_data_i[11]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(wr_data_i[12]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(wr_data_i[13]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(wr_data_i[14]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(wr_data_i[15]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(wr_data_i[1]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(wr_data_i[2]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(wr_data_i[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(wr_data_i[4]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(wr_data_i[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(wr_data_i[6]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(wr_data_i[7]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(wr_data_i[8]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(wr_data_i[9]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(wr_en_i),
    .X(net19));
 sky130_fd_sc_hd__buf_4 output20 (.A(net20),
    .X(empty_o));
 sky130_fd_sc_hd__buf_4 output21 (.A(net21),
    .X(full_o));
 sky130_fd_sc_hd__buf_4 output22 (.A(net22),
    .X(rd_data_o[0]));
 sky130_fd_sc_hd__buf_4 output23 (.A(net23),
    .X(rd_data_o[10]));
 sky130_fd_sc_hd__buf_4 output24 (.A(net24),
    .X(rd_data_o[11]));
 sky130_fd_sc_hd__buf_4 output25 (.A(net25),
    .X(rd_data_o[12]));
 sky130_fd_sc_hd__buf_4 output26 (.A(net26),
    .X(rd_data_o[13]));
 sky130_fd_sc_hd__buf_4 output27 (.A(net27),
    .X(rd_data_o[14]));
 sky130_fd_sc_hd__buf_4 output28 (.A(net28),
    .X(rd_data_o[15]));
 sky130_fd_sc_hd__buf_4 output29 (.A(net29),
    .X(rd_data_o[1]));
 sky130_fd_sc_hd__buf_4 output30 (.A(net30),
    .X(rd_data_o[2]));
 sky130_fd_sc_hd__buf_4 output31 (.A(net31),
    .X(rd_data_o[3]));
 sky130_fd_sc_hd__buf_4 output32 (.A(net32),
    .X(rd_data_o[4]));
 sky130_fd_sc_hd__buf_4 output33 (.A(net33),
    .X(rd_data_o[5]));
 sky130_fd_sc_hd__buf_4 output34 (.A(net34),
    .X(rd_data_o[6]));
 sky130_fd_sc_hd__buf_4 output35 (.A(net35),
    .X(rd_data_o[7]));
 sky130_fd_sc_hd__buf_4 output36 (.A(net36),
    .X(rd_data_o[8]));
 sky130_fd_sc_hd__buf_4 output37 (.A(net37),
    .X(rd_data_o[9]));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(net40),
    .X(net38));
 sky130_fd_sc_hd__buf_2 fanout39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__buf_2 fanout40 (.A(_0291_),
    .X(net40));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(net44),
    .X(net41));
 sky130_fd_sc_hd__buf_1 fanout42 (.A(net44),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(_0290_),
    .X(net44));
 sky130_fd_sc_hd__buf_2 fanout45 (.A(net47),
    .X(net45));
 sky130_fd_sc_hd__buf_2 fanout46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(_0289_),
    .X(net47));
 sky130_fd_sc_hd__buf_2 fanout48 (.A(net51),
    .X(net48));
 sky130_fd_sc_hd__buf_2 fanout49 (.A(net51),
    .X(net49));
 sky130_fd_sc_hd__buf_1 fanout50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 fanout51 (.A(_0288_),
    .X(net51));
 sky130_fd_sc_hd__buf_2 fanout52 (.A(net54),
    .X(net52));
 sky130_fd_sc_hd__buf_2 fanout53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__buf_2 fanout54 (.A(_0286_),
    .X(net54));
 sky130_fd_sc_hd__buf_2 fanout55 (.A(net57),
    .X(net55));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout56 (.A(net57),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 fanout57 (.A(_0285_),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 fanout58 (.A(_0518_),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 fanout59 (.A(_0518_),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 fanout60 (.A(_0518_),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 fanout61 (.A(net63),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(_0517_),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 fanout64 (.A(net66),
    .X(net64));
 sky130_fd_sc_hd__buf_2 fanout65 (.A(net66),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 fanout66 (.A(_0515_),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 fanout67 (.A(net69),
    .X(net67));
 sky130_fd_sc_hd__buf_2 fanout68 (.A(net69),
    .X(net68));
 sky130_fd_sc_hd__buf_4 fanout69 (.A(_0514_),
    .X(net69));
 sky130_fd_sc_hd__buf_2 fanout70 (.A(net73),
    .X(net70));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout71 (.A(net73),
    .X(net71));
 sky130_fd_sc_hd__buf_2 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 fanout73 (.A(_0513_),
    .X(net73));
 sky130_fd_sc_hd__buf_2 fanout74 (.A(net77),
    .X(net74));
 sky130_fd_sc_hd__buf_2 fanout75 (.A(net77),
    .X(net75));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout77 (.A(_0512_),
    .X(net77));
 sky130_fd_sc_hd__buf_2 fanout78 (.A(net80),
    .X(net78));
 sky130_fd_sc_hd__buf_2 fanout79 (.A(net80),
    .X(net79));
 sky130_fd_sc_hd__buf_2 fanout80 (.A(_0510_),
    .X(net80));
 sky130_fd_sc_hd__buf_2 fanout81 (.A(_0509_),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 fanout82 (.A(_0509_),
    .X(net82));
 sky130_fd_sc_hd__buf_2 fanout83 (.A(_0509_),
    .X(net83));
 sky130_fd_sc_hd__buf_2 fanout84 (.A(net86),
    .X(net84));
 sky130_fd_sc_hd__buf_2 fanout85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__buf_2 fanout86 (.A(_0507_),
    .X(net86));
 sky130_fd_sc_hd__buf_2 fanout87 (.A(net90),
    .X(net87));
 sky130_fd_sc_hd__buf_2 fanout88 (.A(net90),
    .X(net88));
 sky130_fd_sc_hd__buf_1 fanout89 (.A(net90),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 fanout90 (.A(_0505_),
    .X(net90));
 sky130_fd_sc_hd__buf_2 fanout91 (.A(net94),
    .X(net91));
 sky130_fd_sc_hd__buf_2 fanout92 (.A(net94),
    .X(net92));
 sky130_fd_sc_hd__buf_1 fanout93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout94 (.A(_0334_),
    .X(net94));
 sky130_fd_sc_hd__buf_2 fanout95 (.A(net98),
    .X(net95));
 sky130_fd_sc_hd__buf_1 fanout96 (.A(net98),
    .X(net96));
 sky130_fd_sc_hd__buf_2 fanout97 (.A(net98),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 fanout98 (.A(_0333_),
    .X(net98));
 sky130_fd_sc_hd__buf_2 fanout99 (.A(net102),
    .X(net99));
 sky130_fd_sc_hd__buf_1 fanout100 (.A(net102),
    .X(net100));
 sky130_fd_sc_hd__buf_2 fanout101 (.A(net102),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 fanout102 (.A(_0332_),
    .X(net102));
 sky130_fd_sc_hd__buf_2 fanout103 (.A(net105),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 fanout105 (.A(_0330_),
    .X(net105));
 sky130_fd_sc_hd__buf_2 fanout106 (.A(net109),
    .X(net106));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout107 (.A(net109),
    .X(net107));
 sky130_fd_sc_hd__buf_2 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 fanout109 (.A(_0329_),
    .X(net109));
 sky130_fd_sc_hd__buf_2 fanout110 (.A(net113),
    .X(net110));
 sky130_fd_sc_hd__buf_2 fanout111 (.A(net113),
    .X(net111));
 sky130_fd_sc_hd__buf_1 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout113 (.A(_0328_),
    .X(net113));
 sky130_fd_sc_hd__buf_2 fanout114 (.A(net116),
    .X(net114));
 sky130_fd_sc_hd__buf_2 fanout115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 fanout116 (.A(_0326_),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 fanout117 (.A(net119),
    .X(net117));
 sky130_fd_sc_hd__buf_2 fanout118 (.A(net119),
    .X(net118));
 sky130_fd_sc_hd__buf_2 fanout119 (.A(_0318_),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 fanout120 (.A(_0299_),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 fanout121 (.A(net125),
    .X(net121));
 sky130_fd_sc_hd__buf_1 fanout122 (.A(net125),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 fanout123 (.A(net125),
    .X(net123));
 sky130_fd_sc_hd__buf_1 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 fanout125 (.A(_0297_),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 fanout126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 fanout127 (.A(net130),
    .X(net127));
 sky130_fd_sc_hd__buf_2 fanout128 (.A(net130),
    .X(net128));
 sky130_fd_sc_hd__buf_1 fanout129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 fanout130 (.A(_0296_),
    .X(net130));
 sky130_fd_sc_hd__buf_2 fanout131 (.A(net133),
    .X(net131));
 sky130_fd_sc_hd__buf_2 fanout132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__buf_2 fanout133 (.A(_0335_),
    .X(net133));
 sky130_fd_sc_hd__buf_2 fanout134 (.A(net136),
    .X(net134));
 sky130_fd_sc_hd__buf_2 fanout135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 fanout136 (.A(_0331_),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 fanout137 (.A(net139),
    .X(net137));
 sky130_fd_sc_hd__buf_1 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__buf_2 fanout139 (.A(_0325_),
    .X(net139));
 sky130_fd_sc_hd__buf_2 fanout140 (.A(net142),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_2 fanout141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__buf_2 fanout142 (.A(_0324_),
    .X(net142));
 sky130_fd_sc_hd__buf_2 fanout143 (.A(net146),
    .X(net143));
 sky130_fd_sc_hd__buf_2 fanout144 (.A(net146),
    .X(net144));
 sky130_fd_sc_hd__buf_1 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 fanout146 (.A(_0323_),
    .X(net146));
 sky130_fd_sc_hd__buf_2 fanout147 (.A(net150),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 fanout148 (.A(net150),
    .X(net148));
 sky130_fd_sc_hd__buf_2 fanout149 (.A(net150),
    .X(net149));
 sky130_fd_sc_hd__buf_2 fanout150 (.A(_0322_),
    .X(net150));
 sky130_fd_sc_hd__buf_2 fanout151 (.A(net153),
    .X(net151));
 sky130_fd_sc_hd__buf_2 fanout152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 fanout153 (.A(_0321_),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 fanout154 (.A(net156),
    .X(net154));
 sky130_fd_sc_hd__buf_2 fanout155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__buf_2 fanout156 (.A(_0320_),
    .X(net156));
 sky130_fd_sc_hd__buf_2 fanout157 (.A(net159),
    .X(net157));
 sky130_fd_sc_hd__buf_2 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__buf_2 fanout159 (.A(_0319_),
    .X(net159));
 sky130_fd_sc_hd__buf_1 fanout160 (.A(_0294_),
    .X(net160));
 sky130_fd_sc_hd__buf_1 fanout161 (.A(\wr_ptr[1] ),
    .X(net161));
 sky130_fd_sc_hd__buf_1 fanout162 (.A(\wr_ptr[1] ),
    .X(net162));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout163 (.A(\wr_ptr[0] ),
    .X(net163));
 sky130_fd_sc_hd__buf_1 fanout164 (.A(\wr_ptr[0] ),
    .X(net164));
 sky130_fd_sc_hd__buf_1 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout166 (.A(\rd_ptr[3] ),
    .X(net166));
 sky130_fd_sc_hd__buf_1 fanout167 (.A(net170),
    .X(net167));
 sky130_fd_sc_hd__buf_1 fanout168 (.A(net170),
    .X(net168));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__buf_1 fanout170 (.A(\rd_ptr[2] ),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__buf_1 fanout172 (.A(net174),
    .X(net172));
 sky130_fd_sc_hd__buf_1 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__buf_1 fanout174 (.A(\rd_ptr[1] ),
    .X(net174));
 sky130_fd_sc_hd__buf_1 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__buf_1 fanout176 (.A(net178),
    .X(net176));
 sky130_fd_sc_hd__buf_1 fanout177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 fanout178 (.A(\rd_ptr[0] ),
    .X(net178));
 sky130_fd_sc_hd__buf_1 fanout179 (.A(net181),
    .X(net179));
 sky130_fd_sc_hd__buf_1 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout181 (.A(net9),
    .X(net181));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout182 (.A(net184),
    .X(net182));
 sky130_fd_sc_hd__buf_1 fanout183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__buf_1 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 fanout185 (.A(net8),
    .X(net185));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout186 (.A(net189),
    .X(net186));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout187 (.A(net189),
    .X(net187));
 sky130_fd_sc_hd__buf_1 fanout188 (.A(net189),
    .X(net188));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout189 (.A(net7),
    .X(net189));
 sky130_fd_sc_hd__buf_1 fanout190 (.A(net192),
    .X(net190));
 sky130_fd_sc_hd__buf_1 fanout191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout192 (.A(net6),
    .X(net192));
 sky130_fd_sc_hd__buf_1 fanout193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 fanout195 (.A(net5),
    .X(net195));
 sky130_fd_sc_hd__buf_1 fanout196 (.A(net198),
    .X(net196));
 sky130_fd_sc_hd__buf_1 fanout197 (.A(net198),
    .X(net197));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__buf_1 fanout199 (.A(net4),
    .X(net199));
 sky130_fd_sc_hd__buf_1 fanout200 (.A(net202),
    .X(net200));
 sky130_fd_sc_hd__buf_1 fanout201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 fanout202 (.A(net3),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 fanout203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout204 (.A(net206),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_2 fanout205 (.A(net206),
    .X(net205));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout206 (.A(net208),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 fanout207 (.A(net208),
    .X(net207));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout208 (.A(net211),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 fanout209 (.A(net211),
    .X(net209));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 fanout211 (.A(net2),
    .X(net211));
 sky130_fd_sc_hd__buf_1 fanout212 (.A(net214),
    .X(net212));
 sky130_fd_sc_hd__buf_1 fanout213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout214 (.A(net18),
    .X(net214));
 sky130_fd_sc_hd__buf_1 fanout215 (.A(net218),
    .X(net215));
 sky130_fd_sc_hd__buf_1 fanout216 (.A(net218),
    .X(net216));
 sky130_fd_sc_hd__buf_1 fanout217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__buf_1 fanout218 (.A(net17),
    .X(net218));
 sky130_fd_sc_hd__buf_1 fanout219 (.A(net221),
    .X(net219));
 sky130_fd_sc_hd__buf_1 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout221 (.A(net16),
    .X(net221));
 sky130_fd_sc_hd__buf_1 fanout222 (.A(net225),
    .X(net222));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout223 (.A(net225),
    .X(net223));
 sky130_fd_sc_hd__buf_1 fanout224 (.A(net225),
    .X(net224));
 sky130_fd_sc_hd__buf_1 fanout225 (.A(net15),
    .X(net225));
 sky130_fd_sc_hd__buf_1 fanout226 (.A(net229),
    .X(net226));
 sky130_fd_sc_hd__buf_1 fanout227 (.A(net229),
    .X(net227));
 sky130_fd_sc_hd__buf_1 fanout228 (.A(net229),
    .X(net228));
 sky130_fd_sc_hd__buf_1 fanout229 (.A(net14),
    .X(net229));
 sky130_fd_sc_hd__buf_1 fanout230 (.A(net233),
    .X(net230));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout231 (.A(net233),
    .X(net231));
 sky130_fd_sc_hd__buf_1 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__buf_1 fanout233 (.A(net13),
    .X(net233));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout234 (.A(net237),
    .X(net234));
 sky130_fd_sc_hd__buf_1 fanout235 (.A(net237),
    .X(net235));
 sky130_fd_sc_hd__buf_1 fanout236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__buf_1 fanout237 (.A(net12),
    .X(net237));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout238 (.A(net11),
    .X(net238));
 sky130_fd_sc_hd__buf_1 fanout239 (.A(net11),
    .X(net239));
 sky130_fd_sc_hd__buf_1 fanout240 (.A(net11),
    .X(net240));
 sky130_fd_sc_hd__buf_1 fanout241 (.A(net10),
    .X(net241));
 sky130_fd_sc_hd__buf_1 fanout242 (.A(net243),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_2 fanout243 (.A(net10),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload1 (.A(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload3 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__inv_6 clkload4 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload5 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__inv_6 clkload6 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__inv_8 clkload7 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkinv_2 clkload8 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload9 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkinv_2 clkload10 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload11 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkinv_2 clkload12 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__inv_6 clkload13 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkinv_2 clkload14 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload15 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__bufinv_16 clkload16 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__bufinv_16 clkload17 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload18 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkinv_4 clkload19 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__inv_4 clkload20 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__inv_6 clkload21 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkinv_4 clkload22 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload23 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload24 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__inv_6 clkload25 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__inv_6 clkload26 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__inv_8 clkload27 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_A (.DIODE(_0285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0943__S (.DIODE(_0285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0950__S (.DIODE(_0285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0937__Y (.DIODE(_0285_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(_0325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0702__A2 (.DIODE(_0325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0627__A2 (.DIODE(_0325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0559__X (.DIODE(_0325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0624__B1 (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0623__X (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(_0509_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(_0509_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(_0509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0799__Y (.DIODE(_0509_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_A (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_A (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0920__Y (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(rd_en_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(rst_n));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(wr_data_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(wr_data_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(wr_data_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(wr_data_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(wr_data_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(wr_data_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(wr_data_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(wr_data_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(wr_data_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(wr_data_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(wr_data_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(wr_data_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(wr_data_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(wr_data_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(wr_data_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(wr_data_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(wr_en_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_X (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__0544__A2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__0526__B1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__0525__B1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_X (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__0950__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__0945__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__0911__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__0982__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__0947__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_X (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__0528__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__0527__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout38_X (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1026__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1029__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1024__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1028__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1025__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout39_X (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__1034__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__1032__S (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout40_X (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1038__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1036__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout39_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1027__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__S (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout38_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout41_X (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1015__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1017__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1011__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1009__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1007__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1013__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout43_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1014__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1019__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1021__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1012__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1010__S (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout44_X (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__1016__S (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout43_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout41_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout42_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout45_X (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__1005__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__1001__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__1003__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__0994__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__0991__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__0990__S (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout46_X (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__1002__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__1004__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__0997__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__0995__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__0992__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__0993__S (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_X (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__1000__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__0999__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout46_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__S (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout45_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_X (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__0976__S (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__0980__S (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__S (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__0974__S (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__0973__S (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__0977__S (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout49_X (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__0987__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__0986__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__0988__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__0983__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__0979__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_X (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout49_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__S (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_X (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__0960__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__0961__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__0957__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__0956__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__0955__S (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_X (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__0964__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__0963__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__0970__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__0968__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__0966__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__0965__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_X (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__0967__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__0969__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__0958__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__0962__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_X (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__0952__S (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__0945__S (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__0947__S (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__0941__S (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_X (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__0930__S (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__0928__S (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__0934__S (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__0936__S (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__0929__S (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__0927__S (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_X (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__0926__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__0924__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__0925__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__0923__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__0921__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__0922__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_X (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__0906__S (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__0911__S (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__0910__S (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__0908__S (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__0905__S (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__0904__S (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_X (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__0916__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__0912__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__0917__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__0915__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__0914__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__0919__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_X (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__0913__S (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__0918__S (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__0909__S (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__0907__S (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_X (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__0887__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__0893__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__0892__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__0890__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__0888__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__0886__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_X (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__0898__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__0896__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__0894__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__0901__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__0899__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__0897__S (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_X (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__0895__S (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__0900__S (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__0891__S (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__0889__S (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout67_X (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__0884__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__0875__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__0871__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__0870__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__0869__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__0881__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__0880__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__0874__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__0876__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__0872__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_X (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__0879__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__0883__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__0877__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__0882__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout67_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_X (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0859__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0860__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0856__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0854__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0852__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_X (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0866__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0862__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0867__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0865__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__0861__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_X (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0838__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0839__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0837__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0836__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0835__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__0841__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_X (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0844__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0848__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0846__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0845__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__0843__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__0840__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0821__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0823__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0820__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0819__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0817__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__0818__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0832__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0830__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0826__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0827__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0825__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__0828__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_X (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0831__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0829__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0824__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__0822__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_X (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0807__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0813__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0811__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0808__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0815__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__0806__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_X (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0801__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0805__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0800__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0803__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0804__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__0802__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0789__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0788__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0784__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0783__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__0782__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_X (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0791__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0797__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0795__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0793__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0792__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__0790__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_X (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0796__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0794__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0787__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__0785__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_X (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0770__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0768__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0766__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0765__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__0764__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_X (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0773__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0777__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0774__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__0772__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_X (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__0769__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_X (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0603__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0584__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0574__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0640__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0615__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__0592__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_X (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0648__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0715__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0695__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0662__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__0741__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_X (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0605__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0584__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0642__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0621__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0596__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__0575__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_X (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0706__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0740__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0697__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0687__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__0658__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0672__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__0726__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_X (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0648__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0660__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0614__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0597__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0573__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__0637__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_X (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__0728__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__0681__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__0735__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_X (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__0702__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_X (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0629__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0638__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0593__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0586__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0575__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__0617__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_X (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0724__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0707__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0714__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0659__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0742__A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__0686__A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_X (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0691__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0672__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0652__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__0610__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_X (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0680__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0736__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0641__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0620__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0585__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__0576__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_X (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0659__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0720__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__0696__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_X (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0705__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0632__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0606__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0595__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0649__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_X (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__0731__A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_X (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0605__A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0621__A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0599__A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0588__A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0571__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__0637__A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_X (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0714__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0738__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0680__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__0665__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_X (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__0632__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_X (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0738__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0643__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0598__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0585__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0576__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__0617__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_X (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0691__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0630__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0651__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__0606__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_X (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0724__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0708__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0662__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__0718__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_X (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0625__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0636__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0618__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0596__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0574__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__0587__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_X (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0671__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0684__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0716__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0694__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0736__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__0658__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_X (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0706__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0654__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__0609__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_X (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_X (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0623__C1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0645__C1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0590__C1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0579__C1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__0601__C1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__C1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0656__C1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0744__C1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0722__C1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__C1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__0667__C1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_X (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0634__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__0752__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_X (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0719__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0638__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0695__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0615__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0582__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0570__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0703__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0728__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0651__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0627__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0604__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__0595__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0686__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0676__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0664__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__0739__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__0604__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__0593__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__0639__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__0577__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__0619__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__0583__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0676__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0682__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0737__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0715__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0693__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0661__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_X (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0727__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0705__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0631__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0725__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0647__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0669__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__0608__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_X (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__0626__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__0641__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__0618__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__0594__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__0583__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__0572__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_X (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__0735__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__0661__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__0718__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__0693__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__0708__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__0650__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__0603__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_X (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__0607__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__0639__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__0594__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__0571__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__0616__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__0587__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_X (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__0730__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__0739__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__0660__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__0628__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_X (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__0663__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__0616__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__0597__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__0572__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__0636__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_X (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__0650__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__0709__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__0725__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__0581__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__0629__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__0609__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_X (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__0656__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__0601__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__0590__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__0579__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__0645__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__0623__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_X (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__0711__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__0667__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__0744__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__0722__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_X (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__0700__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__0634__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__0612__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_X (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__0610__D1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__0643__C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__0622__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__0599__C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__0588__C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__0577__C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_X (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__0671__C1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__0742__C1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__0716__C1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__0694__C1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__0687__C1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__0665__C1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_X (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__0731__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__0709__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__0626__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__0654__B1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_X (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__0607__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__0642__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__0620__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__0598__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__0573__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__0586__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_X (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__0703__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__0741__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__0716__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__0694__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__0684__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__0664__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_X (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__0727__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__0671__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__0625__B1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__0652__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_X (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__0984__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__0932__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__0880__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__0775__A0 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_X (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__1064__RESET_B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_X (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_X (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__0991__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__0974__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__0939__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__0905__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__0870__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload0_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload1_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload2_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net139));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_5 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_5 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_365 ();
endmodule
