magic
tech sky130A
magscale 1 2
timestamp 1769196144
<< viali >>
rect 28089 27421 28123 27455
rect 28365 27353 28399 27387
rect 28089 25857 28123 25891
rect 28365 25789 28399 25823
rect 27721 24361 27755 24395
rect 27537 24157 27571 24191
rect 28089 24157 28123 24191
rect 28365 24089 28399 24123
rect 27721 22729 27755 22763
rect 1501 22593 1535 22627
rect 27537 22593 27571 22627
rect 28089 22593 28123 22627
rect 28365 22525 28399 22559
rect 1777 22389 1811 22423
rect 27721 22185 27755 22219
rect 27537 21981 27571 22015
rect 28089 20893 28123 20927
rect 28365 20825 28399 20859
rect 28089 19329 28123 19363
rect 28365 19329 28399 19363
rect 27721 18921 27755 18955
rect 27537 18717 27571 18751
rect 27721 18377 27755 18411
rect 27537 18241 27571 18275
rect 28089 17629 28123 17663
rect 28365 17561 28399 17595
rect 27445 17289 27479 17323
rect 26985 17085 27019 17119
rect 27353 17017 27387 17051
rect 27537 17017 27571 17051
rect 27353 16745 27387 16779
rect 27169 16677 27203 16711
rect 26893 16609 26927 16643
rect 28089 16201 28123 16235
rect 27261 16065 27295 16099
rect 27169 15997 27203 16031
rect 28365 15521 28399 15555
rect 28089 15453 28123 15487
rect 28089 14365 28123 14399
rect 28365 14297 28399 14331
rect 27721 13481 27755 13515
rect 27537 13277 27571 13311
rect 27077 12801 27111 12835
rect 27169 12801 27203 12835
rect 28089 12801 28123 12835
rect 28365 12733 28399 12767
rect 27353 12597 27387 12631
rect 27721 11849 27755 11883
rect 27537 11713 27571 11747
rect 28089 11101 28123 11135
rect 28365 11033 28399 11067
rect 27813 10693 27847 10727
rect 26617 10625 26651 10659
rect 26801 10625 26835 10659
rect 27077 10625 27111 10659
rect 26801 10489 26835 10523
rect 27537 9537 27571 9571
rect 28089 9537 28123 9571
rect 28365 9469 28399 9503
rect 27721 9401 27755 9435
rect 27721 9129 27755 9163
rect 27537 8925 27571 8959
rect 28089 7837 28123 7871
rect 1501 7769 1535 7803
rect 28365 7769 28399 7803
rect 1777 7701 1811 7735
rect 28089 6273 28123 6307
rect 28365 6205 28399 6239
rect 27721 5865 27755 5899
rect 27537 5661 27571 5695
rect 28089 4573 28123 4607
rect 28365 4505 28399 4539
rect 28089 3009 28123 3043
rect 28365 2941 28399 2975
<< metal1 >>
rect 1104 27770 28888 27792
rect 1104 27718 1950 27770
rect 2002 27718 2014 27770
rect 2066 27718 2078 27770
rect 2130 27718 2142 27770
rect 2194 27718 2206 27770
rect 2258 27718 9950 27770
rect 10002 27718 10014 27770
rect 10066 27718 10078 27770
rect 10130 27718 10142 27770
rect 10194 27718 10206 27770
rect 10258 27718 17950 27770
rect 18002 27718 18014 27770
rect 18066 27718 18078 27770
rect 18130 27718 18142 27770
rect 18194 27718 18206 27770
rect 18258 27718 25950 27770
rect 26002 27718 26014 27770
rect 26066 27718 26078 27770
rect 26130 27718 26142 27770
rect 26194 27718 26206 27770
rect 26258 27718 28888 27770
rect 1104 27696 28888 27718
rect 27614 27412 27620 27464
rect 27672 27452 27678 27464
rect 28077 27455 28135 27461
rect 28077 27452 28089 27455
rect 27672 27424 28089 27452
rect 27672 27412 27678 27424
rect 28077 27421 28089 27424
rect 28123 27421 28135 27455
rect 28077 27415 28135 27421
rect 28350 27344 28356 27396
rect 28408 27344 28414 27396
rect 1104 27226 28888 27248
rect 1104 27174 2610 27226
rect 2662 27174 2674 27226
rect 2726 27174 2738 27226
rect 2790 27174 2802 27226
rect 2854 27174 2866 27226
rect 2918 27174 10610 27226
rect 10662 27174 10674 27226
rect 10726 27174 10738 27226
rect 10790 27174 10802 27226
rect 10854 27174 10866 27226
rect 10918 27174 18610 27226
rect 18662 27174 18674 27226
rect 18726 27174 18738 27226
rect 18790 27174 18802 27226
rect 18854 27174 18866 27226
rect 18918 27174 26610 27226
rect 26662 27174 26674 27226
rect 26726 27174 26738 27226
rect 26790 27174 26802 27226
rect 26854 27174 26866 27226
rect 26918 27174 28888 27226
rect 1104 27152 28888 27174
rect 1104 26682 28888 26704
rect 1104 26630 1950 26682
rect 2002 26630 2014 26682
rect 2066 26630 2078 26682
rect 2130 26630 2142 26682
rect 2194 26630 2206 26682
rect 2258 26630 9950 26682
rect 10002 26630 10014 26682
rect 10066 26630 10078 26682
rect 10130 26630 10142 26682
rect 10194 26630 10206 26682
rect 10258 26630 17950 26682
rect 18002 26630 18014 26682
rect 18066 26630 18078 26682
rect 18130 26630 18142 26682
rect 18194 26630 18206 26682
rect 18258 26630 25950 26682
rect 26002 26630 26014 26682
rect 26066 26630 26078 26682
rect 26130 26630 26142 26682
rect 26194 26630 26206 26682
rect 26258 26630 28888 26682
rect 1104 26608 28888 26630
rect 1104 26138 28888 26160
rect 1104 26086 2610 26138
rect 2662 26086 2674 26138
rect 2726 26086 2738 26138
rect 2790 26086 2802 26138
rect 2854 26086 2866 26138
rect 2918 26086 10610 26138
rect 10662 26086 10674 26138
rect 10726 26086 10738 26138
rect 10790 26086 10802 26138
rect 10854 26086 10866 26138
rect 10918 26086 18610 26138
rect 18662 26086 18674 26138
rect 18726 26086 18738 26138
rect 18790 26086 18802 26138
rect 18854 26086 18866 26138
rect 18918 26086 26610 26138
rect 26662 26086 26674 26138
rect 26726 26086 26738 26138
rect 26790 26086 26802 26138
rect 26854 26086 26866 26138
rect 26918 26086 28888 26138
rect 1104 26064 28888 26086
rect 28074 25848 28080 25900
rect 28132 25848 28138 25900
rect 28350 25780 28356 25832
rect 28408 25780 28414 25832
rect 1104 25594 28888 25616
rect 1104 25542 1950 25594
rect 2002 25542 2014 25594
rect 2066 25542 2078 25594
rect 2130 25542 2142 25594
rect 2194 25542 2206 25594
rect 2258 25542 9950 25594
rect 10002 25542 10014 25594
rect 10066 25542 10078 25594
rect 10130 25542 10142 25594
rect 10194 25542 10206 25594
rect 10258 25542 17950 25594
rect 18002 25542 18014 25594
rect 18066 25542 18078 25594
rect 18130 25542 18142 25594
rect 18194 25542 18206 25594
rect 18258 25542 25950 25594
rect 26002 25542 26014 25594
rect 26066 25542 26078 25594
rect 26130 25542 26142 25594
rect 26194 25542 26206 25594
rect 26258 25542 28888 25594
rect 1104 25520 28888 25542
rect 1104 25050 28888 25072
rect 1104 24998 2610 25050
rect 2662 24998 2674 25050
rect 2726 24998 2738 25050
rect 2790 24998 2802 25050
rect 2854 24998 2866 25050
rect 2918 24998 10610 25050
rect 10662 24998 10674 25050
rect 10726 24998 10738 25050
rect 10790 24998 10802 25050
rect 10854 24998 10866 25050
rect 10918 24998 18610 25050
rect 18662 24998 18674 25050
rect 18726 24998 18738 25050
rect 18790 24998 18802 25050
rect 18854 24998 18866 25050
rect 18918 24998 26610 25050
rect 26662 24998 26674 25050
rect 26726 24998 26738 25050
rect 26790 24998 26802 25050
rect 26854 24998 26866 25050
rect 26918 24998 28888 25050
rect 1104 24976 28888 24998
rect 1104 24506 28888 24528
rect 1104 24454 1950 24506
rect 2002 24454 2014 24506
rect 2066 24454 2078 24506
rect 2130 24454 2142 24506
rect 2194 24454 2206 24506
rect 2258 24454 9950 24506
rect 10002 24454 10014 24506
rect 10066 24454 10078 24506
rect 10130 24454 10142 24506
rect 10194 24454 10206 24506
rect 10258 24454 17950 24506
rect 18002 24454 18014 24506
rect 18066 24454 18078 24506
rect 18130 24454 18142 24506
rect 18194 24454 18206 24506
rect 18258 24454 25950 24506
rect 26002 24454 26014 24506
rect 26066 24454 26078 24506
rect 26130 24454 26142 24506
rect 26194 24454 26206 24506
rect 26258 24454 28888 24506
rect 1104 24432 28888 24454
rect 27709 24395 27767 24401
rect 27709 24361 27721 24395
rect 27755 24392 27767 24395
rect 28074 24392 28080 24404
rect 27755 24364 28080 24392
rect 27755 24361 27767 24364
rect 27709 24355 27767 24361
rect 28074 24352 28080 24364
rect 28132 24352 28138 24404
rect 27522 24148 27528 24200
rect 27580 24148 27586 24200
rect 28074 24148 28080 24200
rect 28132 24148 28138 24200
rect 28350 24080 28356 24132
rect 28408 24080 28414 24132
rect 1104 23962 28888 23984
rect 1104 23910 2610 23962
rect 2662 23910 2674 23962
rect 2726 23910 2738 23962
rect 2790 23910 2802 23962
rect 2854 23910 2866 23962
rect 2918 23910 10610 23962
rect 10662 23910 10674 23962
rect 10726 23910 10738 23962
rect 10790 23910 10802 23962
rect 10854 23910 10866 23962
rect 10918 23910 18610 23962
rect 18662 23910 18674 23962
rect 18726 23910 18738 23962
rect 18790 23910 18802 23962
rect 18854 23910 18866 23962
rect 18918 23910 26610 23962
rect 26662 23910 26674 23962
rect 26726 23910 26738 23962
rect 26790 23910 26802 23962
rect 26854 23910 26866 23962
rect 26918 23910 28888 23962
rect 1104 23888 28888 23910
rect 1104 23418 28888 23440
rect 1104 23366 1950 23418
rect 2002 23366 2014 23418
rect 2066 23366 2078 23418
rect 2130 23366 2142 23418
rect 2194 23366 2206 23418
rect 2258 23366 9950 23418
rect 10002 23366 10014 23418
rect 10066 23366 10078 23418
rect 10130 23366 10142 23418
rect 10194 23366 10206 23418
rect 10258 23366 17950 23418
rect 18002 23366 18014 23418
rect 18066 23366 18078 23418
rect 18130 23366 18142 23418
rect 18194 23366 18206 23418
rect 18258 23366 25950 23418
rect 26002 23366 26014 23418
rect 26066 23366 26078 23418
rect 26130 23366 26142 23418
rect 26194 23366 26206 23418
rect 26258 23366 28888 23418
rect 1104 23344 28888 23366
rect 1104 22874 28888 22896
rect 1104 22822 2610 22874
rect 2662 22822 2674 22874
rect 2726 22822 2738 22874
rect 2790 22822 2802 22874
rect 2854 22822 2866 22874
rect 2918 22822 10610 22874
rect 10662 22822 10674 22874
rect 10726 22822 10738 22874
rect 10790 22822 10802 22874
rect 10854 22822 10866 22874
rect 10918 22822 18610 22874
rect 18662 22822 18674 22874
rect 18726 22822 18738 22874
rect 18790 22822 18802 22874
rect 18854 22822 18866 22874
rect 18918 22822 26610 22874
rect 26662 22822 26674 22874
rect 26726 22822 26738 22874
rect 26790 22822 26802 22874
rect 26854 22822 26866 22874
rect 26918 22822 28888 22874
rect 1104 22800 28888 22822
rect 27709 22763 27767 22769
rect 27709 22729 27721 22763
rect 27755 22760 27767 22763
rect 28074 22760 28080 22772
rect 27755 22732 28080 22760
rect 27755 22729 27767 22732
rect 27709 22723 27767 22729
rect 28074 22720 28080 22732
rect 28132 22720 28138 22772
rect 842 22584 848 22636
rect 900 22624 906 22636
rect 1489 22627 1547 22633
rect 1489 22624 1501 22627
rect 900 22596 1501 22624
rect 900 22584 906 22596
rect 1489 22593 1501 22596
rect 1535 22593 1547 22627
rect 1489 22587 1547 22593
rect 27430 22584 27436 22636
rect 27488 22624 27494 22636
rect 27525 22627 27583 22633
rect 27525 22624 27537 22627
rect 27488 22596 27537 22624
rect 27488 22584 27494 22596
rect 27525 22593 27537 22596
rect 27571 22593 27583 22627
rect 27525 22587 27583 22593
rect 28074 22584 28080 22636
rect 28132 22584 28138 22636
rect 28350 22516 28356 22568
rect 28408 22516 28414 22568
rect 1762 22380 1768 22432
rect 1820 22380 1826 22432
rect 1104 22330 28888 22352
rect 1104 22278 1950 22330
rect 2002 22278 2014 22330
rect 2066 22278 2078 22330
rect 2130 22278 2142 22330
rect 2194 22278 2206 22330
rect 2258 22278 9950 22330
rect 10002 22278 10014 22330
rect 10066 22278 10078 22330
rect 10130 22278 10142 22330
rect 10194 22278 10206 22330
rect 10258 22278 17950 22330
rect 18002 22278 18014 22330
rect 18066 22278 18078 22330
rect 18130 22278 18142 22330
rect 18194 22278 18206 22330
rect 18258 22278 25950 22330
rect 26002 22278 26014 22330
rect 26066 22278 26078 22330
rect 26130 22278 26142 22330
rect 26194 22278 26206 22330
rect 26258 22278 28888 22330
rect 1104 22256 28888 22278
rect 27709 22219 27767 22225
rect 27709 22185 27721 22219
rect 27755 22216 27767 22219
rect 28074 22216 28080 22228
rect 27755 22188 28080 22216
rect 27755 22185 27767 22188
rect 27709 22179 27767 22185
rect 28074 22176 28080 22188
rect 28132 22176 28138 22228
rect 27522 21972 27528 22024
rect 27580 21972 27586 22024
rect 1104 21786 28888 21808
rect 1104 21734 2610 21786
rect 2662 21734 2674 21786
rect 2726 21734 2738 21786
rect 2790 21734 2802 21786
rect 2854 21734 2866 21786
rect 2918 21734 10610 21786
rect 10662 21734 10674 21786
rect 10726 21734 10738 21786
rect 10790 21734 10802 21786
rect 10854 21734 10866 21786
rect 10918 21734 18610 21786
rect 18662 21734 18674 21786
rect 18726 21734 18738 21786
rect 18790 21734 18802 21786
rect 18854 21734 18866 21786
rect 18918 21734 26610 21786
rect 26662 21734 26674 21786
rect 26726 21734 26738 21786
rect 26790 21734 26802 21786
rect 26854 21734 26866 21786
rect 26918 21734 28888 21786
rect 1104 21712 28888 21734
rect 1104 21242 28888 21264
rect 1104 21190 1950 21242
rect 2002 21190 2014 21242
rect 2066 21190 2078 21242
rect 2130 21190 2142 21242
rect 2194 21190 2206 21242
rect 2258 21190 9950 21242
rect 10002 21190 10014 21242
rect 10066 21190 10078 21242
rect 10130 21190 10142 21242
rect 10194 21190 10206 21242
rect 10258 21190 17950 21242
rect 18002 21190 18014 21242
rect 18066 21190 18078 21242
rect 18130 21190 18142 21242
rect 18194 21190 18206 21242
rect 18258 21190 25950 21242
rect 26002 21190 26014 21242
rect 26066 21190 26078 21242
rect 26130 21190 26142 21242
rect 26194 21190 26206 21242
rect 26258 21190 28888 21242
rect 1104 21168 28888 21190
rect 27430 20884 27436 20936
rect 27488 20924 27494 20936
rect 28077 20927 28135 20933
rect 28077 20924 28089 20927
rect 27488 20896 28089 20924
rect 27488 20884 27494 20896
rect 28077 20893 28089 20896
rect 28123 20893 28135 20927
rect 28077 20887 28135 20893
rect 28350 20816 28356 20868
rect 28408 20816 28414 20868
rect 1104 20698 28888 20720
rect 1104 20646 2610 20698
rect 2662 20646 2674 20698
rect 2726 20646 2738 20698
rect 2790 20646 2802 20698
rect 2854 20646 2866 20698
rect 2918 20646 10610 20698
rect 10662 20646 10674 20698
rect 10726 20646 10738 20698
rect 10790 20646 10802 20698
rect 10854 20646 10866 20698
rect 10918 20646 18610 20698
rect 18662 20646 18674 20698
rect 18726 20646 18738 20698
rect 18790 20646 18802 20698
rect 18854 20646 18866 20698
rect 18918 20646 26610 20698
rect 26662 20646 26674 20698
rect 26726 20646 26738 20698
rect 26790 20646 26802 20698
rect 26854 20646 26866 20698
rect 26918 20646 28888 20698
rect 1104 20624 28888 20646
rect 1104 20154 28888 20176
rect 1104 20102 1950 20154
rect 2002 20102 2014 20154
rect 2066 20102 2078 20154
rect 2130 20102 2142 20154
rect 2194 20102 2206 20154
rect 2258 20102 9950 20154
rect 10002 20102 10014 20154
rect 10066 20102 10078 20154
rect 10130 20102 10142 20154
rect 10194 20102 10206 20154
rect 10258 20102 17950 20154
rect 18002 20102 18014 20154
rect 18066 20102 18078 20154
rect 18130 20102 18142 20154
rect 18194 20102 18206 20154
rect 18258 20102 25950 20154
rect 26002 20102 26014 20154
rect 26066 20102 26078 20154
rect 26130 20102 26142 20154
rect 26194 20102 26206 20154
rect 26258 20102 28888 20154
rect 1104 20080 28888 20102
rect 1104 19610 28888 19632
rect 1104 19558 2610 19610
rect 2662 19558 2674 19610
rect 2726 19558 2738 19610
rect 2790 19558 2802 19610
rect 2854 19558 2866 19610
rect 2918 19558 10610 19610
rect 10662 19558 10674 19610
rect 10726 19558 10738 19610
rect 10790 19558 10802 19610
rect 10854 19558 10866 19610
rect 10918 19558 18610 19610
rect 18662 19558 18674 19610
rect 18726 19558 18738 19610
rect 18790 19558 18802 19610
rect 18854 19558 18866 19610
rect 18918 19558 26610 19610
rect 26662 19558 26674 19610
rect 26726 19558 26738 19610
rect 26790 19558 26802 19610
rect 26854 19558 26866 19610
rect 26918 19558 28888 19610
rect 1104 19536 28888 19558
rect 28074 19320 28080 19372
rect 28132 19320 28138 19372
rect 28350 19320 28356 19372
rect 28408 19320 28414 19372
rect 1104 19066 28888 19088
rect 1104 19014 1950 19066
rect 2002 19014 2014 19066
rect 2066 19014 2078 19066
rect 2130 19014 2142 19066
rect 2194 19014 2206 19066
rect 2258 19014 9950 19066
rect 10002 19014 10014 19066
rect 10066 19014 10078 19066
rect 10130 19014 10142 19066
rect 10194 19014 10206 19066
rect 10258 19014 17950 19066
rect 18002 19014 18014 19066
rect 18066 19014 18078 19066
rect 18130 19014 18142 19066
rect 18194 19014 18206 19066
rect 18258 19014 25950 19066
rect 26002 19014 26014 19066
rect 26066 19014 26078 19066
rect 26130 19014 26142 19066
rect 26194 19014 26206 19066
rect 26258 19014 28888 19066
rect 1104 18992 28888 19014
rect 27709 18955 27767 18961
rect 27709 18921 27721 18955
rect 27755 18952 27767 18955
rect 28074 18952 28080 18964
rect 27755 18924 28080 18952
rect 27755 18921 27767 18924
rect 27709 18915 27767 18921
rect 28074 18912 28080 18924
rect 28132 18912 28138 18964
rect 27522 18708 27528 18760
rect 27580 18708 27586 18760
rect 1104 18522 28888 18544
rect 1104 18470 2610 18522
rect 2662 18470 2674 18522
rect 2726 18470 2738 18522
rect 2790 18470 2802 18522
rect 2854 18470 2866 18522
rect 2918 18470 10610 18522
rect 10662 18470 10674 18522
rect 10726 18470 10738 18522
rect 10790 18470 10802 18522
rect 10854 18470 10866 18522
rect 10918 18470 18610 18522
rect 18662 18470 18674 18522
rect 18726 18470 18738 18522
rect 18790 18470 18802 18522
rect 18854 18470 18866 18522
rect 18918 18470 26610 18522
rect 26662 18470 26674 18522
rect 26726 18470 26738 18522
rect 26790 18470 26802 18522
rect 26854 18470 26866 18522
rect 26918 18470 28888 18522
rect 1104 18448 28888 18470
rect 27614 18368 27620 18420
rect 27672 18408 27678 18420
rect 27709 18411 27767 18417
rect 27709 18408 27721 18411
rect 27672 18380 27721 18408
rect 27672 18368 27678 18380
rect 27709 18377 27721 18380
rect 27755 18377 27767 18411
rect 27709 18371 27767 18377
rect 27338 18232 27344 18284
rect 27396 18272 27402 18284
rect 27525 18275 27583 18281
rect 27525 18272 27537 18275
rect 27396 18244 27537 18272
rect 27396 18232 27402 18244
rect 27525 18241 27537 18244
rect 27571 18241 27583 18275
rect 27525 18235 27583 18241
rect 1104 17978 28888 18000
rect 1104 17926 1950 17978
rect 2002 17926 2014 17978
rect 2066 17926 2078 17978
rect 2130 17926 2142 17978
rect 2194 17926 2206 17978
rect 2258 17926 9950 17978
rect 10002 17926 10014 17978
rect 10066 17926 10078 17978
rect 10130 17926 10142 17978
rect 10194 17926 10206 17978
rect 10258 17926 17950 17978
rect 18002 17926 18014 17978
rect 18066 17926 18078 17978
rect 18130 17926 18142 17978
rect 18194 17926 18206 17978
rect 18258 17926 25950 17978
rect 26002 17926 26014 17978
rect 26066 17926 26078 17978
rect 26130 17926 26142 17978
rect 26194 17926 26206 17978
rect 26258 17926 28888 17978
rect 1104 17904 28888 17926
rect 27338 17620 27344 17672
rect 27396 17660 27402 17672
rect 28077 17663 28135 17669
rect 28077 17660 28089 17663
rect 27396 17632 28089 17660
rect 27396 17620 27402 17632
rect 28077 17629 28089 17632
rect 28123 17629 28135 17663
rect 28077 17623 28135 17629
rect 28350 17552 28356 17604
rect 28408 17552 28414 17604
rect 1104 17434 28888 17456
rect 1104 17382 2610 17434
rect 2662 17382 2674 17434
rect 2726 17382 2738 17434
rect 2790 17382 2802 17434
rect 2854 17382 2866 17434
rect 2918 17382 10610 17434
rect 10662 17382 10674 17434
rect 10726 17382 10738 17434
rect 10790 17382 10802 17434
rect 10854 17382 10866 17434
rect 10918 17382 18610 17434
rect 18662 17382 18674 17434
rect 18726 17382 18738 17434
rect 18790 17382 18802 17434
rect 18854 17382 18866 17434
rect 18918 17382 26610 17434
rect 26662 17382 26674 17434
rect 26726 17382 26738 17434
rect 26790 17382 26802 17434
rect 26854 17382 26866 17434
rect 26918 17382 28888 17434
rect 1104 17360 28888 17382
rect 27430 17280 27436 17332
rect 27488 17280 27494 17332
rect 26970 17076 26976 17128
rect 27028 17076 27034 17128
rect 26878 17048 26884 17060
rect 26206 17020 26884 17048
rect 1762 16940 1768 16992
rect 1820 16980 1826 16992
rect 26206 16980 26234 17020
rect 26878 17008 26884 17020
rect 26936 17048 26942 17060
rect 27341 17051 27399 17057
rect 27341 17048 27353 17051
rect 26936 17020 27353 17048
rect 26936 17008 26942 17020
rect 27341 17017 27353 17020
rect 27387 17048 27399 17051
rect 27525 17051 27583 17057
rect 27525 17048 27537 17051
rect 27387 17020 27537 17048
rect 27387 17017 27399 17020
rect 27341 17011 27399 17017
rect 27525 17017 27537 17020
rect 27571 17017 27583 17051
rect 27525 17011 27583 17017
rect 1820 16952 26234 16980
rect 1820 16940 1826 16952
rect 1104 16890 28888 16912
rect 1104 16838 1950 16890
rect 2002 16838 2014 16890
rect 2066 16838 2078 16890
rect 2130 16838 2142 16890
rect 2194 16838 2206 16890
rect 2258 16838 9950 16890
rect 10002 16838 10014 16890
rect 10066 16838 10078 16890
rect 10130 16838 10142 16890
rect 10194 16838 10206 16890
rect 10258 16838 17950 16890
rect 18002 16838 18014 16890
rect 18066 16838 18078 16890
rect 18130 16838 18142 16890
rect 18194 16838 18206 16890
rect 18258 16838 25950 16890
rect 26002 16838 26014 16890
rect 26066 16838 26078 16890
rect 26130 16838 26142 16890
rect 26194 16838 26206 16890
rect 26258 16838 28888 16890
rect 1104 16816 28888 16838
rect 27338 16736 27344 16788
rect 27396 16736 27402 16788
rect 26970 16668 26976 16720
rect 27028 16708 27034 16720
rect 27157 16711 27215 16717
rect 27157 16708 27169 16711
rect 27028 16680 27169 16708
rect 27028 16668 27034 16680
rect 27157 16677 27169 16680
rect 27203 16677 27215 16711
rect 27157 16671 27215 16677
rect 26878 16600 26884 16652
rect 26936 16640 26942 16652
rect 27062 16640 27068 16652
rect 26936 16612 27068 16640
rect 26936 16600 26942 16612
rect 27062 16600 27068 16612
rect 27120 16600 27126 16652
rect 1104 16346 28888 16368
rect 1104 16294 2610 16346
rect 2662 16294 2674 16346
rect 2726 16294 2738 16346
rect 2790 16294 2802 16346
rect 2854 16294 2866 16346
rect 2918 16294 10610 16346
rect 10662 16294 10674 16346
rect 10726 16294 10738 16346
rect 10790 16294 10802 16346
rect 10854 16294 10866 16346
rect 10918 16294 18610 16346
rect 18662 16294 18674 16346
rect 18726 16294 18738 16346
rect 18790 16294 18802 16346
rect 18854 16294 18866 16346
rect 18918 16294 26610 16346
rect 26662 16294 26674 16346
rect 26726 16294 26738 16346
rect 26790 16294 26802 16346
rect 26854 16294 26866 16346
rect 26918 16294 28888 16346
rect 1104 16272 28888 16294
rect 27522 16192 27528 16244
rect 27580 16232 27586 16244
rect 28077 16235 28135 16241
rect 28077 16232 28089 16235
rect 27580 16204 28089 16232
rect 27580 16192 27586 16204
rect 28077 16201 28089 16204
rect 28123 16201 28135 16235
rect 28077 16195 28135 16201
rect 27062 16056 27068 16108
rect 27120 16096 27126 16108
rect 27249 16099 27307 16105
rect 27249 16096 27261 16099
rect 27120 16068 27261 16096
rect 27120 16056 27126 16068
rect 27249 16065 27261 16068
rect 27295 16065 27307 16099
rect 27249 16059 27307 16065
rect 27154 15988 27160 16040
rect 27212 15988 27218 16040
rect 1104 15802 28888 15824
rect 1104 15750 1950 15802
rect 2002 15750 2014 15802
rect 2066 15750 2078 15802
rect 2130 15750 2142 15802
rect 2194 15750 2206 15802
rect 2258 15750 9950 15802
rect 10002 15750 10014 15802
rect 10066 15750 10078 15802
rect 10130 15750 10142 15802
rect 10194 15750 10206 15802
rect 10258 15750 17950 15802
rect 18002 15750 18014 15802
rect 18066 15750 18078 15802
rect 18130 15750 18142 15802
rect 18194 15750 18206 15802
rect 18258 15750 25950 15802
rect 26002 15750 26014 15802
rect 26066 15750 26078 15802
rect 26130 15750 26142 15802
rect 26194 15750 26206 15802
rect 26258 15750 28888 15802
rect 1104 15728 28888 15750
rect 28350 15512 28356 15564
rect 28408 15512 28414 15564
rect 27522 15444 27528 15496
rect 27580 15484 27586 15496
rect 28077 15487 28135 15493
rect 28077 15484 28089 15487
rect 27580 15456 28089 15484
rect 27580 15444 27586 15456
rect 28077 15453 28089 15456
rect 28123 15453 28135 15487
rect 28077 15447 28135 15453
rect 1104 15258 28888 15280
rect 1104 15206 2610 15258
rect 2662 15206 2674 15258
rect 2726 15206 2738 15258
rect 2790 15206 2802 15258
rect 2854 15206 2866 15258
rect 2918 15206 10610 15258
rect 10662 15206 10674 15258
rect 10726 15206 10738 15258
rect 10790 15206 10802 15258
rect 10854 15206 10866 15258
rect 10918 15206 18610 15258
rect 18662 15206 18674 15258
rect 18726 15206 18738 15258
rect 18790 15206 18802 15258
rect 18854 15206 18866 15258
rect 18918 15206 26610 15258
rect 26662 15206 26674 15258
rect 26726 15206 26738 15258
rect 26790 15206 26802 15258
rect 26854 15206 26866 15258
rect 26918 15206 28888 15258
rect 1104 15184 28888 15206
rect 1104 14714 28888 14736
rect 1104 14662 1950 14714
rect 2002 14662 2014 14714
rect 2066 14662 2078 14714
rect 2130 14662 2142 14714
rect 2194 14662 2206 14714
rect 2258 14662 9950 14714
rect 10002 14662 10014 14714
rect 10066 14662 10078 14714
rect 10130 14662 10142 14714
rect 10194 14662 10206 14714
rect 10258 14662 17950 14714
rect 18002 14662 18014 14714
rect 18066 14662 18078 14714
rect 18130 14662 18142 14714
rect 18194 14662 18206 14714
rect 18258 14662 25950 14714
rect 26002 14662 26014 14714
rect 26066 14662 26078 14714
rect 26130 14662 26142 14714
rect 26194 14662 26206 14714
rect 26258 14662 28888 14714
rect 1104 14640 28888 14662
rect 28074 14356 28080 14408
rect 28132 14356 28138 14408
rect 28350 14288 28356 14340
rect 28408 14288 28414 14340
rect 1104 14170 28888 14192
rect 1104 14118 2610 14170
rect 2662 14118 2674 14170
rect 2726 14118 2738 14170
rect 2790 14118 2802 14170
rect 2854 14118 2866 14170
rect 2918 14118 10610 14170
rect 10662 14118 10674 14170
rect 10726 14118 10738 14170
rect 10790 14118 10802 14170
rect 10854 14118 10866 14170
rect 10918 14118 18610 14170
rect 18662 14118 18674 14170
rect 18726 14118 18738 14170
rect 18790 14118 18802 14170
rect 18854 14118 18866 14170
rect 18918 14118 26610 14170
rect 26662 14118 26674 14170
rect 26726 14118 26738 14170
rect 26790 14118 26802 14170
rect 26854 14118 26866 14170
rect 26918 14118 28888 14170
rect 1104 14096 28888 14118
rect 1104 13626 28888 13648
rect 1104 13574 1950 13626
rect 2002 13574 2014 13626
rect 2066 13574 2078 13626
rect 2130 13574 2142 13626
rect 2194 13574 2206 13626
rect 2258 13574 9950 13626
rect 10002 13574 10014 13626
rect 10066 13574 10078 13626
rect 10130 13574 10142 13626
rect 10194 13574 10206 13626
rect 10258 13574 17950 13626
rect 18002 13574 18014 13626
rect 18066 13574 18078 13626
rect 18130 13574 18142 13626
rect 18194 13574 18206 13626
rect 18258 13574 25950 13626
rect 26002 13574 26014 13626
rect 26066 13574 26078 13626
rect 26130 13574 26142 13626
rect 26194 13574 26206 13626
rect 26258 13574 28888 13626
rect 1104 13552 28888 13574
rect 27709 13515 27767 13521
rect 27709 13481 27721 13515
rect 27755 13512 27767 13515
rect 28074 13512 28080 13524
rect 27755 13484 28080 13512
rect 27755 13481 27767 13484
rect 27709 13475 27767 13481
rect 28074 13472 28080 13484
rect 28132 13472 28138 13524
rect 27525 13311 27583 13317
rect 27525 13277 27537 13311
rect 27571 13308 27583 13311
rect 27614 13308 27620 13320
rect 27571 13280 27620 13308
rect 27571 13277 27583 13280
rect 27525 13271 27583 13277
rect 27614 13268 27620 13280
rect 27672 13268 27678 13320
rect 1104 13082 28888 13104
rect 1104 13030 2610 13082
rect 2662 13030 2674 13082
rect 2726 13030 2738 13082
rect 2790 13030 2802 13082
rect 2854 13030 2866 13082
rect 2918 13030 10610 13082
rect 10662 13030 10674 13082
rect 10726 13030 10738 13082
rect 10790 13030 10802 13082
rect 10854 13030 10866 13082
rect 10918 13030 18610 13082
rect 18662 13030 18674 13082
rect 18726 13030 18738 13082
rect 18790 13030 18802 13082
rect 18854 13030 18866 13082
rect 18918 13030 26610 13082
rect 26662 13030 26674 13082
rect 26726 13030 26738 13082
rect 26790 13030 26802 13082
rect 26854 13030 26866 13082
rect 26918 13030 28888 13082
rect 1104 13008 28888 13030
rect 27062 12792 27068 12844
rect 27120 12792 27126 12844
rect 27154 12792 27160 12844
rect 27212 12792 27218 12844
rect 28074 12792 28080 12844
rect 28132 12792 28138 12844
rect 28350 12724 28356 12776
rect 28408 12724 28414 12776
rect 27341 12631 27399 12637
rect 27341 12597 27353 12631
rect 27387 12628 27399 12631
rect 27614 12628 27620 12640
rect 27387 12600 27620 12628
rect 27387 12597 27399 12600
rect 27341 12591 27399 12597
rect 27614 12588 27620 12600
rect 27672 12628 27678 12640
rect 28166 12628 28172 12640
rect 27672 12600 28172 12628
rect 27672 12588 27678 12600
rect 28166 12588 28172 12600
rect 28224 12588 28230 12640
rect 1104 12538 28888 12560
rect 1104 12486 1950 12538
rect 2002 12486 2014 12538
rect 2066 12486 2078 12538
rect 2130 12486 2142 12538
rect 2194 12486 2206 12538
rect 2258 12486 9950 12538
rect 10002 12486 10014 12538
rect 10066 12486 10078 12538
rect 10130 12486 10142 12538
rect 10194 12486 10206 12538
rect 10258 12486 17950 12538
rect 18002 12486 18014 12538
rect 18066 12486 18078 12538
rect 18130 12486 18142 12538
rect 18194 12486 18206 12538
rect 18258 12486 25950 12538
rect 26002 12486 26014 12538
rect 26066 12486 26078 12538
rect 26130 12486 26142 12538
rect 26194 12486 26206 12538
rect 26258 12486 28888 12538
rect 1104 12464 28888 12486
rect 1104 11994 28888 12016
rect 1104 11942 2610 11994
rect 2662 11942 2674 11994
rect 2726 11942 2738 11994
rect 2790 11942 2802 11994
rect 2854 11942 2866 11994
rect 2918 11942 10610 11994
rect 10662 11942 10674 11994
rect 10726 11942 10738 11994
rect 10790 11942 10802 11994
rect 10854 11942 10866 11994
rect 10918 11942 18610 11994
rect 18662 11942 18674 11994
rect 18726 11942 18738 11994
rect 18790 11942 18802 11994
rect 18854 11942 18866 11994
rect 18918 11942 26610 11994
rect 26662 11942 26674 11994
rect 26726 11942 26738 11994
rect 26790 11942 26802 11994
rect 26854 11942 26866 11994
rect 26918 11942 28888 11994
rect 1104 11920 28888 11942
rect 27709 11883 27767 11889
rect 27709 11849 27721 11883
rect 27755 11880 27767 11883
rect 28074 11880 28080 11892
rect 27755 11852 28080 11880
rect 27755 11849 27767 11852
rect 27709 11843 27767 11849
rect 28074 11840 28080 11852
rect 28132 11840 28138 11892
rect 27430 11704 27436 11756
rect 27488 11744 27494 11756
rect 27525 11747 27583 11753
rect 27525 11744 27537 11747
rect 27488 11716 27537 11744
rect 27488 11704 27494 11716
rect 27525 11713 27537 11716
rect 27571 11713 27583 11747
rect 27525 11707 27583 11713
rect 1104 11450 28888 11472
rect 1104 11398 1950 11450
rect 2002 11398 2014 11450
rect 2066 11398 2078 11450
rect 2130 11398 2142 11450
rect 2194 11398 2206 11450
rect 2258 11398 9950 11450
rect 10002 11398 10014 11450
rect 10066 11398 10078 11450
rect 10130 11398 10142 11450
rect 10194 11398 10206 11450
rect 10258 11398 17950 11450
rect 18002 11398 18014 11450
rect 18066 11398 18078 11450
rect 18130 11398 18142 11450
rect 18194 11398 18206 11450
rect 18258 11398 25950 11450
rect 26002 11398 26014 11450
rect 26066 11398 26078 11450
rect 26130 11398 26142 11450
rect 26194 11398 26206 11450
rect 26258 11398 28888 11450
rect 1104 11376 28888 11398
rect 28074 11092 28080 11144
rect 28132 11092 28138 11144
rect 28350 11024 28356 11076
rect 28408 11024 28414 11076
rect 1104 10906 28888 10928
rect 1104 10854 2610 10906
rect 2662 10854 2674 10906
rect 2726 10854 2738 10906
rect 2790 10854 2802 10906
rect 2854 10854 2866 10906
rect 2918 10854 10610 10906
rect 10662 10854 10674 10906
rect 10726 10854 10738 10906
rect 10790 10854 10802 10906
rect 10854 10854 10866 10906
rect 10918 10854 18610 10906
rect 18662 10854 18674 10906
rect 18726 10854 18738 10906
rect 18790 10854 18802 10906
rect 18854 10854 18866 10906
rect 18918 10854 26610 10906
rect 26662 10854 26674 10906
rect 26726 10854 26738 10906
rect 26790 10854 26802 10906
rect 26854 10854 26866 10906
rect 26918 10854 28888 10906
rect 1104 10832 28888 10854
rect 27246 10792 27252 10804
rect 26804 10764 27252 10792
rect 26510 10616 26516 10668
rect 26568 10656 26574 10668
rect 26804 10665 26832 10764
rect 27246 10752 27252 10764
rect 27304 10752 27310 10804
rect 27430 10684 27436 10736
rect 27488 10724 27494 10736
rect 27801 10727 27859 10733
rect 27801 10724 27813 10727
rect 27488 10696 27813 10724
rect 27488 10684 27494 10696
rect 27801 10693 27813 10696
rect 27847 10693 27859 10727
rect 27801 10687 27859 10693
rect 26605 10659 26663 10665
rect 26605 10656 26617 10659
rect 26568 10628 26617 10656
rect 26568 10616 26574 10628
rect 26605 10625 26617 10628
rect 26651 10625 26663 10659
rect 26605 10619 26663 10625
rect 26789 10659 26847 10665
rect 26789 10625 26801 10659
rect 26835 10625 26847 10659
rect 26789 10619 26847 10625
rect 26620 10588 26648 10619
rect 27062 10616 27068 10668
rect 27120 10616 27126 10668
rect 27246 10616 27252 10668
rect 27304 10616 27310 10668
rect 27080 10588 27108 10616
rect 26620 10560 27108 10588
rect 26789 10523 26847 10529
rect 26789 10489 26801 10523
rect 26835 10520 26847 10523
rect 27522 10520 27528 10532
rect 26835 10492 27528 10520
rect 26835 10489 26847 10492
rect 26789 10483 26847 10489
rect 27522 10480 27528 10492
rect 27580 10480 27586 10532
rect 1104 10362 28888 10384
rect 1104 10310 1950 10362
rect 2002 10310 2014 10362
rect 2066 10310 2078 10362
rect 2130 10310 2142 10362
rect 2194 10310 2206 10362
rect 2258 10310 9950 10362
rect 10002 10310 10014 10362
rect 10066 10310 10078 10362
rect 10130 10310 10142 10362
rect 10194 10310 10206 10362
rect 10258 10310 17950 10362
rect 18002 10310 18014 10362
rect 18066 10310 18078 10362
rect 18130 10310 18142 10362
rect 18194 10310 18206 10362
rect 18258 10310 25950 10362
rect 26002 10310 26014 10362
rect 26066 10310 26078 10362
rect 26130 10310 26142 10362
rect 26194 10310 26206 10362
rect 26258 10310 28888 10362
rect 1104 10288 28888 10310
rect 1104 9818 28888 9840
rect 1104 9766 2610 9818
rect 2662 9766 2674 9818
rect 2726 9766 2738 9818
rect 2790 9766 2802 9818
rect 2854 9766 2866 9818
rect 2918 9766 10610 9818
rect 10662 9766 10674 9818
rect 10726 9766 10738 9818
rect 10790 9766 10802 9818
rect 10854 9766 10866 9818
rect 10918 9766 18610 9818
rect 18662 9766 18674 9818
rect 18726 9766 18738 9818
rect 18790 9766 18802 9818
rect 18854 9766 18866 9818
rect 18918 9766 26610 9818
rect 26662 9766 26674 9818
rect 26726 9766 26738 9818
rect 26790 9766 26802 9818
rect 26854 9766 26866 9818
rect 26918 9766 28888 9818
rect 1104 9744 28888 9766
rect 27522 9528 27528 9580
rect 27580 9528 27586 9580
rect 27706 9528 27712 9580
rect 27764 9568 27770 9580
rect 28077 9571 28135 9577
rect 28077 9568 28089 9571
rect 27764 9540 28089 9568
rect 27764 9528 27770 9540
rect 28077 9537 28089 9540
rect 28123 9537 28135 9571
rect 28077 9531 28135 9537
rect 28350 9460 28356 9512
rect 28408 9460 28414 9512
rect 27709 9435 27767 9441
rect 27709 9401 27721 9435
rect 27755 9432 27767 9435
rect 28074 9432 28080 9444
rect 27755 9404 28080 9432
rect 27755 9401 27767 9404
rect 27709 9395 27767 9401
rect 28074 9392 28080 9404
rect 28132 9392 28138 9444
rect 1104 9274 28888 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 9950 9274
rect 10002 9222 10014 9274
rect 10066 9222 10078 9274
rect 10130 9222 10142 9274
rect 10194 9222 10206 9274
rect 10258 9222 17950 9274
rect 18002 9222 18014 9274
rect 18066 9222 18078 9274
rect 18130 9222 18142 9274
rect 18194 9222 18206 9274
rect 18258 9222 25950 9274
rect 26002 9222 26014 9274
rect 26066 9222 26078 9274
rect 26130 9222 26142 9274
rect 26194 9222 26206 9274
rect 26258 9222 28888 9274
rect 1104 9200 28888 9222
rect 27706 9120 27712 9172
rect 27764 9120 27770 9172
rect 27430 8916 27436 8968
rect 27488 8956 27494 8968
rect 27525 8959 27583 8965
rect 27525 8956 27537 8959
rect 27488 8928 27537 8956
rect 27488 8916 27494 8928
rect 27525 8925 27537 8928
rect 27571 8925 27583 8959
rect 27525 8919 27583 8925
rect 1104 8730 28888 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 10610 8730
rect 10662 8678 10674 8730
rect 10726 8678 10738 8730
rect 10790 8678 10802 8730
rect 10854 8678 10866 8730
rect 10918 8678 18610 8730
rect 18662 8678 18674 8730
rect 18726 8678 18738 8730
rect 18790 8678 18802 8730
rect 18854 8678 18866 8730
rect 18918 8678 26610 8730
rect 26662 8678 26674 8730
rect 26726 8678 26738 8730
rect 26790 8678 26802 8730
rect 26854 8678 26866 8730
rect 26918 8678 28888 8730
rect 1104 8656 28888 8678
rect 1104 8186 28888 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 9950 8186
rect 10002 8134 10014 8186
rect 10066 8134 10078 8186
rect 10130 8134 10142 8186
rect 10194 8134 10206 8186
rect 10258 8134 17950 8186
rect 18002 8134 18014 8186
rect 18066 8134 18078 8186
rect 18130 8134 18142 8186
rect 18194 8134 18206 8186
rect 18258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 28888 8186
rect 1104 8112 28888 8134
rect 27522 7828 27528 7880
rect 27580 7868 27586 7880
rect 28077 7871 28135 7877
rect 28077 7868 28089 7871
rect 27580 7840 28089 7868
rect 27580 7828 27586 7840
rect 28077 7837 28089 7840
rect 28123 7837 28135 7871
rect 28077 7831 28135 7837
rect 842 7760 848 7812
rect 900 7800 906 7812
rect 1489 7803 1547 7809
rect 1489 7800 1501 7803
rect 900 7772 1501 7800
rect 900 7760 906 7772
rect 1489 7769 1501 7772
rect 1535 7769 1547 7803
rect 1489 7763 1547 7769
rect 28350 7760 28356 7812
rect 28408 7760 28414 7812
rect 1765 7735 1823 7741
rect 1765 7701 1777 7735
rect 1811 7732 1823 7735
rect 26510 7732 26516 7744
rect 1811 7704 26516 7732
rect 1811 7701 1823 7704
rect 1765 7695 1823 7701
rect 26510 7692 26516 7704
rect 26568 7692 26574 7744
rect 1104 7642 28888 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 10610 7642
rect 10662 7590 10674 7642
rect 10726 7590 10738 7642
rect 10790 7590 10802 7642
rect 10854 7590 10866 7642
rect 10918 7590 18610 7642
rect 18662 7590 18674 7642
rect 18726 7590 18738 7642
rect 18790 7590 18802 7642
rect 18854 7590 18866 7642
rect 18918 7590 26610 7642
rect 26662 7590 26674 7642
rect 26726 7590 26738 7642
rect 26790 7590 26802 7642
rect 26854 7590 26866 7642
rect 26918 7590 28888 7642
rect 1104 7568 28888 7590
rect 1104 7098 28888 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 9950 7098
rect 10002 7046 10014 7098
rect 10066 7046 10078 7098
rect 10130 7046 10142 7098
rect 10194 7046 10206 7098
rect 10258 7046 17950 7098
rect 18002 7046 18014 7098
rect 18066 7046 18078 7098
rect 18130 7046 18142 7098
rect 18194 7046 18206 7098
rect 18258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 28888 7098
rect 1104 7024 28888 7046
rect 1104 6554 28888 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 10610 6554
rect 10662 6502 10674 6554
rect 10726 6502 10738 6554
rect 10790 6502 10802 6554
rect 10854 6502 10866 6554
rect 10918 6502 18610 6554
rect 18662 6502 18674 6554
rect 18726 6502 18738 6554
rect 18790 6502 18802 6554
rect 18854 6502 18866 6554
rect 18918 6502 26610 6554
rect 26662 6502 26674 6554
rect 26726 6502 26738 6554
rect 26790 6502 26802 6554
rect 26854 6502 26866 6554
rect 26918 6502 28888 6554
rect 1104 6480 28888 6502
rect 27706 6264 27712 6316
rect 27764 6304 27770 6316
rect 28077 6307 28135 6313
rect 28077 6304 28089 6307
rect 27764 6276 28089 6304
rect 27764 6264 27770 6276
rect 28077 6273 28089 6276
rect 28123 6273 28135 6307
rect 28077 6267 28135 6273
rect 28350 6196 28356 6248
rect 28408 6196 28414 6248
rect 1104 6010 28888 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 9950 6010
rect 10002 5958 10014 6010
rect 10066 5958 10078 6010
rect 10130 5958 10142 6010
rect 10194 5958 10206 6010
rect 10258 5958 17950 6010
rect 18002 5958 18014 6010
rect 18066 5958 18078 6010
rect 18130 5958 18142 6010
rect 18194 5958 18206 6010
rect 18258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 28888 6010
rect 1104 5936 28888 5958
rect 27706 5856 27712 5908
rect 27764 5856 27770 5908
rect 27522 5652 27528 5704
rect 27580 5652 27586 5704
rect 1104 5466 28888 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 10610 5466
rect 10662 5414 10674 5466
rect 10726 5414 10738 5466
rect 10790 5414 10802 5466
rect 10854 5414 10866 5466
rect 10918 5414 18610 5466
rect 18662 5414 18674 5466
rect 18726 5414 18738 5466
rect 18790 5414 18802 5466
rect 18854 5414 18866 5466
rect 18918 5414 26610 5466
rect 26662 5414 26674 5466
rect 26726 5414 26738 5466
rect 26790 5414 26802 5466
rect 26854 5414 26866 5466
rect 26918 5414 28888 5466
rect 1104 5392 28888 5414
rect 1104 4922 28888 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 9950 4922
rect 10002 4870 10014 4922
rect 10066 4870 10078 4922
rect 10130 4870 10142 4922
rect 10194 4870 10206 4922
rect 10258 4870 17950 4922
rect 18002 4870 18014 4922
rect 18066 4870 18078 4922
rect 18130 4870 18142 4922
rect 18194 4870 18206 4922
rect 18258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 28888 4922
rect 1104 4848 28888 4870
rect 28077 4607 28135 4613
rect 28077 4573 28089 4607
rect 28123 4604 28135 4607
rect 28166 4604 28172 4616
rect 28123 4576 28172 4604
rect 28123 4573 28135 4576
rect 28077 4567 28135 4573
rect 28166 4564 28172 4576
rect 28224 4564 28230 4616
rect 28350 4496 28356 4548
rect 28408 4496 28414 4548
rect 1104 4378 28888 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 10610 4378
rect 10662 4326 10674 4378
rect 10726 4326 10738 4378
rect 10790 4326 10802 4378
rect 10854 4326 10866 4378
rect 10918 4326 18610 4378
rect 18662 4326 18674 4378
rect 18726 4326 18738 4378
rect 18790 4326 18802 4378
rect 18854 4326 18866 4378
rect 18918 4326 26610 4378
rect 26662 4326 26674 4378
rect 26726 4326 26738 4378
rect 26790 4326 26802 4378
rect 26854 4326 26866 4378
rect 26918 4326 28888 4378
rect 1104 4304 28888 4326
rect 1104 3834 28888 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 9950 3834
rect 10002 3782 10014 3834
rect 10066 3782 10078 3834
rect 10130 3782 10142 3834
rect 10194 3782 10206 3834
rect 10258 3782 17950 3834
rect 18002 3782 18014 3834
rect 18066 3782 18078 3834
rect 18130 3782 18142 3834
rect 18194 3782 18206 3834
rect 18258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 28888 3834
rect 1104 3760 28888 3782
rect 1104 3290 28888 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 10610 3290
rect 10662 3238 10674 3290
rect 10726 3238 10738 3290
rect 10790 3238 10802 3290
rect 10854 3238 10866 3290
rect 10918 3238 18610 3290
rect 18662 3238 18674 3290
rect 18726 3238 18738 3290
rect 18790 3238 18802 3290
rect 18854 3238 18866 3290
rect 18918 3238 26610 3290
rect 26662 3238 26674 3290
rect 26726 3238 26738 3290
rect 26790 3238 26802 3290
rect 26854 3238 26866 3290
rect 26918 3238 28888 3290
rect 1104 3216 28888 3238
rect 27522 3000 27528 3052
rect 27580 3040 27586 3052
rect 28077 3043 28135 3049
rect 28077 3040 28089 3043
rect 27580 3012 28089 3040
rect 27580 3000 27586 3012
rect 28077 3009 28089 3012
rect 28123 3009 28135 3043
rect 28077 3003 28135 3009
rect 28350 2932 28356 2984
rect 28408 2932 28414 2984
rect 1104 2746 28888 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 9950 2746
rect 10002 2694 10014 2746
rect 10066 2694 10078 2746
rect 10130 2694 10142 2746
rect 10194 2694 10206 2746
rect 10258 2694 17950 2746
rect 18002 2694 18014 2746
rect 18066 2694 18078 2746
rect 18130 2694 18142 2746
rect 18194 2694 18206 2746
rect 18258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 28888 2746
rect 1104 2672 28888 2694
rect 1104 2202 28888 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 10610 2202
rect 10662 2150 10674 2202
rect 10726 2150 10738 2202
rect 10790 2150 10802 2202
rect 10854 2150 10866 2202
rect 10918 2150 18610 2202
rect 18662 2150 18674 2202
rect 18726 2150 18738 2202
rect 18790 2150 18802 2202
rect 18854 2150 18866 2202
rect 18918 2150 26610 2202
rect 26662 2150 26674 2202
rect 26726 2150 26738 2202
rect 26790 2150 26802 2202
rect 26854 2150 26866 2202
rect 26918 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 1950 27718 2002 27770
rect 2014 27718 2066 27770
rect 2078 27718 2130 27770
rect 2142 27718 2194 27770
rect 2206 27718 2258 27770
rect 9950 27718 10002 27770
rect 10014 27718 10066 27770
rect 10078 27718 10130 27770
rect 10142 27718 10194 27770
rect 10206 27718 10258 27770
rect 17950 27718 18002 27770
rect 18014 27718 18066 27770
rect 18078 27718 18130 27770
rect 18142 27718 18194 27770
rect 18206 27718 18258 27770
rect 25950 27718 26002 27770
rect 26014 27718 26066 27770
rect 26078 27718 26130 27770
rect 26142 27718 26194 27770
rect 26206 27718 26258 27770
rect 27620 27412 27672 27464
rect 28356 27387 28408 27396
rect 28356 27353 28365 27387
rect 28365 27353 28399 27387
rect 28399 27353 28408 27387
rect 28356 27344 28408 27353
rect 2610 27174 2662 27226
rect 2674 27174 2726 27226
rect 2738 27174 2790 27226
rect 2802 27174 2854 27226
rect 2866 27174 2918 27226
rect 10610 27174 10662 27226
rect 10674 27174 10726 27226
rect 10738 27174 10790 27226
rect 10802 27174 10854 27226
rect 10866 27174 10918 27226
rect 18610 27174 18662 27226
rect 18674 27174 18726 27226
rect 18738 27174 18790 27226
rect 18802 27174 18854 27226
rect 18866 27174 18918 27226
rect 26610 27174 26662 27226
rect 26674 27174 26726 27226
rect 26738 27174 26790 27226
rect 26802 27174 26854 27226
rect 26866 27174 26918 27226
rect 1950 26630 2002 26682
rect 2014 26630 2066 26682
rect 2078 26630 2130 26682
rect 2142 26630 2194 26682
rect 2206 26630 2258 26682
rect 9950 26630 10002 26682
rect 10014 26630 10066 26682
rect 10078 26630 10130 26682
rect 10142 26630 10194 26682
rect 10206 26630 10258 26682
rect 17950 26630 18002 26682
rect 18014 26630 18066 26682
rect 18078 26630 18130 26682
rect 18142 26630 18194 26682
rect 18206 26630 18258 26682
rect 25950 26630 26002 26682
rect 26014 26630 26066 26682
rect 26078 26630 26130 26682
rect 26142 26630 26194 26682
rect 26206 26630 26258 26682
rect 2610 26086 2662 26138
rect 2674 26086 2726 26138
rect 2738 26086 2790 26138
rect 2802 26086 2854 26138
rect 2866 26086 2918 26138
rect 10610 26086 10662 26138
rect 10674 26086 10726 26138
rect 10738 26086 10790 26138
rect 10802 26086 10854 26138
rect 10866 26086 10918 26138
rect 18610 26086 18662 26138
rect 18674 26086 18726 26138
rect 18738 26086 18790 26138
rect 18802 26086 18854 26138
rect 18866 26086 18918 26138
rect 26610 26086 26662 26138
rect 26674 26086 26726 26138
rect 26738 26086 26790 26138
rect 26802 26086 26854 26138
rect 26866 26086 26918 26138
rect 28080 25891 28132 25900
rect 28080 25857 28089 25891
rect 28089 25857 28123 25891
rect 28123 25857 28132 25891
rect 28080 25848 28132 25857
rect 28356 25823 28408 25832
rect 28356 25789 28365 25823
rect 28365 25789 28399 25823
rect 28399 25789 28408 25823
rect 28356 25780 28408 25789
rect 1950 25542 2002 25594
rect 2014 25542 2066 25594
rect 2078 25542 2130 25594
rect 2142 25542 2194 25594
rect 2206 25542 2258 25594
rect 9950 25542 10002 25594
rect 10014 25542 10066 25594
rect 10078 25542 10130 25594
rect 10142 25542 10194 25594
rect 10206 25542 10258 25594
rect 17950 25542 18002 25594
rect 18014 25542 18066 25594
rect 18078 25542 18130 25594
rect 18142 25542 18194 25594
rect 18206 25542 18258 25594
rect 25950 25542 26002 25594
rect 26014 25542 26066 25594
rect 26078 25542 26130 25594
rect 26142 25542 26194 25594
rect 26206 25542 26258 25594
rect 2610 24998 2662 25050
rect 2674 24998 2726 25050
rect 2738 24998 2790 25050
rect 2802 24998 2854 25050
rect 2866 24998 2918 25050
rect 10610 24998 10662 25050
rect 10674 24998 10726 25050
rect 10738 24998 10790 25050
rect 10802 24998 10854 25050
rect 10866 24998 10918 25050
rect 18610 24998 18662 25050
rect 18674 24998 18726 25050
rect 18738 24998 18790 25050
rect 18802 24998 18854 25050
rect 18866 24998 18918 25050
rect 26610 24998 26662 25050
rect 26674 24998 26726 25050
rect 26738 24998 26790 25050
rect 26802 24998 26854 25050
rect 26866 24998 26918 25050
rect 1950 24454 2002 24506
rect 2014 24454 2066 24506
rect 2078 24454 2130 24506
rect 2142 24454 2194 24506
rect 2206 24454 2258 24506
rect 9950 24454 10002 24506
rect 10014 24454 10066 24506
rect 10078 24454 10130 24506
rect 10142 24454 10194 24506
rect 10206 24454 10258 24506
rect 17950 24454 18002 24506
rect 18014 24454 18066 24506
rect 18078 24454 18130 24506
rect 18142 24454 18194 24506
rect 18206 24454 18258 24506
rect 25950 24454 26002 24506
rect 26014 24454 26066 24506
rect 26078 24454 26130 24506
rect 26142 24454 26194 24506
rect 26206 24454 26258 24506
rect 28080 24352 28132 24404
rect 27528 24191 27580 24200
rect 27528 24157 27537 24191
rect 27537 24157 27571 24191
rect 27571 24157 27580 24191
rect 27528 24148 27580 24157
rect 28080 24191 28132 24200
rect 28080 24157 28089 24191
rect 28089 24157 28123 24191
rect 28123 24157 28132 24191
rect 28080 24148 28132 24157
rect 28356 24123 28408 24132
rect 28356 24089 28365 24123
rect 28365 24089 28399 24123
rect 28399 24089 28408 24123
rect 28356 24080 28408 24089
rect 2610 23910 2662 23962
rect 2674 23910 2726 23962
rect 2738 23910 2790 23962
rect 2802 23910 2854 23962
rect 2866 23910 2918 23962
rect 10610 23910 10662 23962
rect 10674 23910 10726 23962
rect 10738 23910 10790 23962
rect 10802 23910 10854 23962
rect 10866 23910 10918 23962
rect 18610 23910 18662 23962
rect 18674 23910 18726 23962
rect 18738 23910 18790 23962
rect 18802 23910 18854 23962
rect 18866 23910 18918 23962
rect 26610 23910 26662 23962
rect 26674 23910 26726 23962
rect 26738 23910 26790 23962
rect 26802 23910 26854 23962
rect 26866 23910 26918 23962
rect 1950 23366 2002 23418
rect 2014 23366 2066 23418
rect 2078 23366 2130 23418
rect 2142 23366 2194 23418
rect 2206 23366 2258 23418
rect 9950 23366 10002 23418
rect 10014 23366 10066 23418
rect 10078 23366 10130 23418
rect 10142 23366 10194 23418
rect 10206 23366 10258 23418
rect 17950 23366 18002 23418
rect 18014 23366 18066 23418
rect 18078 23366 18130 23418
rect 18142 23366 18194 23418
rect 18206 23366 18258 23418
rect 25950 23366 26002 23418
rect 26014 23366 26066 23418
rect 26078 23366 26130 23418
rect 26142 23366 26194 23418
rect 26206 23366 26258 23418
rect 2610 22822 2662 22874
rect 2674 22822 2726 22874
rect 2738 22822 2790 22874
rect 2802 22822 2854 22874
rect 2866 22822 2918 22874
rect 10610 22822 10662 22874
rect 10674 22822 10726 22874
rect 10738 22822 10790 22874
rect 10802 22822 10854 22874
rect 10866 22822 10918 22874
rect 18610 22822 18662 22874
rect 18674 22822 18726 22874
rect 18738 22822 18790 22874
rect 18802 22822 18854 22874
rect 18866 22822 18918 22874
rect 26610 22822 26662 22874
rect 26674 22822 26726 22874
rect 26738 22822 26790 22874
rect 26802 22822 26854 22874
rect 26866 22822 26918 22874
rect 28080 22720 28132 22772
rect 848 22584 900 22636
rect 27436 22584 27488 22636
rect 28080 22627 28132 22636
rect 28080 22593 28089 22627
rect 28089 22593 28123 22627
rect 28123 22593 28132 22627
rect 28080 22584 28132 22593
rect 28356 22559 28408 22568
rect 28356 22525 28365 22559
rect 28365 22525 28399 22559
rect 28399 22525 28408 22559
rect 28356 22516 28408 22525
rect 1768 22423 1820 22432
rect 1768 22389 1777 22423
rect 1777 22389 1811 22423
rect 1811 22389 1820 22423
rect 1768 22380 1820 22389
rect 1950 22278 2002 22330
rect 2014 22278 2066 22330
rect 2078 22278 2130 22330
rect 2142 22278 2194 22330
rect 2206 22278 2258 22330
rect 9950 22278 10002 22330
rect 10014 22278 10066 22330
rect 10078 22278 10130 22330
rect 10142 22278 10194 22330
rect 10206 22278 10258 22330
rect 17950 22278 18002 22330
rect 18014 22278 18066 22330
rect 18078 22278 18130 22330
rect 18142 22278 18194 22330
rect 18206 22278 18258 22330
rect 25950 22278 26002 22330
rect 26014 22278 26066 22330
rect 26078 22278 26130 22330
rect 26142 22278 26194 22330
rect 26206 22278 26258 22330
rect 28080 22176 28132 22228
rect 27528 22015 27580 22024
rect 27528 21981 27537 22015
rect 27537 21981 27571 22015
rect 27571 21981 27580 22015
rect 27528 21972 27580 21981
rect 2610 21734 2662 21786
rect 2674 21734 2726 21786
rect 2738 21734 2790 21786
rect 2802 21734 2854 21786
rect 2866 21734 2918 21786
rect 10610 21734 10662 21786
rect 10674 21734 10726 21786
rect 10738 21734 10790 21786
rect 10802 21734 10854 21786
rect 10866 21734 10918 21786
rect 18610 21734 18662 21786
rect 18674 21734 18726 21786
rect 18738 21734 18790 21786
rect 18802 21734 18854 21786
rect 18866 21734 18918 21786
rect 26610 21734 26662 21786
rect 26674 21734 26726 21786
rect 26738 21734 26790 21786
rect 26802 21734 26854 21786
rect 26866 21734 26918 21786
rect 1950 21190 2002 21242
rect 2014 21190 2066 21242
rect 2078 21190 2130 21242
rect 2142 21190 2194 21242
rect 2206 21190 2258 21242
rect 9950 21190 10002 21242
rect 10014 21190 10066 21242
rect 10078 21190 10130 21242
rect 10142 21190 10194 21242
rect 10206 21190 10258 21242
rect 17950 21190 18002 21242
rect 18014 21190 18066 21242
rect 18078 21190 18130 21242
rect 18142 21190 18194 21242
rect 18206 21190 18258 21242
rect 25950 21190 26002 21242
rect 26014 21190 26066 21242
rect 26078 21190 26130 21242
rect 26142 21190 26194 21242
rect 26206 21190 26258 21242
rect 27436 20884 27488 20936
rect 28356 20859 28408 20868
rect 28356 20825 28365 20859
rect 28365 20825 28399 20859
rect 28399 20825 28408 20859
rect 28356 20816 28408 20825
rect 2610 20646 2662 20698
rect 2674 20646 2726 20698
rect 2738 20646 2790 20698
rect 2802 20646 2854 20698
rect 2866 20646 2918 20698
rect 10610 20646 10662 20698
rect 10674 20646 10726 20698
rect 10738 20646 10790 20698
rect 10802 20646 10854 20698
rect 10866 20646 10918 20698
rect 18610 20646 18662 20698
rect 18674 20646 18726 20698
rect 18738 20646 18790 20698
rect 18802 20646 18854 20698
rect 18866 20646 18918 20698
rect 26610 20646 26662 20698
rect 26674 20646 26726 20698
rect 26738 20646 26790 20698
rect 26802 20646 26854 20698
rect 26866 20646 26918 20698
rect 1950 20102 2002 20154
rect 2014 20102 2066 20154
rect 2078 20102 2130 20154
rect 2142 20102 2194 20154
rect 2206 20102 2258 20154
rect 9950 20102 10002 20154
rect 10014 20102 10066 20154
rect 10078 20102 10130 20154
rect 10142 20102 10194 20154
rect 10206 20102 10258 20154
rect 17950 20102 18002 20154
rect 18014 20102 18066 20154
rect 18078 20102 18130 20154
rect 18142 20102 18194 20154
rect 18206 20102 18258 20154
rect 25950 20102 26002 20154
rect 26014 20102 26066 20154
rect 26078 20102 26130 20154
rect 26142 20102 26194 20154
rect 26206 20102 26258 20154
rect 2610 19558 2662 19610
rect 2674 19558 2726 19610
rect 2738 19558 2790 19610
rect 2802 19558 2854 19610
rect 2866 19558 2918 19610
rect 10610 19558 10662 19610
rect 10674 19558 10726 19610
rect 10738 19558 10790 19610
rect 10802 19558 10854 19610
rect 10866 19558 10918 19610
rect 18610 19558 18662 19610
rect 18674 19558 18726 19610
rect 18738 19558 18790 19610
rect 18802 19558 18854 19610
rect 18866 19558 18918 19610
rect 26610 19558 26662 19610
rect 26674 19558 26726 19610
rect 26738 19558 26790 19610
rect 26802 19558 26854 19610
rect 26866 19558 26918 19610
rect 28080 19363 28132 19372
rect 28080 19329 28089 19363
rect 28089 19329 28123 19363
rect 28123 19329 28132 19363
rect 28080 19320 28132 19329
rect 28356 19363 28408 19372
rect 28356 19329 28365 19363
rect 28365 19329 28399 19363
rect 28399 19329 28408 19363
rect 28356 19320 28408 19329
rect 1950 19014 2002 19066
rect 2014 19014 2066 19066
rect 2078 19014 2130 19066
rect 2142 19014 2194 19066
rect 2206 19014 2258 19066
rect 9950 19014 10002 19066
rect 10014 19014 10066 19066
rect 10078 19014 10130 19066
rect 10142 19014 10194 19066
rect 10206 19014 10258 19066
rect 17950 19014 18002 19066
rect 18014 19014 18066 19066
rect 18078 19014 18130 19066
rect 18142 19014 18194 19066
rect 18206 19014 18258 19066
rect 25950 19014 26002 19066
rect 26014 19014 26066 19066
rect 26078 19014 26130 19066
rect 26142 19014 26194 19066
rect 26206 19014 26258 19066
rect 28080 18912 28132 18964
rect 27528 18751 27580 18760
rect 27528 18717 27537 18751
rect 27537 18717 27571 18751
rect 27571 18717 27580 18751
rect 27528 18708 27580 18717
rect 2610 18470 2662 18522
rect 2674 18470 2726 18522
rect 2738 18470 2790 18522
rect 2802 18470 2854 18522
rect 2866 18470 2918 18522
rect 10610 18470 10662 18522
rect 10674 18470 10726 18522
rect 10738 18470 10790 18522
rect 10802 18470 10854 18522
rect 10866 18470 10918 18522
rect 18610 18470 18662 18522
rect 18674 18470 18726 18522
rect 18738 18470 18790 18522
rect 18802 18470 18854 18522
rect 18866 18470 18918 18522
rect 26610 18470 26662 18522
rect 26674 18470 26726 18522
rect 26738 18470 26790 18522
rect 26802 18470 26854 18522
rect 26866 18470 26918 18522
rect 27620 18368 27672 18420
rect 27344 18232 27396 18284
rect 1950 17926 2002 17978
rect 2014 17926 2066 17978
rect 2078 17926 2130 17978
rect 2142 17926 2194 17978
rect 2206 17926 2258 17978
rect 9950 17926 10002 17978
rect 10014 17926 10066 17978
rect 10078 17926 10130 17978
rect 10142 17926 10194 17978
rect 10206 17926 10258 17978
rect 17950 17926 18002 17978
rect 18014 17926 18066 17978
rect 18078 17926 18130 17978
rect 18142 17926 18194 17978
rect 18206 17926 18258 17978
rect 25950 17926 26002 17978
rect 26014 17926 26066 17978
rect 26078 17926 26130 17978
rect 26142 17926 26194 17978
rect 26206 17926 26258 17978
rect 27344 17620 27396 17672
rect 28356 17595 28408 17604
rect 28356 17561 28365 17595
rect 28365 17561 28399 17595
rect 28399 17561 28408 17595
rect 28356 17552 28408 17561
rect 2610 17382 2662 17434
rect 2674 17382 2726 17434
rect 2738 17382 2790 17434
rect 2802 17382 2854 17434
rect 2866 17382 2918 17434
rect 10610 17382 10662 17434
rect 10674 17382 10726 17434
rect 10738 17382 10790 17434
rect 10802 17382 10854 17434
rect 10866 17382 10918 17434
rect 18610 17382 18662 17434
rect 18674 17382 18726 17434
rect 18738 17382 18790 17434
rect 18802 17382 18854 17434
rect 18866 17382 18918 17434
rect 26610 17382 26662 17434
rect 26674 17382 26726 17434
rect 26738 17382 26790 17434
rect 26802 17382 26854 17434
rect 26866 17382 26918 17434
rect 27436 17323 27488 17332
rect 27436 17289 27445 17323
rect 27445 17289 27479 17323
rect 27479 17289 27488 17323
rect 27436 17280 27488 17289
rect 26976 17119 27028 17128
rect 26976 17085 26985 17119
rect 26985 17085 27019 17119
rect 27019 17085 27028 17119
rect 26976 17076 27028 17085
rect 1768 16940 1820 16992
rect 26884 17008 26936 17060
rect 1950 16838 2002 16890
rect 2014 16838 2066 16890
rect 2078 16838 2130 16890
rect 2142 16838 2194 16890
rect 2206 16838 2258 16890
rect 9950 16838 10002 16890
rect 10014 16838 10066 16890
rect 10078 16838 10130 16890
rect 10142 16838 10194 16890
rect 10206 16838 10258 16890
rect 17950 16838 18002 16890
rect 18014 16838 18066 16890
rect 18078 16838 18130 16890
rect 18142 16838 18194 16890
rect 18206 16838 18258 16890
rect 25950 16838 26002 16890
rect 26014 16838 26066 16890
rect 26078 16838 26130 16890
rect 26142 16838 26194 16890
rect 26206 16838 26258 16890
rect 27344 16779 27396 16788
rect 27344 16745 27353 16779
rect 27353 16745 27387 16779
rect 27387 16745 27396 16779
rect 27344 16736 27396 16745
rect 26976 16668 27028 16720
rect 26884 16643 26936 16652
rect 26884 16609 26893 16643
rect 26893 16609 26927 16643
rect 26927 16609 26936 16643
rect 26884 16600 26936 16609
rect 27068 16600 27120 16652
rect 2610 16294 2662 16346
rect 2674 16294 2726 16346
rect 2738 16294 2790 16346
rect 2802 16294 2854 16346
rect 2866 16294 2918 16346
rect 10610 16294 10662 16346
rect 10674 16294 10726 16346
rect 10738 16294 10790 16346
rect 10802 16294 10854 16346
rect 10866 16294 10918 16346
rect 18610 16294 18662 16346
rect 18674 16294 18726 16346
rect 18738 16294 18790 16346
rect 18802 16294 18854 16346
rect 18866 16294 18918 16346
rect 26610 16294 26662 16346
rect 26674 16294 26726 16346
rect 26738 16294 26790 16346
rect 26802 16294 26854 16346
rect 26866 16294 26918 16346
rect 27528 16192 27580 16244
rect 27068 16056 27120 16108
rect 27160 16031 27212 16040
rect 27160 15997 27169 16031
rect 27169 15997 27203 16031
rect 27203 15997 27212 16031
rect 27160 15988 27212 15997
rect 1950 15750 2002 15802
rect 2014 15750 2066 15802
rect 2078 15750 2130 15802
rect 2142 15750 2194 15802
rect 2206 15750 2258 15802
rect 9950 15750 10002 15802
rect 10014 15750 10066 15802
rect 10078 15750 10130 15802
rect 10142 15750 10194 15802
rect 10206 15750 10258 15802
rect 17950 15750 18002 15802
rect 18014 15750 18066 15802
rect 18078 15750 18130 15802
rect 18142 15750 18194 15802
rect 18206 15750 18258 15802
rect 25950 15750 26002 15802
rect 26014 15750 26066 15802
rect 26078 15750 26130 15802
rect 26142 15750 26194 15802
rect 26206 15750 26258 15802
rect 28356 15555 28408 15564
rect 28356 15521 28365 15555
rect 28365 15521 28399 15555
rect 28399 15521 28408 15555
rect 28356 15512 28408 15521
rect 27528 15444 27580 15496
rect 2610 15206 2662 15258
rect 2674 15206 2726 15258
rect 2738 15206 2790 15258
rect 2802 15206 2854 15258
rect 2866 15206 2918 15258
rect 10610 15206 10662 15258
rect 10674 15206 10726 15258
rect 10738 15206 10790 15258
rect 10802 15206 10854 15258
rect 10866 15206 10918 15258
rect 18610 15206 18662 15258
rect 18674 15206 18726 15258
rect 18738 15206 18790 15258
rect 18802 15206 18854 15258
rect 18866 15206 18918 15258
rect 26610 15206 26662 15258
rect 26674 15206 26726 15258
rect 26738 15206 26790 15258
rect 26802 15206 26854 15258
rect 26866 15206 26918 15258
rect 1950 14662 2002 14714
rect 2014 14662 2066 14714
rect 2078 14662 2130 14714
rect 2142 14662 2194 14714
rect 2206 14662 2258 14714
rect 9950 14662 10002 14714
rect 10014 14662 10066 14714
rect 10078 14662 10130 14714
rect 10142 14662 10194 14714
rect 10206 14662 10258 14714
rect 17950 14662 18002 14714
rect 18014 14662 18066 14714
rect 18078 14662 18130 14714
rect 18142 14662 18194 14714
rect 18206 14662 18258 14714
rect 25950 14662 26002 14714
rect 26014 14662 26066 14714
rect 26078 14662 26130 14714
rect 26142 14662 26194 14714
rect 26206 14662 26258 14714
rect 28080 14399 28132 14408
rect 28080 14365 28089 14399
rect 28089 14365 28123 14399
rect 28123 14365 28132 14399
rect 28080 14356 28132 14365
rect 28356 14331 28408 14340
rect 28356 14297 28365 14331
rect 28365 14297 28399 14331
rect 28399 14297 28408 14331
rect 28356 14288 28408 14297
rect 2610 14118 2662 14170
rect 2674 14118 2726 14170
rect 2738 14118 2790 14170
rect 2802 14118 2854 14170
rect 2866 14118 2918 14170
rect 10610 14118 10662 14170
rect 10674 14118 10726 14170
rect 10738 14118 10790 14170
rect 10802 14118 10854 14170
rect 10866 14118 10918 14170
rect 18610 14118 18662 14170
rect 18674 14118 18726 14170
rect 18738 14118 18790 14170
rect 18802 14118 18854 14170
rect 18866 14118 18918 14170
rect 26610 14118 26662 14170
rect 26674 14118 26726 14170
rect 26738 14118 26790 14170
rect 26802 14118 26854 14170
rect 26866 14118 26918 14170
rect 1950 13574 2002 13626
rect 2014 13574 2066 13626
rect 2078 13574 2130 13626
rect 2142 13574 2194 13626
rect 2206 13574 2258 13626
rect 9950 13574 10002 13626
rect 10014 13574 10066 13626
rect 10078 13574 10130 13626
rect 10142 13574 10194 13626
rect 10206 13574 10258 13626
rect 17950 13574 18002 13626
rect 18014 13574 18066 13626
rect 18078 13574 18130 13626
rect 18142 13574 18194 13626
rect 18206 13574 18258 13626
rect 25950 13574 26002 13626
rect 26014 13574 26066 13626
rect 26078 13574 26130 13626
rect 26142 13574 26194 13626
rect 26206 13574 26258 13626
rect 28080 13472 28132 13524
rect 27620 13268 27672 13320
rect 2610 13030 2662 13082
rect 2674 13030 2726 13082
rect 2738 13030 2790 13082
rect 2802 13030 2854 13082
rect 2866 13030 2918 13082
rect 10610 13030 10662 13082
rect 10674 13030 10726 13082
rect 10738 13030 10790 13082
rect 10802 13030 10854 13082
rect 10866 13030 10918 13082
rect 18610 13030 18662 13082
rect 18674 13030 18726 13082
rect 18738 13030 18790 13082
rect 18802 13030 18854 13082
rect 18866 13030 18918 13082
rect 26610 13030 26662 13082
rect 26674 13030 26726 13082
rect 26738 13030 26790 13082
rect 26802 13030 26854 13082
rect 26866 13030 26918 13082
rect 27068 12835 27120 12844
rect 27068 12801 27077 12835
rect 27077 12801 27111 12835
rect 27111 12801 27120 12835
rect 27068 12792 27120 12801
rect 27160 12835 27212 12844
rect 27160 12801 27169 12835
rect 27169 12801 27203 12835
rect 27203 12801 27212 12835
rect 27160 12792 27212 12801
rect 28080 12835 28132 12844
rect 28080 12801 28089 12835
rect 28089 12801 28123 12835
rect 28123 12801 28132 12835
rect 28080 12792 28132 12801
rect 28356 12767 28408 12776
rect 28356 12733 28365 12767
rect 28365 12733 28399 12767
rect 28399 12733 28408 12767
rect 28356 12724 28408 12733
rect 27620 12588 27672 12640
rect 28172 12588 28224 12640
rect 1950 12486 2002 12538
rect 2014 12486 2066 12538
rect 2078 12486 2130 12538
rect 2142 12486 2194 12538
rect 2206 12486 2258 12538
rect 9950 12486 10002 12538
rect 10014 12486 10066 12538
rect 10078 12486 10130 12538
rect 10142 12486 10194 12538
rect 10206 12486 10258 12538
rect 17950 12486 18002 12538
rect 18014 12486 18066 12538
rect 18078 12486 18130 12538
rect 18142 12486 18194 12538
rect 18206 12486 18258 12538
rect 25950 12486 26002 12538
rect 26014 12486 26066 12538
rect 26078 12486 26130 12538
rect 26142 12486 26194 12538
rect 26206 12486 26258 12538
rect 2610 11942 2662 11994
rect 2674 11942 2726 11994
rect 2738 11942 2790 11994
rect 2802 11942 2854 11994
rect 2866 11942 2918 11994
rect 10610 11942 10662 11994
rect 10674 11942 10726 11994
rect 10738 11942 10790 11994
rect 10802 11942 10854 11994
rect 10866 11942 10918 11994
rect 18610 11942 18662 11994
rect 18674 11942 18726 11994
rect 18738 11942 18790 11994
rect 18802 11942 18854 11994
rect 18866 11942 18918 11994
rect 26610 11942 26662 11994
rect 26674 11942 26726 11994
rect 26738 11942 26790 11994
rect 26802 11942 26854 11994
rect 26866 11942 26918 11994
rect 28080 11840 28132 11892
rect 27436 11704 27488 11756
rect 1950 11398 2002 11450
rect 2014 11398 2066 11450
rect 2078 11398 2130 11450
rect 2142 11398 2194 11450
rect 2206 11398 2258 11450
rect 9950 11398 10002 11450
rect 10014 11398 10066 11450
rect 10078 11398 10130 11450
rect 10142 11398 10194 11450
rect 10206 11398 10258 11450
rect 17950 11398 18002 11450
rect 18014 11398 18066 11450
rect 18078 11398 18130 11450
rect 18142 11398 18194 11450
rect 18206 11398 18258 11450
rect 25950 11398 26002 11450
rect 26014 11398 26066 11450
rect 26078 11398 26130 11450
rect 26142 11398 26194 11450
rect 26206 11398 26258 11450
rect 28080 11135 28132 11144
rect 28080 11101 28089 11135
rect 28089 11101 28123 11135
rect 28123 11101 28132 11135
rect 28080 11092 28132 11101
rect 28356 11067 28408 11076
rect 28356 11033 28365 11067
rect 28365 11033 28399 11067
rect 28399 11033 28408 11067
rect 28356 11024 28408 11033
rect 2610 10854 2662 10906
rect 2674 10854 2726 10906
rect 2738 10854 2790 10906
rect 2802 10854 2854 10906
rect 2866 10854 2918 10906
rect 10610 10854 10662 10906
rect 10674 10854 10726 10906
rect 10738 10854 10790 10906
rect 10802 10854 10854 10906
rect 10866 10854 10918 10906
rect 18610 10854 18662 10906
rect 18674 10854 18726 10906
rect 18738 10854 18790 10906
rect 18802 10854 18854 10906
rect 18866 10854 18918 10906
rect 26610 10854 26662 10906
rect 26674 10854 26726 10906
rect 26738 10854 26790 10906
rect 26802 10854 26854 10906
rect 26866 10854 26918 10906
rect 26516 10616 26568 10668
rect 27252 10752 27304 10804
rect 27436 10684 27488 10736
rect 27068 10659 27120 10668
rect 27068 10625 27077 10659
rect 27077 10625 27111 10659
rect 27111 10625 27120 10659
rect 27068 10616 27120 10625
rect 27252 10616 27304 10668
rect 27528 10480 27580 10532
rect 1950 10310 2002 10362
rect 2014 10310 2066 10362
rect 2078 10310 2130 10362
rect 2142 10310 2194 10362
rect 2206 10310 2258 10362
rect 9950 10310 10002 10362
rect 10014 10310 10066 10362
rect 10078 10310 10130 10362
rect 10142 10310 10194 10362
rect 10206 10310 10258 10362
rect 17950 10310 18002 10362
rect 18014 10310 18066 10362
rect 18078 10310 18130 10362
rect 18142 10310 18194 10362
rect 18206 10310 18258 10362
rect 25950 10310 26002 10362
rect 26014 10310 26066 10362
rect 26078 10310 26130 10362
rect 26142 10310 26194 10362
rect 26206 10310 26258 10362
rect 2610 9766 2662 9818
rect 2674 9766 2726 9818
rect 2738 9766 2790 9818
rect 2802 9766 2854 9818
rect 2866 9766 2918 9818
rect 10610 9766 10662 9818
rect 10674 9766 10726 9818
rect 10738 9766 10790 9818
rect 10802 9766 10854 9818
rect 10866 9766 10918 9818
rect 18610 9766 18662 9818
rect 18674 9766 18726 9818
rect 18738 9766 18790 9818
rect 18802 9766 18854 9818
rect 18866 9766 18918 9818
rect 26610 9766 26662 9818
rect 26674 9766 26726 9818
rect 26738 9766 26790 9818
rect 26802 9766 26854 9818
rect 26866 9766 26918 9818
rect 27528 9571 27580 9580
rect 27528 9537 27537 9571
rect 27537 9537 27571 9571
rect 27571 9537 27580 9571
rect 27528 9528 27580 9537
rect 27712 9528 27764 9580
rect 28356 9503 28408 9512
rect 28356 9469 28365 9503
rect 28365 9469 28399 9503
rect 28399 9469 28408 9503
rect 28356 9460 28408 9469
rect 28080 9392 28132 9444
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 9950 9222 10002 9274
rect 10014 9222 10066 9274
rect 10078 9222 10130 9274
rect 10142 9222 10194 9274
rect 10206 9222 10258 9274
rect 17950 9222 18002 9274
rect 18014 9222 18066 9274
rect 18078 9222 18130 9274
rect 18142 9222 18194 9274
rect 18206 9222 18258 9274
rect 25950 9222 26002 9274
rect 26014 9222 26066 9274
rect 26078 9222 26130 9274
rect 26142 9222 26194 9274
rect 26206 9222 26258 9274
rect 27712 9163 27764 9172
rect 27712 9129 27721 9163
rect 27721 9129 27755 9163
rect 27755 9129 27764 9163
rect 27712 9120 27764 9129
rect 27436 8916 27488 8968
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 10610 8678 10662 8730
rect 10674 8678 10726 8730
rect 10738 8678 10790 8730
rect 10802 8678 10854 8730
rect 10866 8678 10918 8730
rect 18610 8678 18662 8730
rect 18674 8678 18726 8730
rect 18738 8678 18790 8730
rect 18802 8678 18854 8730
rect 18866 8678 18918 8730
rect 26610 8678 26662 8730
rect 26674 8678 26726 8730
rect 26738 8678 26790 8730
rect 26802 8678 26854 8730
rect 26866 8678 26918 8730
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 9950 8134 10002 8186
rect 10014 8134 10066 8186
rect 10078 8134 10130 8186
rect 10142 8134 10194 8186
rect 10206 8134 10258 8186
rect 17950 8134 18002 8186
rect 18014 8134 18066 8186
rect 18078 8134 18130 8186
rect 18142 8134 18194 8186
rect 18206 8134 18258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 27528 7828 27580 7880
rect 848 7760 900 7812
rect 28356 7803 28408 7812
rect 28356 7769 28365 7803
rect 28365 7769 28399 7803
rect 28399 7769 28408 7803
rect 28356 7760 28408 7769
rect 26516 7692 26568 7744
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 10610 7590 10662 7642
rect 10674 7590 10726 7642
rect 10738 7590 10790 7642
rect 10802 7590 10854 7642
rect 10866 7590 10918 7642
rect 18610 7590 18662 7642
rect 18674 7590 18726 7642
rect 18738 7590 18790 7642
rect 18802 7590 18854 7642
rect 18866 7590 18918 7642
rect 26610 7590 26662 7642
rect 26674 7590 26726 7642
rect 26738 7590 26790 7642
rect 26802 7590 26854 7642
rect 26866 7590 26918 7642
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 9950 7046 10002 7098
rect 10014 7046 10066 7098
rect 10078 7046 10130 7098
rect 10142 7046 10194 7098
rect 10206 7046 10258 7098
rect 17950 7046 18002 7098
rect 18014 7046 18066 7098
rect 18078 7046 18130 7098
rect 18142 7046 18194 7098
rect 18206 7046 18258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 10610 6502 10662 6554
rect 10674 6502 10726 6554
rect 10738 6502 10790 6554
rect 10802 6502 10854 6554
rect 10866 6502 10918 6554
rect 18610 6502 18662 6554
rect 18674 6502 18726 6554
rect 18738 6502 18790 6554
rect 18802 6502 18854 6554
rect 18866 6502 18918 6554
rect 26610 6502 26662 6554
rect 26674 6502 26726 6554
rect 26738 6502 26790 6554
rect 26802 6502 26854 6554
rect 26866 6502 26918 6554
rect 27712 6264 27764 6316
rect 28356 6239 28408 6248
rect 28356 6205 28365 6239
rect 28365 6205 28399 6239
rect 28399 6205 28408 6239
rect 28356 6196 28408 6205
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 9950 5958 10002 6010
rect 10014 5958 10066 6010
rect 10078 5958 10130 6010
rect 10142 5958 10194 6010
rect 10206 5958 10258 6010
rect 17950 5958 18002 6010
rect 18014 5958 18066 6010
rect 18078 5958 18130 6010
rect 18142 5958 18194 6010
rect 18206 5958 18258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 27712 5899 27764 5908
rect 27712 5865 27721 5899
rect 27721 5865 27755 5899
rect 27755 5865 27764 5899
rect 27712 5856 27764 5865
rect 27528 5695 27580 5704
rect 27528 5661 27537 5695
rect 27537 5661 27571 5695
rect 27571 5661 27580 5695
rect 27528 5652 27580 5661
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 10610 5414 10662 5466
rect 10674 5414 10726 5466
rect 10738 5414 10790 5466
rect 10802 5414 10854 5466
rect 10866 5414 10918 5466
rect 18610 5414 18662 5466
rect 18674 5414 18726 5466
rect 18738 5414 18790 5466
rect 18802 5414 18854 5466
rect 18866 5414 18918 5466
rect 26610 5414 26662 5466
rect 26674 5414 26726 5466
rect 26738 5414 26790 5466
rect 26802 5414 26854 5466
rect 26866 5414 26918 5466
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 9950 4870 10002 4922
rect 10014 4870 10066 4922
rect 10078 4870 10130 4922
rect 10142 4870 10194 4922
rect 10206 4870 10258 4922
rect 17950 4870 18002 4922
rect 18014 4870 18066 4922
rect 18078 4870 18130 4922
rect 18142 4870 18194 4922
rect 18206 4870 18258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 28172 4564 28224 4616
rect 28356 4539 28408 4548
rect 28356 4505 28365 4539
rect 28365 4505 28399 4539
rect 28399 4505 28408 4539
rect 28356 4496 28408 4505
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 10610 4326 10662 4378
rect 10674 4326 10726 4378
rect 10738 4326 10790 4378
rect 10802 4326 10854 4378
rect 10866 4326 10918 4378
rect 18610 4326 18662 4378
rect 18674 4326 18726 4378
rect 18738 4326 18790 4378
rect 18802 4326 18854 4378
rect 18866 4326 18918 4378
rect 26610 4326 26662 4378
rect 26674 4326 26726 4378
rect 26738 4326 26790 4378
rect 26802 4326 26854 4378
rect 26866 4326 26918 4378
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 9950 3782 10002 3834
rect 10014 3782 10066 3834
rect 10078 3782 10130 3834
rect 10142 3782 10194 3834
rect 10206 3782 10258 3834
rect 17950 3782 18002 3834
rect 18014 3782 18066 3834
rect 18078 3782 18130 3834
rect 18142 3782 18194 3834
rect 18206 3782 18258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 10610 3238 10662 3290
rect 10674 3238 10726 3290
rect 10738 3238 10790 3290
rect 10802 3238 10854 3290
rect 10866 3238 10918 3290
rect 18610 3238 18662 3290
rect 18674 3238 18726 3290
rect 18738 3238 18790 3290
rect 18802 3238 18854 3290
rect 18866 3238 18918 3290
rect 26610 3238 26662 3290
rect 26674 3238 26726 3290
rect 26738 3238 26790 3290
rect 26802 3238 26854 3290
rect 26866 3238 26918 3290
rect 27528 3000 27580 3052
rect 28356 2975 28408 2984
rect 28356 2941 28365 2975
rect 28365 2941 28399 2975
rect 28399 2941 28408 2975
rect 28356 2932 28408 2941
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 9950 2694 10002 2746
rect 10014 2694 10066 2746
rect 10078 2694 10130 2746
rect 10142 2694 10194 2746
rect 10206 2694 10258 2746
rect 17950 2694 18002 2746
rect 18014 2694 18066 2746
rect 18078 2694 18130 2746
rect 18142 2694 18194 2746
rect 18206 2694 18258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
rect 10610 2150 10662 2202
rect 10674 2150 10726 2202
rect 10738 2150 10790 2202
rect 10802 2150 10854 2202
rect 10866 2150 10918 2202
rect 18610 2150 18662 2202
rect 18674 2150 18726 2202
rect 18738 2150 18790 2202
rect 18802 2150 18854 2202
rect 18866 2150 18918 2202
rect 26610 2150 26662 2202
rect 26674 2150 26726 2202
rect 26738 2150 26790 2202
rect 26802 2150 26854 2202
rect 26866 2150 26918 2202
<< metal2 >>
rect 1950 27772 2258 27781
rect 1950 27770 1956 27772
rect 2012 27770 2036 27772
rect 2092 27770 2116 27772
rect 2172 27770 2196 27772
rect 2252 27770 2258 27772
rect 2012 27718 2014 27770
rect 2194 27718 2196 27770
rect 1950 27716 1956 27718
rect 2012 27716 2036 27718
rect 2092 27716 2116 27718
rect 2172 27716 2196 27718
rect 2252 27716 2258 27718
rect 1950 27707 2258 27716
rect 9950 27772 10258 27781
rect 9950 27770 9956 27772
rect 10012 27770 10036 27772
rect 10092 27770 10116 27772
rect 10172 27770 10196 27772
rect 10252 27770 10258 27772
rect 10012 27718 10014 27770
rect 10194 27718 10196 27770
rect 9950 27716 9956 27718
rect 10012 27716 10036 27718
rect 10092 27716 10116 27718
rect 10172 27716 10196 27718
rect 10252 27716 10258 27718
rect 9950 27707 10258 27716
rect 17950 27772 18258 27781
rect 17950 27770 17956 27772
rect 18012 27770 18036 27772
rect 18092 27770 18116 27772
rect 18172 27770 18196 27772
rect 18252 27770 18258 27772
rect 18012 27718 18014 27770
rect 18194 27718 18196 27770
rect 17950 27716 17956 27718
rect 18012 27716 18036 27718
rect 18092 27716 18116 27718
rect 18172 27716 18196 27718
rect 18252 27716 18258 27718
rect 17950 27707 18258 27716
rect 25950 27772 26258 27781
rect 25950 27770 25956 27772
rect 26012 27770 26036 27772
rect 26092 27770 26116 27772
rect 26172 27770 26196 27772
rect 26252 27770 26258 27772
rect 26012 27718 26014 27770
rect 26194 27718 26196 27770
rect 25950 27716 25956 27718
rect 26012 27716 26036 27718
rect 26092 27716 26116 27718
rect 26172 27716 26196 27718
rect 26252 27716 26258 27718
rect 25950 27707 26258 27716
rect 27620 27464 27672 27470
rect 27620 27406 27672 27412
rect 2610 27228 2918 27237
rect 2610 27226 2616 27228
rect 2672 27226 2696 27228
rect 2752 27226 2776 27228
rect 2832 27226 2856 27228
rect 2912 27226 2918 27228
rect 2672 27174 2674 27226
rect 2854 27174 2856 27226
rect 2610 27172 2616 27174
rect 2672 27172 2696 27174
rect 2752 27172 2776 27174
rect 2832 27172 2856 27174
rect 2912 27172 2918 27174
rect 2610 27163 2918 27172
rect 10610 27228 10918 27237
rect 10610 27226 10616 27228
rect 10672 27226 10696 27228
rect 10752 27226 10776 27228
rect 10832 27226 10856 27228
rect 10912 27226 10918 27228
rect 10672 27174 10674 27226
rect 10854 27174 10856 27226
rect 10610 27172 10616 27174
rect 10672 27172 10696 27174
rect 10752 27172 10776 27174
rect 10832 27172 10856 27174
rect 10912 27172 10918 27174
rect 10610 27163 10918 27172
rect 18610 27228 18918 27237
rect 18610 27226 18616 27228
rect 18672 27226 18696 27228
rect 18752 27226 18776 27228
rect 18832 27226 18856 27228
rect 18912 27226 18918 27228
rect 18672 27174 18674 27226
rect 18854 27174 18856 27226
rect 18610 27172 18616 27174
rect 18672 27172 18696 27174
rect 18752 27172 18776 27174
rect 18832 27172 18856 27174
rect 18912 27172 18918 27174
rect 18610 27163 18918 27172
rect 26610 27228 26918 27237
rect 26610 27226 26616 27228
rect 26672 27226 26696 27228
rect 26752 27226 26776 27228
rect 26832 27226 26856 27228
rect 26912 27226 26918 27228
rect 26672 27174 26674 27226
rect 26854 27174 26856 27226
rect 26610 27172 26616 27174
rect 26672 27172 26696 27174
rect 26752 27172 26776 27174
rect 26832 27172 26856 27174
rect 26912 27172 26918 27174
rect 26610 27163 26918 27172
rect 1950 26684 2258 26693
rect 1950 26682 1956 26684
rect 2012 26682 2036 26684
rect 2092 26682 2116 26684
rect 2172 26682 2196 26684
rect 2252 26682 2258 26684
rect 2012 26630 2014 26682
rect 2194 26630 2196 26682
rect 1950 26628 1956 26630
rect 2012 26628 2036 26630
rect 2092 26628 2116 26630
rect 2172 26628 2196 26630
rect 2252 26628 2258 26630
rect 1950 26619 2258 26628
rect 9950 26684 10258 26693
rect 9950 26682 9956 26684
rect 10012 26682 10036 26684
rect 10092 26682 10116 26684
rect 10172 26682 10196 26684
rect 10252 26682 10258 26684
rect 10012 26630 10014 26682
rect 10194 26630 10196 26682
rect 9950 26628 9956 26630
rect 10012 26628 10036 26630
rect 10092 26628 10116 26630
rect 10172 26628 10196 26630
rect 10252 26628 10258 26630
rect 9950 26619 10258 26628
rect 17950 26684 18258 26693
rect 17950 26682 17956 26684
rect 18012 26682 18036 26684
rect 18092 26682 18116 26684
rect 18172 26682 18196 26684
rect 18252 26682 18258 26684
rect 18012 26630 18014 26682
rect 18194 26630 18196 26682
rect 17950 26628 17956 26630
rect 18012 26628 18036 26630
rect 18092 26628 18116 26630
rect 18172 26628 18196 26630
rect 18252 26628 18258 26630
rect 17950 26619 18258 26628
rect 25950 26684 26258 26693
rect 25950 26682 25956 26684
rect 26012 26682 26036 26684
rect 26092 26682 26116 26684
rect 26172 26682 26196 26684
rect 26252 26682 26258 26684
rect 26012 26630 26014 26682
rect 26194 26630 26196 26682
rect 25950 26628 25956 26630
rect 26012 26628 26036 26630
rect 26092 26628 26116 26630
rect 26172 26628 26196 26630
rect 26252 26628 26258 26630
rect 25950 26619 26258 26628
rect 2610 26140 2918 26149
rect 2610 26138 2616 26140
rect 2672 26138 2696 26140
rect 2752 26138 2776 26140
rect 2832 26138 2856 26140
rect 2912 26138 2918 26140
rect 2672 26086 2674 26138
rect 2854 26086 2856 26138
rect 2610 26084 2616 26086
rect 2672 26084 2696 26086
rect 2752 26084 2776 26086
rect 2832 26084 2856 26086
rect 2912 26084 2918 26086
rect 2610 26075 2918 26084
rect 10610 26140 10918 26149
rect 10610 26138 10616 26140
rect 10672 26138 10696 26140
rect 10752 26138 10776 26140
rect 10832 26138 10856 26140
rect 10912 26138 10918 26140
rect 10672 26086 10674 26138
rect 10854 26086 10856 26138
rect 10610 26084 10616 26086
rect 10672 26084 10696 26086
rect 10752 26084 10776 26086
rect 10832 26084 10856 26086
rect 10912 26084 10918 26086
rect 10610 26075 10918 26084
rect 18610 26140 18918 26149
rect 18610 26138 18616 26140
rect 18672 26138 18696 26140
rect 18752 26138 18776 26140
rect 18832 26138 18856 26140
rect 18912 26138 18918 26140
rect 18672 26086 18674 26138
rect 18854 26086 18856 26138
rect 18610 26084 18616 26086
rect 18672 26084 18696 26086
rect 18752 26084 18776 26086
rect 18832 26084 18856 26086
rect 18912 26084 18918 26086
rect 18610 26075 18918 26084
rect 26610 26140 26918 26149
rect 26610 26138 26616 26140
rect 26672 26138 26696 26140
rect 26752 26138 26776 26140
rect 26832 26138 26856 26140
rect 26912 26138 26918 26140
rect 26672 26086 26674 26138
rect 26854 26086 26856 26138
rect 26610 26084 26616 26086
rect 26672 26084 26696 26086
rect 26752 26084 26776 26086
rect 26832 26084 26856 26086
rect 26912 26084 26918 26086
rect 26610 26075 26918 26084
rect 1950 25596 2258 25605
rect 1950 25594 1956 25596
rect 2012 25594 2036 25596
rect 2092 25594 2116 25596
rect 2172 25594 2196 25596
rect 2252 25594 2258 25596
rect 2012 25542 2014 25594
rect 2194 25542 2196 25594
rect 1950 25540 1956 25542
rect 2012 25540 2036 25542
rect 2092 25540 2116 25542
rect 2172 25540 2196 25542
rect 2252 25540 2258 25542
rect 1950 25531 2258 25540
rect 9950 25596 10258 25605
rect 9950 25594 9956 25596
rect 10012 25594 10036 25596
rect 10092 25594 10116 25596
rect 10172 25594 10196 25596
rect 10252 25594 10258 25596
rect 10012 25542 10014 25594
rect 10194 25542 10196 25594
rect 9950 25540 9956 25542
rect 10012 25540 10036 25542
rect 10092 25540 10116 25542
rect 10172 25540 10196 25542
rect 10252 25540 10258 25542
rect 9950 25531 10258 25540
rect 17950 25596 18258 25605
rect 17950 25594 17956 25596
rect 18012 25594 18036 25596
rect 18092 25594 18116 25596
rect 18172 25594 18196 25596
rect 18252 25594 18258 25596
rect 18012 25542 18014 25594
rect 18194 25542 18196 25594
rect 17950 25540 17956 25542
rect 18012 25540 18036 25542
rect 18092 25540 18116 25542
rect 18172 25540 18196 25542
rect 18252 25540 18258 25542
rect 17950 25531 18258 25540
rect 25950 25596 26258 25605
rect 25950 25594 25956 25596
rect 26012 25594 26036 25596
rect 26092 25594 26116 25596
rect 26172 25594 26196 25596
rect 26252 25594 26258 25596
rect 26012 25542 26014 25594
rect 26194 25542 26196 25594
rect 25950 25540 25956 25542
rect 26012 25540 26036 25542
rect 26092 25540 26116 25542
rect 26172 25540 26196 25542
rect 26252 25540 26258 25542
rect 25950 25531 26258 25540
rect 2610 25052 2918 25061
rect 2610 25050 2616 25052
rect 2672 25050 2696 25052
rect 2752 25050 2776 25052
rect 2832 25050 2856 25052
rect 2912 25050 2918 25052
rect 2672 24998 2674 25050
rect 2854 24998 2856 25050
rect 2610 24996 2616 24998
rect 2672 24996 2696 24998
rect 2752 24996 2776 24998
rect 2832 24996 2856 24998
rect 2912 24996 2918 24998
rect 2610 24987 2918 24996
rect 10610 25052 10918 25061
rect 10610 25050 10616 25052
rect 10672 25050 10696 25052
rect 10752 25050 10776 25052
rect 10832 25050 10856 25052
rect 10912 25050 10918 25052
rect 10672 24998 10674 25050
rect 10854 24998 10856 25050
rect 10610 24996 10616 24998
rect 10672 24996 10696 24998
rect 10752 24996 10776 24998
rect 10832 24996 10856 24998
rect 10912 24996 10918 24998
rect 10610 24987 10918 24996
rect 18610 25052 18918 25061
rect 18610 25050 18616 25052
rect 18672 25050 18696 25052
rect 18752 25050 18776 25052
rect 18832 25050 18856 25052
rect 18912 25050 18918 25052
rect 18672 24998 18674 25050
rect 18854 24998 18856 25050
rect 18610 24996 18616 24998
rect 18672 24996 18696 24998
rect 18752 24996 18776 24998
rect 18832 24996 18856 24998
rect 18912 24996 18918 24998
rect 18610 24987 18918 24996
rect 26610 25052 26918 25061
rect 26610 25050 26616 25052
rect 26672 25050 26696 25052
rect 26752 25050 26776 25052
rect 26832 25050 26856 25052
rect 26912 25050 26918 25052
rect 26672 24998 26674 25050
rect 26854 24998 26856 25050
rect 26610 24996 26616 24998
rect 26672 24996 26696 24998
rect 26752 24996 26776 24998
rect 26832 24996 26856 24998
rect 26912 24996 26918 24998
rect 26610 24987 26918 24996
rect 1950 24508 2258 24517
rect 1950 24506 1956 24508
rect 2012 24506 2036 24508
rect 2092 24506 2116 24508
rect 2172 24506 2196 24508
rect 2252 24506 2258 24508
rect 2012 24454 2014 24506
rect 2194 24454 2196 24506
rect 1950 24452 1956 24454
rect 2012 24452 2036 24454
rect 2092 24452 2116 24454
rect 2172 24452 2196 24454
rect 2252 24452 2258 24454
rect 1950 24443 2258 24452
rect 9950 24508 10258 24517
rect 9950 24506 9956 24508
rect 10012 24506 10036 24508
rect 10092 24506 10116 24508
rect 10172 24506 10196 24508
rect 10252 24506 10258 24508
rect 10012 24454 10014 24506
rect 10194 24454 10196 24506
rect 9950 24452 9956 24454
rect 10012 24452 10036 24454
rect 10092 24452 10116 24454
rect 10172 24452 10196 24454
rect 10252 24452 10258 24454
rect 9950 24443 10258 24452
rect 17950 24508 18258 24517
rect 17950 24506 17956 24508
rect 18012 24506 18036 24508
rect 18092 24506 18116 24508
rect 18172 24506 18196 24508
rect 18252 24506 18258 24508
rect 18012 24454 18014 24506
rect 18194 24454 18196 24506
rect 17950 24452 17956 24454
rect 18012 24452 18036 24454
rect 18092 24452 18116 24454
rect 18172 24452 18196 24454
rect 18252 24452 18258 24454
rect 17950 24443 18258 24452
rect 25950 24508 26258 24517
rect 25950 24506 25956 24508
rect 26012 24506 26036 24508
rect 26092 24506 26116 24508
rect 26172 24506 26196 24508
rect 26252 24506 26258 24508
rect 26012 24454 26014 24506
rect 26194 24454 26196 24506
rect 25950 24452 25956 24454
rect 26012 24452 26036 24454
rect 26092 24452 26116 24454
rect 26172 24452 26196 24454
rect 26252 24452 26258 24454
rect 25950 24443 26258 24452
rect 27528 24200 27580 24206
rect 27528 24142 27580 24148
rect 2610 23964 2918 23973
rect 2610 23962 2616 23964
rect 2672 23962 2696 23964
rect 2752 23962 2776 23964
rect 2832 23962 2856 23964
rect 2912 23962 2918 23964
rect 2672 23910 2674 23962
rect 2854 23910 2856 23962
rect 2610 23908 2616 23910
rect 2672 23908 2696 23910
rect 2752 23908 2776 23910
rect 2832 23908 2856 23910
rect 2912 23908 2918 23910
rect 2610 23899 2918 23908
rect 10610 23964 10918 23973
rect 10610 23962 10616 23964
rect 10672 23962 10696 23964
rect 10752 23962 10776 23964
rect 10832 23962 10856 23964
rect 10912 23962 10918 23964
rect 10672 23910 10674 23962
rect 10854 23910 10856 23962
rect 10610 23908 10616 23910
rect 10672 23908 10696 23910
rect 10752 23908 10776 23910
rect 10832 23908 10856 23910
rect 10912 23908 10918 23910
rect 10610 23899 10918 23908
rect 18610 23964 18918 23973
rect 18610 23962 18616 23964
rect 18672 23962 18696 23964
rect 18752 23962 18776 23964
rect 18832 23962 18856 23964
rect 18912 23962 18918 23964
rect 18672 23910 18674 23962
rect 18854 23910 18856 23962
rect 18610 23908 18616 23910
rect 18672 23908 18696 23910
rect 18752 23908 18776 23910
rect 18832 23908 18856 23910
rect 18912 23908 18918 23910
rect 18610 23899 18918 23908
rect 26610 23964 26918 23973
rect 26610 23962 26616 23964
rect 26672 23962 26696 23964
rect 26752 23962 26776 23964
rect 26832 23962 26856 23964
rect 26912 23962 26918 23964
rect 26672 23910 26674 23962
rect 26854 23910 26856 23962
rect 26610 23908 26616 23910
rect 26672 23908 26696 23910
rect 26752 23908 26776 23910
rect 26832 23908 26856 23910
rect 26912 23908 26918 23910
rect 26610 23899 26918 23908
rect 1950 23420 2258 23429
rect 1950 23418 1956 23420
rect 2012 23418 2036 23420
rect 2092 23418 2116 23420
rect 2172 23418 2196 23420
rect 2252 23418 2258 23420
rect 2012 23366 2014 23418
rect 2194 23366 2196 23418
rect 1950 23364 1956 23366
rect 2012 23364 2036 23366
rect 2092 23364 2116 23366
rect 2172 23364 2196 23366
rect 2252 23364 2258 23366
rect 1950 23355 2258 23364
rect 9950 23420 10258 23429
rect 9950 23418 9956 23420
rect 10012 23418 10036 23420
rect 10092 23418 10116 23420
rect 10172 23418 10196 23420
rect 10252 23418 10258 23420
rect 10012 23366 10014 23418
rect 10194 23366 10196 23418
rect 9950 23364 9956 23366
rect 10012 23364 10036 23366
rect 10092 23364 10116 23366
rect 10172 23364 10196 23366
rect 10252 23364 10258 23366
rect 9950 23355 10258 23364
rect 17950 23420 18258 23429
rect 17950 23418 17956 23420
rect 18012 23418 18036 23420
rect 18092 23418 18116 23420
rect 18172 23418 18196 23420
rect 18252 23418 18258 23420
rect 18012 23366 18014 23418
rect 18194 23366 18196 23418
rect 17950 23364 17956 23366
rect 18012 23364 18036 23366
rect 18092 23364 18116 23366
rect 18172 23364 18196 23366
rect 18252 23364 18258 23366
rect 17950 23355 18258 23364
rect 25950 23420 26258 23429
rect 25950 23418 25956 23420
rect 26012 23418 26036 23420
rect 26092 23418 26116 23420
rect 26172 23418 26196 23420
rect 26252 23418 26258 23420
rect 26012 23366 26014 23418
rect 26194 23366 26196 23418
rect 25950 23364 25956 23366
rect 26012 23364 26036 23366
rect 26092 23364 26116 23366
rect 26172 23364 26196 23366
rect 26252 23364 26258 23366
rect 25950 23355 26258 23364
rect 2610 22876 2918 22885
rect 2610 22874 2616 22876
rect 2672 22874 2696 22876
rect 2752 22874 2776 22876
rect 2832 22874 2856 22876
rect 2912 22874 2918 22876
rect 2672 22822 2674 22874
rect 2854 22822 2856 22874
rect 2610 22820 2616 22822
rect 2672 22820 2696 22822
rect 2752 22820 2776 22822
rect 2832 22820 2856 22822
rect 2912 22820 2918 22822
rect 2610 22811 2918 22820
rect 10610 22876 10918 22885
rect 10610 22874 10616 22876
rect 10672 22874 10696 22876
rect 10752 22874 10776 22876
rect 10832 22874 10856 22876
rect 10912 22874 10918 22876
rect 10672 22822 10674 22874
rect 10854 22822 10856 22874
rect 10610 22820 10616 22822
rect 10672 22820 10696 22822
rect 10752 22820 10776 22822
rect 10832 22820 10856 22822
rect 10912 22820 10918 22822
rect 10610 22811 10918 22820
rect 18610 22876 18918 22885
rect 18610 22874 18616 22876
rect 18672 22874 18696 22876
rect 18752 22874 18776 22876
rect 18832 22874 18856 22876
rect 18912 22874 18918 22876
rect 18672 22822 18674 22874
rect 18854 22822 18856 22874
rect 18610 22820 18616 22822
rect 18672 22820 18696 22822
rect 18752 22820 18776 22822
rect 18832 22820 18856 22822
rect 18912 22820 18918 22822
rect 18610 22811 18918 22820
rect 26610 22876 26918 22885
rect 26610 22874 26616 22876
rect 26672 22874 26696 22876
rect 26752 22874 26776 22876
rect 26832 22874 26856 22876
rect 26912 22874 26918 22876
rect 26672 22822 26674 22874
rect 26854 22822 26856 22874
rect 26610 22820 26616 22822
rect 26672 22820 26696 22822
rect 26752 22820 26776 22822
rect 26832 22820 26856 22822
rect 26912 22820 26918 22822
rect 26610 22811 26918 22820
rect 848 22636 900 22642
rect 848 22578 900 22584
rect 27436 22636 27488 22642
rect 27436 22578 27488 22584
rect 860 22545 888 22578
rect 846 22536 902 22545
rect 846 22471 902 22480
rect 1768 22432 1820 22438
rect 1768 22374 1820 22380
rect 1780 16998 1808 22374
rect 1950 22332 2258 22341
rect 1950 22330 1956 22332
rect 2012 22330 2036 22332
rect 2092 22330 2116 22332
rect 2172 22330 2196 22332
rect 2252 22330 2258 22332
rect 2012 22278 2014 22330
rect 2194 22278 2196 22330
rect 1950 22276 1956 22278
rect 2012 22276 2036 22278
rect 2092 22276 2116 22278
rect 2172 22276 2196 22278
rect 2252 22276 2258 22278
rect 1950 22267 2258 22276
rect 9950 22332 10258 22341
rect 9950 22330 9956 22332
rect 10012 22330 10036 22332
rect 10092 22330 10116 22332
rect 10172 22330 10196 22332
rect 10252 22330 10258 22332
rect 10012 22278 10014 22330
rect 10194 22278 10196 22330
rect 9950 22276 9956 22278
rect 10012 22276 10036 22278
rect 10092 22276 10116 22278
rect 10172 22276 10196 22278
rect 10252 22276 10258 22278
rect 9950 22267 10258 22276
rect 17950 22332 18258 22341
rect 17950 22330 17956 22332
rect 18012 22330 18036 22332
rect 18092 22330 18116 22332
rect 18172 22330 18196 22332
rect 18252 22330 18258 22332
rect 18012 22278 18014 22330
rect 18194 22278 18196 22330
rect 17950 22276 17956 22278
rect 18012 22276 18036 22278
rect 18092 22276 18116 22278
rect 18172 22276 18196 22278
rect 18252 22276 18258 22278
rect 17950 22267 18258 22276
rect 25950 22332 26258 22341
rect 25950 22330 25956 22332
rect 26012 22330 26036 22332
rect 26092 22330 26116 22332
rect 26172 22330 26196 22332
rect 26252 22330 26258 22332
rect 26012 22278 26014 22330
rect 26194 22278 26196 22330
rect 25950 22276 25956 22278
rect 26012 22276 26036 22278
rect 26092 22276 26116 22278
rect 26172 22276 26196 22278
rect 26252 22276 26258 22278
rect 25950 22267 26258 22276
rect 2610 21788 2918 21797
rect 2610 21786 2616 21788
rect 2672 21786 2696 21788
rect 2752 21786 2776 21788
rect 2832 21786 2856 21788
rect 2912 21786 2918 21788
rect 2672 21734 2674 21786
rect 2854 21734 2856 21786
rect 2610 21732 2616 21734
rect 2672 21732 2696 21734
rect 2752 21732 2776 21734
rect 2832 21732 2856 21734
rect 2912 21732 2918 21734
rect 2610 21723 2918 21732
rect 10610 21788 10918 21797
rect 10610 21786 10616 21788
rect 10672 21786 10696 21788
rect 10752 21786 10776 21788
rect 10832 21786 10856 21788
rect 10912 21786 10918 21788
rect 10672 21734 10674 21786
rect 10854 21734 10856 21786
rect 10610 21732 10616 21734
rect 10672 21732 10696 21734
rect 10752 21732 10776 21734
rect 10832 21732 10856 21734
rect 10912 21732 10918 21734
rect 10610 21723 10918 21732
rect 18610 21788 18918 21797
rect 18610 21786 18616 21788
rect 18672 21786 18696 21788
rect 18752 21786 18776 21788
rect 18832 21786 18856 21788
rect 18912 21786 18918 21788
rect 18672 21734 18674 21786
rect 18854 21734 18856 21786
rect 18610 21732 18616 21734
rect 18672 21732 18696 21734
rect 18752 21732 18776 21734
rect 18832 21732 18856 21734
rect 18912 21732 18918 21734
rect 18610 21723 18918 21732
rect 26610 21788 26918 21797
rect 26610 21786 26616 21788
rect 26672 21786 26696 21788
rect 26752 21786 26776 21788
rect 26832 21786 26856 21788
rect 26912 21786 26918 21788
rect 26672 21734 26674 21786
rect 26854 21734 26856 21786
rect 26610 21732 26616 21734
rect 26672 21732 26696 21734
rect 26752 21732 26776 21734
rect 26832 21732 26856 21734
rect 26912 21732 26918 21734
rect 26610 21723 26918 21732
rect 1950 21244 2258 21253
rect 1950 21242 1956 21244
rect 2012 21242 2036 21244
rect 2092 21242 2116 21244
rect 2172 21242 2196 21244
rect 2252 21242 2258 21244
rect 2012 21190 2014 21242
rect 2194 21190 2196 21242
rect 1950 21188 1956 21190
rect 2012 21188 2036 21190
rect 2092 21188 2116 21190
rect 2172 21188 2196 21190
rect 2252 21188 2258 21190
rect 1950 21179 2258 21188
rect 9950 21244 10258 21253
rect 9950 21242 9956 21244
rect 10012 21242 10036 21244
rect 10092 21242 10116 21244
rect 10172 21242 10196 21244
rect 10252 21242 10258 21244
rect 10012 21190 10014 21242
rect 10194 21190 10196 21242
rect 9950 21188 9956 21190
rect 10012 21188 10036 21190
rect 10092 21188 10116 21190
rect 10172 21188 10196 21190
rect 10252 21188 10258 21190
rect 9950 21179 10258 21188
rect 17950 21244 18258 21253
rect 17950 21242 17956 21244
rect 18012 21242 18036 21244
rect 18092 21242 18116 21244
rect 18172 21242 18196 21244
rect 18252 21242 18258 21244
rect 18012 21190 18014 21242
rect 18194 21190 18196 21242
rect 17950 21188 17956 21190
rect 18012 21188 18036 21190
rect 18092 21188 18116 21190
rect 18172 21188 18196 21190
rect 18252 21188 18258 21190
rect 17950 21179 18258 21188
rect 25950 21244 26258 21253
rect 25950 21242 25956 21244
rect 26012 21242 26036 21244
rect 26092 21242 26116 21244
rect 26172 21242 26196 21244
rect 26252 21242 26258 21244
rect 26012 21190 26014 21242
rect 26194 21190 26196 21242
rect 25950 21188 25956 21190
rect 26012 21188 26036 21190
rect 26092 21188 26116 21190
rect 26172 21188 26196 21190
rect 26252 21188 26258 21190
rect 25950 21179 26258 21188
rect 27448 20942 27476 22578
rect 27540 22030 27568 24142
rect 27528 22024 27580 22030
rect 27528 21966 27580 21972
rect 27436 20936 27488 20942
rect 27436 20878 27488 20884
rect 2610 20700 2918 20709
rect 2610 20698 2616 20700
rect 2672 20698 2696 20700
rect 2752 20698 2776 20700
rect 2832 20698 2856 20700
rect 2912 20698 2918 20700
rect 2672 20646 2674 20698
rect 2854 20646 2856 20698
rect 2610 20644 2616 20646
rect 2672 20644 2696 20646
rect 2752 20644 2776 20646
rect 2832 20644 2856 20646
rect 2912 20644 2918 20646
rect 2610 20635 2918 20644
rect 10610 20700 10918 20709
rect 10610 20698 10616 20700
rect 10672 20698 10696 20700
rect 10752 20698 10776 20700
rect 10832 20698 10856 20700
rect 10912 20698 10918 20700
rect 10672 20646 10674 20698
rect 10854 20646 10856 20698
rect 10610 20644 10616 20646
rect 10672 20644 10696 20646
rect 10752 20644 10776 20646
rect 10832 20644 10856 20646
rect 10912 20644 10918 20646
rect 10610 20635 10918 20644
rect 18610 20700 18918 20709
rect 18610 20698 18616 20700
rect 18672 20698 18696 20700
rect 18752 20698 18776 20700
rect 18832 20698 18856 20700
rect 18912 20698 18918 20700
rect 18672 20646 18674 20698
rect 18854 20646 18856 20698
rect 18610 20644 18616 20646
rect 18672 20644 18696 20646
rect 18752 20644 18776 20646
rect 18832 20644 18856 20646
rect 18912 20644 18918 20646
rect 18610 20635 18918 20644
rect 26610 20700 26918 20709
rect 26610 20698 26616 20700
rect 26672 20698 26696 20700
rect 26752 20698 26776 20700
rect 26832 20698 26856 20700
rect 26912 20698 26918 20700
rect 26672 20646 26674 20698
rect 26854 20646 26856 20698
rect 26610 20644 26616 20646
rect 26672 20644 26696 20646
rect 26752 20644 26776 20646
rect 26832 20644 26856 20646
rect 26912 20644 26918 20646
rect 26610 20635 26918 20644
rect 1950 20156 2258 20165
rect 1950 20154 1956 20156
rect 2012 20154 2036 20156
rect 2092 20154 2116 20156
rect 2172 20154 2196 20156
rect 2252 20154 2258 20156
rect 2012 20102 2014 20154
rect 2194 20102 2196 20154
rect 1950 20100 1956 20102
rect 2012 20100 2036 20102
rect 2092 20100 2116 20102
rect 2172 20100 2196 20102
rect 2252 20100 2258 20102
rect 1950 20091 2258 20100
rect 9950 20156 10258 20165
rect 9950 20154 9956 20156
rect 10012 20154 10036 20156
rect 10092 20154 10116 20156
rect 10172 20154 10196 20156
rect 10252 20154 10258 20156
rect 10012 20102 10014 20154
rect 10194 20102 10196 20154
rect 9950 20100 9956 20102
rect 10012 20100 10036 20102
rect 10092 20100 10116 20102
rect 10172 20100 10196 20102
rect 10252 20100 10258 20102
rect 9950 20091 10258 20100
rect 17950 20156 18258 20165
rect 17950 20154 17956 20156
rect 18012 20154 18036 20156
rect 18092 20154 18116 20156
rect 18172 20154 18196 20156
rect 18252 20154 18258 20156
rect 18012 20102 18014 20154
rect 18194 20102 18196 20154
rect 17950 20100 17956 20102
rect 18012 20100 18036 20102
rect 18092 20100 18116 20102
rect 18172 20100 18196 20102
rect 18252 20100 18258 20102
rect 17950 20091 18258 20100
rect 25950 20156 26258 20165
rect 25950 20154 25956 20156
rect 26012 20154 26036 20156
rect 26092 20154 26116 20156
rect 26172 20154 26196 20156
rect 26252 20154 26258 20156
rect 26012 20102 26014 20154
rect 26194 20102 26196 20154
rect 25950 20100 25956 20102
rect 26012 20100 26036 20102
rect 26092 20100 26116 20102
rect 26172 20100 26196 20102
rect 26252 20100 26258 20102
rect 25950 20091 26258 20100
rect 2610 19612 2918 19621
rect 2610 19610 2616 19612
rect 2672 19610 2696 19612
rect 2752 19610 2776 19612
rect 2832 19610 2856 19612
rect 2912 19610 2918 19612
rect 2672 19558 2674 19610
rect 2854 19558 2856 19610
rect 2610 19556 2616 19558
rect 2672 19556 2696 19558
rect 2752 19556 2776 19558
rect 2832 19556 2856 19558
rect 2912 19556 2918 19558
rect 2610 19547 2918 19556
rect 10610 19612 10918 19621
rect 10610 19610 10616 19612
rect 10672 19610 10696 19612
rect 10752 19610 10776 19612
rect 10832 19610 10856 19612
rect 10912 19610 10918 19612
rect 10672 19558 10674 19610
rect 10854 19558 10856 19610
rect 10610 19556 10616 19558
rect 10672 19556 10696 19558
rect 10752 19556 10776 19558
rect 10832 19556 10856 19558
rect 10912 19556 10918 19558
rect 10610 19547 10918 19556
rect 18610 19612 18918 19621
rect 18610 19610 18616 19612
rect 18672 19610 18696 19612
rect 18752 19610 18776 19612
rect 18832 19610 18856 19612
rect 18912 19610 18918 19612
rect 18672 19558 18674 19610
rect 18854 19558 18856 19610
rect 18610 19556 18616 19558
rect 18672 19556 18696 19558
rect 18752 19556 18776 19558
rect 18832 19556 18856 19558
rect 18912 19556 18918 19558
rect 18610 19547 18918 19556
rect 26610 19612 26918 19621
rect 26610 19610 26616 19612
rect 26672 19610 26696 19612
rect 26752 19610 26776 19612
rect 26832 19610 26856 19612
rect 26912 19610 26918 19612
rect 26672 19558 26674 19610
rect 26854 19558 26856 19610
rect 26610 19556 26616 19558
rect 26672 19556 26696 19558
rect 26752 19556 26776 19558
rect 26832 19556 26856 19558
rect 26912 19556 26918 19558
rect 26610 19547 26918 19556
rect 1950 19068 2258 19077
rect 1950 19066 1956 19068
rect 2012 19066 2036 19068
rect 2092 19066 2116 19068
rect 2172 19066 2196 19068
rect 2252 19066 2258 19068
rect 2012 19014 2014 19066
rect 2194 19014 2196 19066
rect 1950 19012 1956 19014
rect 2012 19012 2036 19014
rect 2092 19012 2116 19014
rect 2172 19012 2196 19014
rect 2252 19012 2258 19014
rect 1950 19003 2258 19012
rect 9950 19068 10258 19077
rect 9950 19066 9956 19068
rect 10012 19066 10036 19068
rect 10092 19066 10116 19068
rect 10172 19066 10196 19068
rect 10252 19066 10258 19068
rect 10012 19014 10014 19066
rect 10194 19014 10196 19066
rect 9950 19012 9956 19014
rect 10012 19012 10036 19014
rect 10092 19012 10116 19014
rect 10172 19012 10196 19014
rect 10252 19012 10258 19014
rect 9950 19003 10258 19012
rect 17950 19068 18258 19077
rect 17950 19066 17956 19068
rect 18012 19066 18036 19068
rect 18092 19066 18116 19068
rect 18172 19066 18196 19068
rect 18252 19066 18258 19068
rect 18012 19014 18014 19066
rect 18194 19014 18196 19066
rect 17950 19012 17956 19014
rect 18012 19012 18036 19014
rect 18092 19012 18116 19014
rect 18172 19012 18196 19014
rect 18252 19012 18258 19014
rect 17950 19003 18258 19012
rect 25950 19068 26258 19077
rect 25950 19066 25956 19068
rect 26012 19066 26036 19068
rect 26092 19066 26116 19068
rect 26172 19066 26196 19068
rect 26252 19066 26258 19068
rect 26012 19014 26014 19066
rect 26194 19014 26196 19066
rect 25950 19012 25956 19014
rect 26012 19012 26036 19014
rect 26092 19012 26116 19014
rect 26172 19012 26196 19014
rect 26252 19012 26258 19014
rect 25950 19003 26258 19012
rect 2610 18524 2918 18533
rect 2610 18522 2616 18524
rect 2672 18522 2696 18524
rect 2752 18522 2776 18524
rect 2832 18522 2856 18524
rect 2912 18522 2918 18524
rect 2672 18470 2674 18522
rect 2854 18470 2856 18522
rect 2610 18468 2616 18470
rect 2672 18468 2696 18470
rect 2752 18468 2776 18470
rect 2832 18468 2856 18470
rect 2912 18468 2918 18470
rect 2610 18459 2918 18468
rect 10610 18524 10918 18533
rect 10610 18522 10616 18524
rect 10672 18522 10696 18524
rect 10752 18522 10776 18524
rect 10832 18522 10856 18524
rect 10912 18522 10918 18524
rect 10672 18470 10674 18522
rect 10854 18470 10856 18522
rect 10610 18468 10616 18470
rect 10672 18468 10696 18470
rect 10752 18468 10776 18470
rect 10832 18468 10856 18470
rect 10912 18468 10918 18470
rect 10610 18459 10918 18468
rect 18610 18524 18918 18533
rect 18610 18522 18616 18524
rect 18672 18522 18696 18524
rect 18752 18522 18776 18524
rect 18832 18522 18856 18524
rect 18912 18522 18918 18524
rect 18672 18470 18674 18522
rect 18854 18470 18856 18522
rect 18610 18468 18616 18470
rect 18672 18468 18696 18470
rect 18752 18468 18776 18470
rect 18832 18468 18856 18470
rect 18912 18468 18918 18470
rect 18610 18459 18918 18468
rect 26610 18524 26918 18533
rect 26610 18522 26616 18524
rect 26672 18522 26696 18524
rect 26752 18522 26776 18524
rect 26832 18522 26856 18524
rect 26912 18522 26918 18524
rect 26672 18470 26674 18522
rect 26854 18470 26856 18522
rect 26610 18468 26616 18470
rect 26672 18468 26696 18470
rect 26752 18468 26776 18470
rect 26832 18468 26856 18470
rect 26912 18468 26918 18470
rect 26610 18459 26918 18468
rect 27344 18284 27396 18290
rect 27344 18226 27396 18232
rect 1950 17980 2258 17989
rect 1950 17978 1956 17980
rect 2012 17978 2036 17980
rect 2092 17978 2116 17980
rect 2172 17978 2196 17980
rect 2252 17978 2258 17980
rect 2012 17926 2014 17978
rect 2194 17926 2196 17978
rect 1950 17924 1956 17926
rect 2012 17924 2036 17926
rect 2092 17924 2116 17926
rect 2172 17924 2196 17926
rect 2252 17924 2258 17926
rect 1950 17915 2258 17924
rect 9950 17980 10258 17989
rect 9950 17978 9956 17980
rect 10012 17978 10036 17980
rect 10092 17978 10116 17980
rect 10172 17978 10196 17980
rect 10252 17978 10258 17980
rect 10012 17926 10014 17978
rect 10194 17926 10196 17978
rect 9950 17924 9956 17926
rect 10012 17924 10036 17926
rect 10092 17924 10116 17926
rect 10172 17924 10196 17926
rect 10252 17924 10258 17926
rect 9950 17915 10258 17924
rect 17950 17980 18258 17989
rect 17950 17978 17956 17980
rect 18012 17978 18036 17980
rect 18092 17978 18116 17980
rect 18172 17978 18196 17980
rect 18252 17978 18258 17980
rect 18012 17926 18014 17978
rect 18194 17926 18196 17978
rect 17950 17924 17956 17926
rect 18012 17924 18036 17926
rect 18092 17924 18116 17926
rect 18172 17924 18196 17926
rect 18252 17924 18258 17926
rect 17950 17915 18258 17924
rect 25950 17980 26258 17989
rect 25950 17978 25956 17980
rect 26012 17978 26036 17980
rect 26092 17978 26116 17980
rect 26172 17978 26196 17980
rect 26252 17978 26258 17980
rect 26012 17926 26014 17978
rect 26194 17926 26196 17978
rect 25950 17924 25956 17926
rect 26012 17924 26036 17926
rect 26092 17924 26116 17926
rect 26172 17924 26196 17926
rect 26252 17924 26258 17926
rect 25950 17915 26258 17924
rect 27356 17678 27384 18226
rect 27344 17672 27396 17678
rect 27344 17614 27396 17620
rect 2610 17436 2918 17445
rect 2610 17434 2616 17436
rect 2672 17434 2696 17436
rect 2752 17434 2776 17436
rect 2832 17434 2856 17436
rect 2912 17434 2918 17436
rect 2672 17382 2674 17434
rect 2854 17382 2856 17434
rect 2610 17380 2616 17382
rect 2672 17380 2696 17382
rect 2752 17380 2776 17382
rect 2832 17380 2856 17382
rect 2912 17380 2918 17382
rect 2610 17371 2918 17380
rect 10610 17436 10918 17445
rect 10610 17434 10616 17436
rect 10672 17434 10696 17436
rect 10752 17434 10776 17436
rect 10832 17434 10856 17436
rect 10912 17434 10918 17436
rect 10672 17382 10674 17434
rect 10854 17382 10856 17434
rect 10610 17380 10616 17382
rect 10672 17380 10696 17382
rect 10752 17380 10776 17382
rect 10832 17380 10856 17382
rect 10912 17380 10918 17382
rect 10610 17371 10918 17380
rect 18610 17436 18918 17445
rect 18610 17434 18616 17436
rect 18672 17434 18696 17436
rect 18752 17434 18776 17436
rect 18832 17434 18856 17436
rect 18912 17434 18918 17436
rect 18672 17382 18674 17434
rect 18854 17382 18856 17434
rect 18610 17380 18616 17382
rect 18672 17380 18696 17382
rect 18752 17380 18776 17382
rect 18832 17380 18856 17382
rect 18912 17380 18918 17382
rect 18610 17371 18918 17380
rect 26610 17436 26918 17445
rect 26610 17434 26616 17436
rect 26672 17434 26696 17436
rect 26752 17434 26776 17436
rect 26832 17434 26856 17436
rect 26912 17434 26918 17436
rect 26672 17382 26674 17434
rect 26854 17382 26856 17434
rect 26610 17380 26616 17382
rect 26672 17380 26696 17382
rect 26752 17380 26776 17382
rect 26832 17380 26856 17382
rect 26912 17380 26918 17382
rect 26610 17371 26918 17380
rect 26976 17128 27028 17134
rect 26976 17070 27028 17076
rect 26884 17060 26936 17066
rect 26884 17002 26936 17008
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1950 16892 2258 16901
rect 1950 16890 1956 16892
rect 2012 16890 2036 16892
rect 2092 16890 2116 16892
rect 2172 16890 2196 16892
rect 2252 16890 2258 16892
rect 2012 16838 2014 16890
rect 2194 16838 2196 16890
rect 1950 16836 1956 16838
rect 2012 16836 2036 16838
rect 2092 16836 2116 16838
rect 2172 16836 2196 16838
rect 2252 16836 2258 16838
rect 1950 16827 2258 16836
rect 9950 16892 10258 16901
rect 9950 16890 9956 16892
rect 10012 16890 10036 16892
rect 10092 16890 10116 16892
rect 10172 16890 10196 16892
rect 10252 16890 10258 16892
rect 10012 16838 10014 16890
rect 10194 16838 10196 16890
rect 9950 16836 9956 16838
rect 10012 16836 10036 16838
rect 10092 16836 10116 16838
rect 10172 16836 10196 16838
rect 10252 16836 10258 16838
rect 9950 16827 10258 16836
rect 17950 16892 18258 16901
rect 17950 16890 17956 16892
rect 18012 16890 18036 16892
rect 18092 16890 18116 16892
rect 18172 16890 18196 16892
rect 18252 16890 18258 16892
rect 18012 16838 18014 16890
rect 18194 16838 18196 16890
rect 17950 16836 17956 16838
rect 18012 16836 18036 16838
rect 18092 16836 18116 16838
rect 18172 16836 18196 16838
rect 18252 16836 18258 16838
rect 17950 16827 18258 16836
rect 25950 16892 26258 16901
rect 25950 16890 25956 16892
rect 26012 16890 26036 16892
rect 26092 16890 26116 16892
rect 26172 16890 26196 16892
rect 26252 16890 26258 16892
rect 26012 16838 26014 16890
rect 26194 16838 26196 16890
rect 25950 16836 25956 16838
rect 26012 16836 26036 16838
rect 26092 16836 26116 16838
rect 26172 16836 26196 16838
rect 26252 16836 26258 16838
rect 25950 16827 26258 16836
rect 26896 16658 26924 17002
rect 26988 16726 27016 17070
rect 27356 16794 27384 17614
rect 27448 17338 27476 20878
rect 27540 18766 27568 21966
rect 27528 18760 27580 18766
rect 27528 18702 27580 18708
rect 27436 17332 27488 17338
rect 27436 17274 27488 17280
rect 27344 16788 27396 16794
rect 27344 16730 27396 16736
rect 26976 16720 27028 16726
rect 26976 16662 27028 16668
rect 26884 16652 26936 16658
rect 26884 16594 26936 16600
rect 2610 16348 2918 16357
rect 2610 16346 2616 16348
rect 2672 16346 2696 16348
rect 2752 16346 2776 16348
rect 2832 16346 2856 16348
rect 2912 16346 2918 16348
rect 2672 16294 2674 16346
rect 2854 16294 2856 16346
rect 2610 16292 2616 16294
rect 2672 16292 2696 16294
rect 2752 16292 2776 16294
rect 2832 16292 2856 16294
rect 2912 16292 2918 16294
rect 2610 16283 2918 16292
rect 10610 16348 10918 16357
rect 10610 16346 10616 16348
rect 10672 16346 10696 16348
rect 10752 16346 10776 16348
rect 10832 16346 10856 16348
rect 10912 16346 10918 16348
rect 10672 16294 10674 16346
rect 10854 16294 10856 16346
rect 10610 16292 10616 16294
rect 10672 16292 10696 16294
rect 10752 16292 10776 16294
rect 10832 16292 10856 16294
rect 10912 16292 10918 16294
rect 10610 16283 10918 16292
rect 18610 16348 18918 16357
rect 18610 16346 18616 16348
rect 18672 16346 18696 16348
rect 18752 16346 18776 16348
rect 18832 16346 18856 16348
rect 18912 16346 18918 16348
rect 18672 16294 18674 16346
rect 18854 16294 18856 16346
rect 18610 16292 18616 16294
rect 18672 16292 18696 16294
rect 18752 16292 18776 16294
rect 18832 16292 18856 16294
rect 18912 16292 18918 16294
rect 18610 16283 18918 16292
rect 26610 16348 26918 16357
rect 26610 16346 26616 16348
rect 26672 16346 26696 16348
rect 26752 16346 26776 16348
rect 26832 16346 26856 16348
rect 26912 16346 26918 16348
rect 26672 16294 26674 16346
rect 26854 16294 26856 16346
rect 26610 16292 26616 16294
rect 26672 16292 26696 16294
rect 26752 16292 26776 16294
rect 26832 16292 26856 16294
rect 26912 16292 26918 16294
rect 26610 16283 26918 16292
rect 26988 16130 27016 16662
rect 27068 16652 27120 16658
rect 27068 16594 27120 16600
rect 27080 16266 27108 16594
rect 27080 16238 27200 16266
rect 27540 16250 27568 18702
rect 27632 18426 27660 27406
rect 28356 27396 28408 27402
rect 28356 27338 28408 27344
rect 28368 27033 28396 27338
rect 28354 27024 28410 27033
rect 28354 26959 28410 26968
rect 28080 25900 28132 25906
rect 28080 25842 28132 25848
rect 28092 24410 28120 25842
rect 28356 25832 28408 25838
rect 28356 25774 28408 25780
rect 28368 25401 28396 25774
rect 28354 25392 28410 25401
rect 28354 25327 28410 25336
rect 28080 24404 28132 24410
rect 28080 24346 28132 24352
rect 28080 24200 28132 24206
rect 28080 24142 28132 24148
rect 28092 22778 28120 24142
rect 28356 24132 28408 24138
rect 28356 24074 28408 24080
rect 28368 23769 28396 24074
rect 28354 23760 28410 23769
rect 28354 23695 28410 23704
rect 28080 22772 28132 22778
rect 28080 22714 28132 22720
rect 28080 22636 28132 22642
rect 28080 22578 28132 22584
rect 28092 22234 28120 22578
rect 28356 22568 28408 22574
rect 28356 22510 28408 22516
rect 28080 22228 28132 22234
rect 28080 22170 28132 22176
rect 28368 22137 28396 22510
rect 28354 22128 28410 22137
rect 28354 22063 28410 22072
rect 28356 20868 28408 20874
rect 28356 20810 28408 20816
rect 28368 20505 28396 20810
rect 28354 20496 28410 20505
rect 28354 20431 28410 20440
rect 28080 19372 28132 19378
rect 28080 19314 28132 19320
rect 28356 19372 28408 19378
rect 28356 19314 28408 19320
rect 28092 18970 28120 19314
rect 28080 18964 28132 18970
rect 28080 18906 28132 18912
rect 28368 18873 28396 19314
rect 28354 18864 28410 18873
rect 28354 18799 28410 18808
rect 27620 18420 27672 18426
rect 27620 18362 27672 18368
rect 28356 17604 28408 17610
rect 28356 17546 28408 17552
rect 28368 17241 28396 17546
rect 28354 17232 28410 17241
rect 28354 17167 28410 17176
rect 26988 16114 27108 16130
rect 26988 16108 27120 16114
rect 26988 16102 27068 16108
rect 27068 16050 27120 16056
rect 1950 15804 2258 15813
rect 1950 15802 1956 15804
rect 2012 15802 2036 15804
rect 2092 15802 2116 15804
rect 2172 15802 2196 15804
rect 2252 15802 2258 15804
rect 2012 15750 2014 15802
rect 2194 15750 2196 15802
rect 1950 15748 1956 15750
rect 2012 15748 2036 15750
rect 2092 15748 2116 15750
rect 2172 15748 2196 15750
rect 2252 15748 2258 15750
rect 1950 15739 2258 15748
rect 9950 15804 10258 15813
rect 9950 15802 9956 15804
rect 10012 15802 10036 15804
rect 10092 15802 10116 15804
rect 10172 15802 10196 15804
rect 10252 15802 10258 15804
rect 10012 15750 10014 15802
rect 10194 15750 10196 15802
rect 9950 15748 9956 15750
rect 10012 15748 10036 15750
rect 10092 15748 10116 15750
rect 10172 15748 10196 15750
rect 10252 15748 10258 15750
rect 9950 15739 10258 15748
rect 17950 15804 18258 15813
rect 17950 15802 17956 15804
rect 18012 15802 18036 15804
rect 18092 15802 18116 15804
rect 18172 15802 18196 15804
rect 18252 15802 18258 15804
rect 18012 15750 18014 15802
rect 18194 15750 18196 15802
rect 17950 15748 17956 15750
rect 18012 15748 18036 15750
rect 18092 15748 18116 15750
rect 18172 15748 18196 15750
rect 18252 15748 18258 15750
rect 17950 15739 18258 15748
rect 25950 15804 26258 15813
rect 25950 15802 25956 15804
rect 26012 15802 26036 15804
rect 26092 15802 26116 15804
rect 26172 15802 26196 15804
rect 26252 15802 26258 15804
rect 26012 15750 26014 15802
rect 26194 15750 26196 15802
rect 25950 15748 25956 15750
rect 26012 15748 26036 15750
rect 26092 15748 26116 15750
rect 26172 15748 26196 15750
rect 26252 15748 26258 15750
rect 25950 15739 26258 15748
rect 2610 15260 2918 15269
rect 2610 15258 2616 15260
rect 2672 15258 2696 15260
rect 2752 15258 2776 15260
rect 2832 15258 2856 15260
rect 2912 15258 2918 15260
rect 2672 15206 2674 15258
rect 2854 15206 2856 15258
rect 2610 15204 2616 15206
rect 2672 15204 2696 15206
rect 2752 15204 2776 15206
rect 2832 15204 2856 15206
rect 2912 15204 2918 15206
rect 2610 15195 2918 15204
rect 10610 15260 10918 15269
rect 10610 15258 10616 15260
rect 10672 15258 10696 15260
rect 10752 15258 10776 15260
rect 10832 15258 10856 15260
rect 10912 15258 10918 15260
rect 10672 15206 10674 15258
rect 10854 15206 10856 15258
rect 10610 15204 10616 15206
rect 10672 15204 10696 15206
rect 10752 15204 10776 15206
rect 10832 15204 10856 15206
rect 10912 15204 10918 15206
rect 10610 15195 10918 15204
rect 18610 15260 18918 15269
rect 18610 15258 18616 15260
rect 18672 15258 18696 15260
rect 18752 15258 18776 15260
rect 18832 15258 18856 15260
rect 18912 15258 18918 15260
rect 18672 15206 18674 15258
rect 18854 15206 18856 15258
rect 18610 15204 18616 15206
rect 18672 15204 18696 15206
rect 18752 15204 18776 15206
rect 18832 15204 18856 15206
rect 18912 15204 18918 15206
rect 18610 15195 18918 15204
rect 26610 15260 26918 15269
rect 26610 15258 26616 15260
rect 26672 15258 26696 15260
rect 26752 15258 26776 15260
rect 26832 15258 26856 15260
rect 26912 15258 26918 15260
rect 26672 15206 26674 15258
rect 26854 15206 26856 15258
rect 26610 15204 26616 15206
rect 26672 15204 26696 15206
rect 26752 15204 26776 15206
rect 26832 15204 26856 15206
rect 26912 15204 26918 15206
rect 26610 15195 26918 15204
rect 1950 14716 2258 14725
rect 1950 14714 1956 14716
rect 2012 14714 2036 14716
rect 2092 14714 2116 14716
rect 2172 14714 2196 14716
rect 2252 14714 2258 14716
rect 2012 14662 2014 14714
rect 2194 14662 2196 14714
rect 1950 14660 1956 14662
rect 2012 14660 2036 14662
rect 2092 14660 2116 14662
rect 2172 14660 2196 14662
rect 2252 14660 2258 14662
rect 1950 14651 2258 14660
rect 9950 14716 10258 14725
rect 9950 14714 9956 14716
rect 10012 14714 10036 14716
rect 10092 14714 10116 14716
rect 10172 14714 10196 14716
rect 10252 14714 10258 14716
rect 10012 14662 10014 14714
rect 10194 14662 10196 14714
rect 9950 14660 9956 14662
rect 10012 14660 10036 14662
rect 10092 14660 10116 14662
rect 10172 14660 10196 14662
rect 10252 14660 10258 14662
rect 9950 14651 10258 14660
rect 17950 14716 18258 14725
rect 17950 14714 17956 14716
rect 18012 14714 18036 14716
rect 18092 14714 18116 14716
rect 18172 14714 18196 14716
rect 18252 14714 18258 14716
rect 18012 14662 18014 14714
rect 18194 14662 18196 14714
rect 17950 14660 17956 14662
rect 18012 14660 18036 14662
rect 18092 14660 18116 14662
rect 18172 14660 18196 14662
rect 18252 14660 18258 14662
rect 17950 14651 18258 14660
rect 25950 14716 26258 14725
rect 25950 14714 25956 14716
rect 26012 14714 26036 14716
rect 26092 14714 26116 14716
rect 26172 14714 26196 14716
rect 26252 14714 26258 14716
rect 26012 14662 26014 14714
rect 26194 14662 26196 14714
rect 25950 14660 25956 14662
rect 26012 14660 26036 14662
rect 26092 14660 26116 14662
rect 26172 14660 26196 14662
rect 26252 14660 26258 14662
rect 25950 14651 26258 14660
rect 2610 14172 2918 14181
rect 2610 14170 2616 14172
rect 2672 14170 2696 14172
rect 2752 14170 2776 14172
rect 2832 14170 2856 14172
rect 2912 14170 2918 14172
rect 2672 14118 2674 14170
rect 2854 14118 2856 14170
rect 2610 14116 2616 14118
rect 2672 14116 2696 14118
rect 2752 14116 2776 14118
rect 2832 14116 2856 14118
rect 2912 14116 2918 14118
rect 2610 14107 2918 14116
rect 10610 14172 10918 14181
rect 10610 14170 10616 14172
rect 10672 14170 10696 14172
rect 10752 14170 10776 14172
rect 10832 14170 10856 14172
rect 10912 14170 10918 14172
rect 10672 14118 10674 14170
rect 10854 14118 10856 14170
rect 10610 14116 10616 14118
rect 10672 14116 10696 14118
rect 10752 14116 10776 14118
rect 10832 14116 10856 14118
rect 10912 14116 10918 14118
rect 10610 14107 10918 14116
rect 18610 14172 18918 14181
rect 18610 14170 18616 14172
rect 18672 14170 18696 14172
rect 18752 14170 18776 14172
rect 18832 14170 18856 14172
rect 18912 14170 18918 14172
rect 18672 14118 18674 14170
rect 18854 14118 18856 14170
rect 18610 14116 18616 14118
rect 18672 14116 18696 14118
rect 18752 14116 18776 14118
rect 18832 14116 18856 14118
rect 18912 14116 18918 14118
rect 18610 14107 18918 14116
rect 26610 14172 26918 14181
rect 26610 14170 26616 14172
rect 26672 14170 26696 14172
rect 26752 14170 26776 14172
rect 26832 14170 26856 14172
rect 26912 14170 26918 14172
rect 26672 14118 26674 14170
rect 26854 14118 26856 14170
rect 26610 14116 26616 14118
rect 26672 14116 26696 14118
rect 26752 14116 26776 14118
rect 26832 14116 26856 14118
rect 26912 14116 26918 14118
rect 26610 14107 26918 14116
rect 1950 13628 2258 13637
rect 1950 13626 1956 13628
rect 2012 13626 2036 13628
rect 2092 13626 2116 13628
rect 2172 13626 2196 13628
rect 2252 13626 2258 13628
rect 2012 13574 2014 13626
rect 2194 13574 2196 13626
rect 1950 13572 1956 13574
rect 2012 13572 2036 13574
rect 2092 13572 2116 13574
rect 2172 13572 2196 13574
rect 2252 13572 2258 13574
rect 1950 13563 2258 13572
rect 9950 13628 10258 13637
rect 9950 13626 9956 13628
rect 10012 13626 10036 13628
rect 10092 13626 10116 13628
rect 10172 13626 10196 13628
rect 10252 13626 10258 13628
rect 10012 13574 10014 13626
rect 10194 13574 10196 13626
rect 9950 13572 9956 13574
rect 10012 13572 10036 13574
rect 10092 13572 10116 13574
rect 10172 13572 10196 13574
rect 10252 13572 10258 13574
rect 9950 13563 10258 13572
rect 17950 13628 18258 13637
rect 17950 13626 17956 13628
rect 18012 13626 18036 13628
rect 18092 13626 18116 13628
rect 18172 13626 18196 13628
rect 18252 13626 18258 13628
rect 18012 13574 18014 13626
rect 18194 13574 18196 13626
rect 17950 13572 17956 13574
rect 18012 13572 18036 13574
rect 18092 13572 18116 13574
rect 18172 13572 18196 13574
rect 18252 13572 18258 13574
rect 17950 13563 18258 13572
rect 25950 13628 26258 13637
rect 25950 13626 25956 13628
rect 26012 13626 26036 13628
rect 26092 13626 26116 13628
rect 26172 13626 26196 13628
rect 26252 13626 26258 13628
rect 26012 13574 26014 13626
rect 26194 13574 26196 13626
rect 25950 13572 25956 13574
rect 26012 13572 26036 13574
rect 26092 13572 26116 13574
rect 26172 13572 26196 13574
rect 26252 13572 26258 13574
rect 25950 13563 26258 13572
rect 2610 13084 2918 13093
rect 2610 13082 2616 13084
rect 2672 13082 2696 13084
rect 2752 13082 2776 13084
rect 2832 13082 2856 13084
rect 2912 13082 2918 13084
rect 2672 13030 2674 13082
rect 2854 13030 2856 13082
rect 2610 13028 2616 13030
rect 2672 13028 2696 13030
rect 2752 13028 2776 13030
rect 2832 13028 2856 13030
rect 2912 13028 2918 13030
rect 2610 13019 2918 13028
rect 10610 13084 10918 13093
rect 10610 13082 10616 13084
rect 10672 13082 10696 13084
rect 10752 13082 10776 13084
rect 10832 13082 10856 13084
rect 10912 13082 10918 13084
rect 10672 13030 10674 13082
rect 10854 13030 10856 13082
rect 10610 13028 10616 13030
rect 10672 13028 10696 13030
rect 10752 13028 10776 13030
rect 10832 13028 10856 13030
rect 10912 13028 10918 13030
rect 10610 13019 10918 13028
rect 18610 13084 18918 13093
rect 18610 13082 18616 13084
rect 18672 13082 18696 13084
rect 18752 13082 18776 13084
rect 18832 13082 18856 13084
rect 18912 13082 18918 13084
rect 18672 13030 18674 13082
rect 18854 13030 18856 13082
rect 18610 13028 18616 13030
rect 18672 13028 18696 13030
rect 18752 13028 18776 13030
rect 18832 13028 18856 13030
rect 18912 13028 18918 13030
rect 18610 13019 18918 13028
rect 26610 13084 26918 13093
rect 26610 13082 26616 13084
rect 26672 13082 26696 13084
rect 26752 13082 26776 13084
rect 26832 13082 26856 13084
rect 26912 13082 26918 13084
rect 26672 13030 26674 13082
rect 26854 13030 26856 13082
rect 26610 13028 26616 13030
rect 26672 13028 26696 13030
rect 26752 13028 26776 13030
rect 26832 13028 26856 13030
rect 26912 13028 26918 13030
rect 26610 13019 26918 13028
rect 27080 12850 27108 16050
rect 27172 16046 27200 16238
rect 27528 16244 27580 16250
rect 27528 16186 27580 16192
rect 27160 16040 27212 16046
rect 27160 15982 27212 15988
rect 27172 12850 27200 15982
rect 27540 15502 27568 16186
rect 28354 15600 28410 15609
rect 28354 15535 28356 15544
rect 28408 15535 28410 15544
rect 28356 15506 28408 15512
rect 27528 15496 27580 15502
rect 27528 15438 27580 15444
rect 28080 14408 28132 14414
rect 28080 14350 28132 14356
rect 28092 13530 28120 14350
rect 28356 14340 28408 14346
rect 28356 14282 28408 14288
rect 28368 13977 28396 14282
rect 28354 13968 28410 13977
rect 28354 13903 28410 13912
rect 28080 13524 28132 13530
rect 28080 13466 28132 13472
rect 27620 13320 27672 13326
rect 27620 13262 27672 13268
rect 27068 12844 27120 12850
rect 27068 12786 27120 12792
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 1950 12540 2258 12549
rect 1950 12538 1956 12540
rect 2012 12538 2036 12540
rect 2092 12538 2116 12540
rect 2172 12538 2196 12540
rect 2252 12538 2258 12540
rect 2012 12486 2014 12538
rect 2194 12486 2196 12538
rect 1950 12484 1956 12486
rect 2012 12484 2036 12486
rect 2092 12484 2116 12486
rect 2172 12484 2196 12486
rect 2252 12484 2258 12486
rect 1950 12475 2258 12484
rect 9950 12540 10258 12549
rect 9950 12538 9956 12540
rect 10012 12538 10036 12540
rect 10092 12538 10116 12540
rect 10172 12538 10196 12540
rect 10252 12538 10258 12540
rect 10012 12486 10014 12538
rect 10194 12486 10196 12538
rect 9950 12484 9956 12486
rect 10012 12484 10036 12486
rect 10092 12484 10116 12486
rect 10172 12484 10196 12486
rect 10252 12484 10258 12486
rect 9950 12475 10258 12484
rect 17950 12540 18258 12549
rect 17950 12538 17956 12540
rect 18012 12538 18036 12540
rect 18092 12538 18116 12540
rect 18172 12538 18196 12540
rect 18252 12538 18258 12540
rect 18012 12486 18014 12538
rect 18194 12486 18196 12538
rect 17950 12484 17956 12486
rect 18012 12484 18036 12486
rect 18092 12484 18116 12486
rect 18172 12484 18196 12486
rect 18252 12484 18258 12486
rect 17950 12475 18258 12484
rect 25950 12540 26258 12549
rect 25950 12538 25956 12540
rect 26012 12538 26036 12540
rect 26092 12538 26116 12540
rect 26172 12538 26196 12540
rect 26252 12538 26258 12540
rect 26012 12486 26014 12538
rect 26194 12486 26196 12538
rect 25950 12484 25956 12486
rect 26012 12484 26036 12486
rect 26092 12484 26116 12486
rect 26172 12484 26196 12486
rect 26252 12484 26258 12486
rect 25950 12475 26258 12484
rect 2610 11996 2918 12005
rect 2610 11994 2616 11996
rect 2672 11994 2696 11996
rect 2752 11994 2776 11996
rect 2832 11994 2856 11996
rect 2912 11994 2918 11996
rect 2672 11942 2674 11994
rect 2854 11942 2856 11994
rect 2610 11940 2616 11942
rect 2672 11940 2696 11942
rect 2752 11940 2776 11942
rect 2832 11940 2856 11942
rect 2912 11940 2918 11942
rect 2610 11931 2918 11940
rect 10610 11996 10918 12005
rect 10610 11994 10616 11996
rect 10672 11994 10696 11996
rect 10752 11994 10776 11996
rect 10832 11994 10856 11996
rect 10912 11994 10918 11996
rect 10672 11942 10674 11994
rect 10854 11942 10856 11994
rect 10610 11940 10616 11942
rect 10672 11940 10696 11942
rect 10752 11940 10776 11942
rect 10832 11940 10856 11942
rect 10912 11940 10918 11942
rect 10610 11931 10918 11940
rect 18610 11996 18918 12005
rect 18610 11994 18616 11996
rect 18672 11994 18696 11996
rect 18752 11994 18776 11996
rect 18832 11994 18856 11996
rect 18912 11994 18918 11996
rect 18672 11942 18674 11994
rect 18854 11942 18856 11994
rect 18610 11940 18616 11942
rect 18672 11940 18696 11942
rect 18752 11940 18776 11942
rect 18832 11940 18856 11942
rect 18912 11940 18918 11942
rect 18610 11931 18918 11940
rect 26610 11996 26918 12005
rect 26610 11994 26616 11996
rect 26672 11994 26696 11996
rect 26752 11994 26776 11996
rect 26832 11994 26856 11996
rect 26912 11994 26918 11996
rect 26672 11942 26674 11994
rect 26854 11942 26856 11994
rect 26610 11940 26616 11942
rect 26672 11940 26696 11942
rect 26752 11940 26776 11942
rect 26832 11940 26856 11942
rect 26912 11940 26918 11942
rect 26610 11931 26918 11940
rect 1950 11452 2258 11461
rect 1950 11450 1956 11452
rect 2012 11450 2036 11452
rect 2092 11450 2116 11452
rect 2172 11450 2196 11452
rect 2252 11450 2258 11452
rect 2012 11398 2014 11450
rect 2194 11398 2196 11450
rect 1950 11396 1956 11398
rect 2012 11396 2036 11398
rect 2092 11396 2116 11398
rect 2172 11396 2196 11398
rect 2252 11396 2258 11398
rect 1950 11387 2258 11396
rect 9950 11452 10258 11461
rect 9950 11450 9956 11452
rect 10012 11450 10036 11452
rect 10092 11450 10116 11452
rect 10172 11450 10196 11452
rect 10252 11450 10258 11452
rect 10012 11398 10014 11450
rect 10194 11398 10196 11450
rect 9950 11396 9956 11398
rect 10012 11396 10036 11398
rect 10092 11396 10116 11398
rect 10172 11396 10196 11398
rect 10252 11396 10258 11398
rect 9950 11387 10258 11396
rect 17950 11452 18258 11461
rect 17950 11450 17956 11452
rect 18012 11450 18036 11452
rect 18092 11450 18116 11452
rect 18172 11450 18196 11452
rect 18252 11450 18258 11452
rect 18012 11398 18014 11450
rect 18194 11398 18196 11450
rect 17950 11396 17956 11398
rect 18012 11396 18036 11398
rect 18092 11396 18116 11398
rect 18172 11396 18196 11398
rect 18252 11396 18258 11398
rect 17950 11387 18258 11396
rect 25950 11452 26258 11461
rect 25950 11450 25956 11452
rect 26012 11450 26036 11452
rect 26092 11450 26116 11452
rect 26172 11450 26196 11452
rect 26252 11450 26258 11452
rect 26012 11398 26014 11450
rect 26194 11398 26196 11450
rect 25950 11396 25956 11398
rect 26012 11396 26036 11398
rect 26092 11396 26116 11398
rect 26172 11396 26196 11398
rect 26252 11396 26258 11398
rect 25950 11387 26258 11396
rect 2610 10908 2918 10917
rect 2610 10906 2616 10908
rect 2672 10906 2696 10908
rect 2752 10906 2776 10908
rect 2832 10906 2856 10908
rect 2912 10906 2918 10908
rect 2672 10854 2674 10906
rect 2854 10854 2856 10906
rect 2610 10852 2616 10854
rect 2672 10852 2696 10854
rect 2752 10852 2776 10854
rect 2832 10852 2856 10854
rect 2912 10852 2918 10854
rect 2610 10843 2918 10852
rect 10610 10908 10918 10917
rect 10610 10906 10616 10908
rect 10672 10906 10696 10908
rect 10752 10906 10776 10908
rect 10832 10906 10856 10908
rect 10912 10906 10918 10908
rect 10672 10854 10674 10906
rect 10854 10854 10856 10906
rect 10610 10852 10616 10854
rect 10672 10852 10696 10854
rect 10752 10852 10776 10854
rect 10832 10852 10856 10854
rect 10912 10852 10918 10854
rect 10610 10843 10918 10852
rect 18610 10908 18918 10917
rect 18610 10906 18616 10908
rect 18672 10906 18696 10908
rect 18752 10906 18776 10908
rect 18832 10906 18856 10908
rect 18912 10906 18918 10908
rect 18672 10854 18674 10906
rect 18854 10854 18856 10906
rect 18610 10852 18616 10854
rect 18672 10852 18696 10854
rect 18752 10852 18776 10854
rect 18832 10852 18856 10854
rect 18912 10852 18918 10854
rect 18610 10843 18918 10852
rect 26610 10908 26918 10917
rect 26610 10906 26616 10908
rect 26672 10906 26696 10908
rect 26752 10906 26776 10908
rect 26832 10906 26856 10908
rect 26912 10906 26918 10908
rect 26672 10854 26674 10906
rect 26854 10854 26856 10906
rect 26610 10852 26616 10854
rect 26672 10852 26696 10854
rect 26752 10852 26776 10854
rect 26832 10852 26856 10854
rect 26912 10852 26918 10854
rect 26610 10843 26918 10852
rect 27080 10674 27108 12786
rect 27172 12730 27200 12786
rect 27172 12702 27292 12730
rect 27264 10810 27292 12702
rect 27632 12646 27660 13262
rect 28080 12844 28132 12850
rect 28080 12786 28132 12792
rect 27620 12640 27672 12646
rect 27620 12582 27672 12588
rect 28092 11898 28120 12786
rect 28356 12776 28408 12782
rect 28356 12718 28408 12724
rect 28172 12640 28224 12646
rect 28172 12582 28224 12588
rect 28080 11892 28132 11898
rect 28080 11834 28132 11840
rect 27436 11756 27488 11762
rect 27436 11698 27488 11704
rect 27252 10804 27304 10810
rect 27252 10746 27304 10752
rect 27264 10674 27292 10746
rect 27448 10742 27476 11698
rect 28080 11144 28132 11150
rect 28080 11086 28132 11092
rect 27436 10736 27488 10742
rect 27436 10678 27488 10684
rect 26516 10668 26568 10674
rect 26516 10610 26568 10616
rect 27068 10668 27120 10674
rect 27068 10610 27120 10616
rect 27252 10668 27304 10674
rect 27252 10610 27304 10616
rect 1950 10364 2258 10373
rect 1950 10362 1956 10364
rect 2012 10362 2036 10364
rect 2092 10362 2116 10364
rect 2172 10362 2196 10364
rect 2252 10362 2258 10364
rect 2012 10310 2014 10362
rect 2194 10310 2196 10362
rect 1950 10308 1956 10310
rect 2012 10308 2036 10310
rect 2092 10308 2116 10310
rect 2172 10308 2196 10310
rect 2252 10308 2258 10310
rect 1950 10299 2258 10308
rect 9950 10364 10258 10373
rect 9950 10362 9956 10364
rect 10012 10362 10036 10364
rect 10092 10362 10116 10364
rect 10172 10362 10196 10364
rect 10252 10362 10258 10364
rect 10012 10310 10014 10362
rect 10194 10310 10196 10362
rect 9950 10308 9956 10310
rect 10012 10308 10036 10310
rect 10092 10308 10116 10310
rect 10172 10308 10196 10310
rect 10252 10308 10258 10310
rect 9950 10299 10258 10308
rect 17950 10364 18258 10373
rect 17950 10362 17956 10364
rect 18012 10362 18036 10364
rect 18092 10362 18116 10364
rect 18172 10362 18196 10364
rect 18252 10362 18258 10364
rect 18012 10310 18014 10362
rect 18194 10310 18196 10362
rect 17950 10308 17956 10310
rect 18012 10308 18036 10310
rect 18092 10308 18116 10310
rect 18172 10308 18196 10310
rect 18252 10308 18258 10310
rect 17950 10299 18258 10308
rect 25950 10364 26258 10373
rect 25950 10362 25956 10364
rect 26012 10362 26036 10364
rect 26092 10362 26116 10364
rect 26172 10362 26196 10364
rect 26252 10362 26258 10364
rect 26012 10310 26014 10362
rect 26194 10310 26196 10362
rect 25950 10308 25956 10310
rect 26012 10308 26036 10310
rect 26092 10308 26116 10310
rect 26172 10308 26196 10310
rect 26252 10308 26258 10310
rect 25950 10299 26258 10308
rect 2610 9820 2918 9829
rect 2610 9818 2616 9820
rect 2672 9818 2696 9820
rect 2752 9818 2776 9820
rect 2832 9818 2856 9820
rect 2912 9818 2918 9820
rect 2672 9766 2674 9818
rect 2854 9766 2856 9818
rect 2610 9764 2616 9766
rect 2672 9764 2696 9766
rect 2752 9764 2776 9766
rect 2832 9764 2856 9766
rect 2912 9764 2918 9766
rect 2610 9755 2918 9764
rect 10610 9820 10918 9829
rect 10610 9818 10616 9820
rect 10672 9818 10696 9820
rect 10752 9818 10776 9820
rect 10832 9818 10856 9820
rect 10912 9818 10918 9820
rect 10672 9766 10674 9818
rect 10854 9766 10856 9818
rect 10610 9764 10616 9766
rect 10672 9764 10696 9766
rect 10752 9764 10776 9766
rect 10832 9764 10856 9766
rect 10912 9764 10918 9766
rect 10610 9755 10918 9764
rect 18610 9820 18918 9829
rect 18610 9818 18616 9820
rect 18672 9818 18696 9820
rect 18752 9818 18776 9820
rect 18832 9818 18856 9820
rect 18912 9818 18918 9820
rect 18672 9766 18674 9818
rect 18854 9766 18856 9818
rect 18610 9764 18616 9766
rect 18672 9764 18696 9766
rect 18752 9764 18776 9766
rect 18832 9764 18856 9766
rect 18912 9764 18918 9766
rect 18610 9755 18918 9764
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 9950 9276 10258 9285
rect 9950 9274 9956 9276
rect 10012 9274 10036 9276
rect 10092 9274 10116 9276
rect 10172 9274 10196 9276
rect 10252 9274 10258 9276
rect 10012 9222 10014 9274
rect 10194 9222 10196 9274
rect 9950 9220 9956 9222
rect 10012 9220 10036 9222
rect 10092 9220 10116 9222
rect 10172 9220 10196 9222
rect 10252 9220 10258 9222
rect 9950 9211 10258 9220
rect 17950 9276 18258 9285
rect 17950 9274 17956 9276
rect 18012 9274 18036 9276
rect 18092 9274 18116 9276
rect 18172 9274 18196 9276
rect 18252 9274 18258 9276
rect 18012 9222 18014 9274
rect 18194 9222 18196 9274
rect 17950 9220 17956 9222
rect 18012 9220 18036 9222
rect 18092 9220 18116 9222
rect 18172 9220 18196 9222
rect 18252 9220 18258 9222
rect 17950 9211 18258 9220
rect 25950 9276 26258 9285
rect 25950 9274 25956 9276
rect 26012 9274 26036 9276
rect 26092 9274 26116 9276
rect 26172 9274 26196 9276
rect 26252 9274 26258 9276
rect 26012 9222 26014 9274
rect 26194 9222 26196 9274
rect 25950 9220 25956 9222
rect 26012 9220 26036 9222
rect 26092 9220 26116 9222
rect 26172 9220 26196 9222
rect 26252 9220 26258 9222
rect 25950 9211 26258 9220
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 10610 8732 10918 8741
rect 10610 8730 10616 8732
rect 10672 8730 10696 8732
rect 10752 8730 10776 8732
rect 10832 8730 10856 8732
rect 10912 8730 10918 8732
rect 10672 8678 10674 8730
rect 10854 8678 10856 8730
rect 10610 8676 10616 8678
rect 10672 8676 10696 8678
rect 10752 8676 10776 8678
rect 10832 8676 10856 8678
rect 10912 8676 10918 8678
rect 10610 8667 10918 8676
rect 18610 8732 18918 8741
rect 18610 8730 18616 8732
rect 18672 8730 18696 8732
rect 18752 8730 18776 8732
rect 18832 8730 18856 8732
rect 18912 8730 18918 8732
rect 18672 8678 18674 8730
rect 18854 8678 18856 8730
rect 18610 8676 18616 8678
rect 18672 8676 18696 8678
rect 18752 8676 18776 8678
rect 18832 8676 18856 8678
rect 18912 8676 18918 8678
rect 18610 8667 18918 8676
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 9950 8188 10258 8197
rect 9950 8186 9956 8188
rect 10012 8186 10036 8188
rect 10092 8186 10116 8188
rect 10172 8186 10196 8188
rect 10252 8186 10258 8188
rect 10012 8134 10014 8186
rect 10194 8134 10196 8186
rect 9950 8132 9956 8134
rect 10012 8132 10036 8134
rect 10092 8132 10116 8134
rect 10172 8132 10196 8134
rect 10252 8132 10258 8134
rect 9950 8123 10258 8132
rect 17950 8188 18258 8197
rect 17950 8186 17956 8188
rect 18012 8186 18036 8188
rect 18092 8186 18116 8188
rect 18172 8186 18196 8188
rect 18252 8186 18258 8188
rect 18012 8134 18014 8186
rect 18194 8134 18196 8186
rect 17950 8132 17956 8134
rect 18012 8132 18036 8134
rect 18092 8132 18116 8134
rect 18172 8132 18196 8134
rect 18252 8132 18258 8134
rect 17950 8123 18258 8132
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 848 7812 900 7818
rect 848 7754 900 7760
rect 860 7585 888 7754
rect 26528 7750 26556 10610
rect 26610 9820 26918 9829
rect 26610 9818 26616 9820
rect 26672 9818 26696 9820
rect 26752 9818 26776 9820
rect 26832 9818 26856 9820
rect 26912 9818 26918 9820
rect 26672 9766 26674 9818
rect 26854 9766 26856 9818
rect 26610 9764 26616 9766
rect 26672 9764 26696 9766
rect 26752 9764 26776 9766
rect 26832 9764 26856 9766
rect 26912 9764 26918 9766
rect 26610 9755 26918 9764
rect 27448 8974 27476 10678
rect 27528 10532 27580 10538
rect 27528 10474 27580 10480
rect 27540 9586 27568 10474
rect 27528 9580 27580 9586
rect 27528 9522 27580 9528
rect 27712 9580 27764 9586
rect 27712 9522 27764 9528
rect 27436 8968 27488 8974
rect 27436 8910 27488 8916
rect 26610 8732 26918 8741
rect 26610 8730 26616 8732
rect 26672 8730 26696 8732
rect 26752 8730 26776 8732
rect 26832 8730 26856 8732
rect 26912 8730 26918 8732
rect 26672 8678 26674 8730
rect 26854 8678 26856 8730
rect 26610 8676 26616 8678
rect 26672 8676 26696 8678
rect 26752 8676 26776 8678
rect 26832 8676 26856 8678
rect 26912 8676 26918 8678
rect 26610 8667 26918 8676
rect 26516 7744 26568 7750
rect 26516 7686 26568 7692
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 846 7576 902 7585
rect 2610 7579 2918 7588
rect 10610 7644 10918 7653
rect 10610 7642 10616 7644
rect 10672 7642 10696 7644
rect 10752 7642 10776 7644
rect 10832 7642 10856 7644
rect 10912 7642 10918 7644
rect 10672 7590 10674 7642
rect 10854 7590 10856 7642
rect 10610 7588 10616 7590
rect 10672 7588 10696 7590
rect 10752 7588 10776 7590
rect 10832 7588 10856 7590
rect 10912 7588 10918 7590
rect 10610 7579 10918 7588
rect 18610 7644 18918 7653
rect 18610 7642 18616 7644
rect 18672 7642 18696 7644
rect 18752 7642 18776 7644
rect 18832 7642 18856 7644
rect 18912 7642 18918 7644
rect 18672 7590 18674 7642
rect 18854 7590 18856 7642
rect 18610 7588 18616 7590
rect 18672 7588 18696 7590
rect 18752 7588 18776 7590
rect 18832 7588 18856 7590
rect 18912 7588 18918 7590
rect 18610 7579 18918 7588
rect 26610 7644 26918 7653
rect 26610 7642 26616 7644
rect 26672 7642 26696 7644
rect 26752 7642 26776 7644
rect 26832 7642 26856 7644
rect 26912 7642 26918 7644
rect 26672 7590 26674 7642
rect 26854 7590 26856 7642
rect 26610 7588 26616 7590
rect 26672 7588 26696 7590
rect 26752 7588 26776 7590
rect 26832 7588 26856 7590
rect 26912 7588 26918 7590
rect 26610 7579 26918 7588
rect 846 7511 902 7520
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 9950 7100 10258 7109
rect 9950 7098 9956 7100
rect 10012 7098 10036 7100
rect 10092 7098 10116 7100
rect 10172 7098 10196 7100
rect 10252 7098 10258 7100
rect 10012 7046 10014 7098
rect 10194 7046 10196 7098
rect 9950 7044 9956 7046
rect 10012 7044 10036 7046
rect 10092 7044 10116 7046
rect 10172 7044 10196 7046
rect 10252 7044 10258 7046
rect 9950 7035 10258 7044
rect 17950 7100 18258 7109
rect 17950 7098 17956 7100
rect 18012 7098 18036 7100
rect 18092 7098 18116 7100
rect 18172 7098 18196 7100
rect 18252 7098 18258 7100
rect 18012 7046 18014 7098
rect 18194 7046 18196 7098
rect 17950 7044 17956 7046
rect 18012 7044 18036 7046
rect 18092 7044 18116 7046
rect 18172 7044 18196 7046
rect 18252 7044 18258 7046
rect 17950 7035 18258 7044
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 27448 6914 27476 8910
rect 27540 7886 27568 9522
rect 27724 9178 27752 9522
rect 28092 9450 28120 11086
rect 28080 9444 28132 9450
rect 28080 9386 28132 9392
rect 27712 9172 27764 9178
rect 27712 9114 27764 9120
rect 27528 7880 27580 7886
rect 27528 7822 27580 7828
rect 27448 6886 27568 6914
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 10610 6556 10918 6565
rect 10610 6554 10616 6556
rect 10672 6554 10696 6556
rect 10752 6554 10776 6556
rect 10832 6554 10856 6556
rect 10912 6554 10918 6556
rect 10672 6502 10674 6554
rect 10854 6502 10856 6554
rect 10610 6500 10616 6502
rect 10672 6500 10696 6502
rect 10752 6500 10776 6502
rect 10832 6500 10856 6502
rect 10912 6500 10918 6502
rect 10610 6491 10918 6500
rect 18610 6556 18918 6565
rect 18610 6554 18616 6556
rect 18672 6554 18696 6556
rect 18752 6554 18776 6556
rect 18832 6554 18856 6556
rect 18912 6554 18918 6556
rect 18672 6502 18674 6554
rect 18854 6502 18856 6554
rect 18610 6500 18616 6502
rect 18672 6500 18696 6502
rect 18752 6500 18776 6502
rect 18832 6500 18856 6502
rect 18912 6500 18918 6502
rect 18610 6491 18918 6500
rect 26610 6556 26918 6565
rect 26610 6554 26616 6556
rect 26672 6554 26696 6556
rect 26752 6554 26776 6556
rect 26832 6554 26856 6556
rect 26912 6554 26918 6556
rect 26672 6502 26674 6554
rect 26854 6502 26856 6554
rect 26610 6500 26616 6502
rect 26672 6500 26696 6502
rect 26752 6500 26776 6502
rect 26832 6500 26856 6502
rect 26912 6500 26918 6502
rect 26610 6491 26918 6500
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 9950 6012 10258 6021
rect 9950 6010 9956 6012
rect 10012 6010 10036 6012
rect 10092 6010 10116 6012
rect 10172 6010 10196 6012
rect 10252 6010 10258 6012
rect 10012 5958 10014 6010
rect 10194 5958 10196 6010
rect 9950 5956 9956 5958
rect 10012 5956 10036 5958
rect 10092 5956 10116 5958
rect 10172 5956 10196 5958
rect 10252 5956 10258 5958
rect 9950 5947 10258 5956
rect 17950 6012 18258 6021
rect 17950 6010 17956 6012
rect 18012 6010 18036 6012
rect 18092 6010 18116 6012
rect 18172 6010 18196 6012
rect 18252 6010 18258 6012
rect 18012 5958 18014 6010
rect 18194 5958 18196 6010
rect 17950 5956 17956 5958
rect 18012 5956 18036 5958
rect 18092 5956 18116 5958
rect 18172 5956 18196 5958
rect 18252 5956 18258 5958
rect 17950 5947 18258 5956
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 27540 5710 27568 6886
rect 27712 6316 27764 6322
rect 27712 6258 27764 6264
rect 27724 5914 27752 6258
rect 27712 5908 27764 5914
rect 27712 5850 27764 5856
rect 27528 5704 27580 5710
rect 27528 5646 27580 5652
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 10610 5468 10918 5477
rect 10610 5466 10616 5468
rect 10672 5466 10696 5468
rect 10752 5466 10776 5468
rect 10832 5466 10856 5468
rect 10912 5466 10918 5468
rect 10672 5414 10674 5466
rect 10854 5414 10856 5466
rect 10610 5412 10616 5414
rect 10672 5412 10696 5414
rect 10752 5412 10776 5414
rect 10832 5412 10856 5414
rect 10912 5412 10918 5414
rect 10610 5403 10918 5412
rect 18610 5468 18918 5477
rect 18610 5466 18616 5468
rect 18672 5466 18696 5468
rect 18752 5466 18776 5468
rect 18832 5466 18856 5468
rect 18912 5466 18918 5468
rect 18672 5414 18674 5466
rect 18854 5414 18856 5466
rect 18610 5412 18616 5414
rect 18672 5412 18696 5414
rect 18752 5412 18776 5414
rect 18832 5412 18856 5414
rect 18912 5412 18918 5414
rect 18610 5403 18918 5412
rect 26610 5468 26918 5477
rect 26610 5466 26616 5468
rect 26672 5466 26696 5468
rect 26752 5466 26776 5468
rect 26832 5466 26856 5468
rect 26912 5466 26918 5468
rect 26672 5414 26674 5466
rect 26854 5414 26856 5466
rect 26610 5412 26616 5414
rect 26672 5412 26696 5414
rect 26752 5412 26776 5414
rect 26832 5412 26856 5414
rect 26912 5412 26918 5414
rect 26610 5403 26918 5412
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 9950 4924 10258 4933
rect 9950 4922 9956 4924
rect 10012 4922 10036 4924
rect 10092 4922 10116 4924
rect 10172 4922 10196 4924
rect 10252 4922 10258 4924
rect 10012 4870 10014 4922
rect 10194 4870 10196 4922
rect 9950 4868 9956 4870
rect 10012 4868 10036 4870
rect 10092 4868 10116 4870
rect 10172 4868 10196 4870
rect 10252 4868 10258 4870
rect 9950 4859 10258 4868
rect 17950 4924 18258 4933
rect 17950 4922 17956 4924
rect 18012 4922 18036 4924
rect 18092 4922 18116 4924
rect 18172 4922 18196 4924
rect 18252 4922 18258 4924
rect 18012 4870 18014 4922
rect 18194 4870 18196 4922
rect 17950 4868 17956 4870
rect 18012 4868 18036 4870
rect 18092 4868 18116 4870
rect 18172 4868 18196 4870
rect 18252 4868 18258 4870
rect 17950 4859 18258 4868
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 10610 4380 10918 4389
rect 10610 4378 10616 4380
rect 10672 4378 10696 4380
rect 10752 4378 10776 4380
rect 10832 4378 10856 4380
rect 10912 4378 10918 4380
rect 10672 4326 10674 4378
rect 10854 4326 10856 4378
rect 10610 4324 10616 4326
rect 10672 4324 10696 4326
rect 10752 4324 10776 4326
rect 10832 4324 10856 4326
rect 10912 4324 10918 4326
rect 10610 4315 10918 4324
rect 18610 4380 18918 4389
rect 18610 4378 18616 4380
rect 18672 4378 18696 4380
rect 18752 4378 18776 4380
rect 18832 4378 18856 4380
rect 18912 4378 18918 4380
rect 18672 4326 18674 4378
rect 18854 4326 18856 4378
rect 18610 4324 18616 4326
rect 18672 4324 18696 4326
rect 18752 4324 18776 4326
rect 18832 4324 18856 4326
rect 18912 4324 18918 4326
rect 18610 4315 18918 4324
rect 26610 4380 26918 4389
rect 26610 4378 26616 4380
rect 26672 4378 26696 4380
rect 26752 4378 26776 4380
rect 26832 4378 26856 4380
rect 26912 4378 26918 4380
rect 26672 4326 26674 4378
rect 26854 4326 26856 4378
rect 26610 4324 26616 4326
rect 26672 4324 26696 4326
rect 26752 4324 26776 4326
rect 26832 4324 26856 4326
rect 26912 4324 26918 4326
rect 26610 4315 26918 4324
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 9950 3836 10258 3845
rect 9950 3834 9956 3836
rect 10012 3834 10036 3836
rect 10092 3834 10116 3836
rect 10172 3834 10196 3836
rect 10252 3834 10258 3836
rect 10012 3782 10014 3834
rect 10194 3782 10196 3834
rect 9950 3780 9956 3782
rect 10012 3780 10036 3782
rect 10092 3780 10116 3782
rect 10172 3780 10196 3782
rect 10252 3780 10258 3782
rect 9950 3771 10258 3780
rect 17950 3836 18258 3845
rect 17950 3834 17956 3836
rect 18012 3834 18036 3836
rect 18092 3834 18116 3836
rect 18172 3834 18196 3836
rect 18252 3834 18258 3836
rect 18012 3782 18014 3834
rect 18194 3782 18196 3834
rect 17950 3780 17956 3782
rect 18012 3780 18036 3782
rect 18092 3780 18116 3782
rect 18172 3780 18196 3782
rect 18252 3780 18258 3782
rect 17950 3771 18258 3780
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 10610 3292 10918 3301
rect 10610 3290 10616 3292
rect 10672 3290 10696 3292
rect 10752 3290 10776 3292
rect 10832 3290 10856 3292
rect 10912 3290 10918 3292
rect 10672 3238 10674 3290
rect 10854 3238 10856 3290
rect 10610 3236 10616 3238
rect 10672 3236 10696 3238
rect 10752 3236 10776 3238
rect 10832 3236 10856 3238
rect 10912 3236 10918 3238
rect 10610 3227 10918 3236
rect 18610 3292 18918 3301
rect 18610 3290 18616 3292
rect 18672 3290 18696 3292
rect 18752 3290 18776 3292
rect 18832 3290 18856 3292
rect 18912 3290 18918 3292
rect 18672 3238 18674 3290
rect 18854 3238 18856 3290
rect 18610 3236 18616 3238
rect 18672 3236 18696 3238
rect 18752 3236 18776 3238
rect 18832 3236 18856 3238
rect 18912 3236 18918 3238
rect 18610 3227 18918 3236
rect 26610 3292 26918 3301
rect 26610 3290 26616 3292
rect 26672 3290 26696 3292
rect 26752 3290 26776 3292
rect 26832 3290 26856 3292
rect 26912 3290 26918 3292
rect 26672 3238 26674 3290
rect 26854 3238 26856 3290
rect 26610 3236 26616 3238
rect 26672 3236 26696 3238
rect 26752 3236 26776 3238
rect 26832 3236 26856 3238
rect 26912 3236 26918 3238
rect 26610 3227 26918 3236
rect 27540 3058 27568 5646
rect 28184 4622 28212 12582
rect 28368 12345 28396 12718
rect 28354 12336 28410 12345
rect 28354 12271 28410 12280
rect 28356 11076 28408 11082
rect 28356 11018 28408 11024
rect 28368 10713 28396 11018
rect 28354 10704 28410 10713
rect 28354 10639 28410 10648
rect 28356 9512 28408 9518
rect 28356 9454 28408 9460
rect 28368 9081 28396 9454
rect 28354 9072 28410 9081
rect 28354 9007 28410 9016
rect 28356 7812 28408 7818
rect 28356 7754 28408 7760
rect 28368 7449 28396 7754
rect 28354 7440 28410 7449
rect 28354 7375 28410 7384
rect 28356 6248 28408 6254
rect 28356 6190 28408 6196
rect 28368 5817 28396 6190
rect 28354 5808 28410 5817
rect 28354 5743 28410 5752
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 28356 4548 28408 4554
rect 28356 4490 28408 4496
rect 28368 4185 28396 4490
rect 28354 4176 28410 4185
rect 28354 4111 28410 4120
rect 27528 3052 27580 3058
rect 27528 2994 27580 3000
rect 28356 2984 28408 2990
rect 28356 2926 28408 2932
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 9950 2748 10258 2757
rect 9950 2746 9956 2748
rect 10012 2746 10036 2748
rect 10092 2746 10116 2748
rect 10172 2746 10196 2748
rect 10252 2746 10258 2748
rect 10012 2694 10014 2746
rect 10194 2694 10196 2746
rect 9950 2692 9956 2694
rect 10012 2692 10036 2694
rect 10092 2692 10116 2694
rect 10172 2692 10196 2694
rect 10252 2692 10258 2694
rect 9950 2683 10258 2692
rect 17950 2748 18258 2757
rect 17950 2746 17956 2748
rect 18012 2746 18036 2748
rect 18092 2746 18116 2748
rect 18172 2746 18196 2748
rect 18252 2746 18258 2748
rect 18012 2694 18014 2746
rect 18194 2694 18196 2746
rect 17950 2692 17956 2694
rect 18012 2692 18036 2694
rect 18092 2692 18116 2694
rect 18172 2692 18196 2694
rect 18252 2692 18258 2694
rect 17950 2683 18258 2692
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 28368 2553 28396 2926
rect 28354 2544 28410 2553
rect 28354 2479 28410 2488
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 10610 2204 10918 2213
rect 10610 2202 10616 2204
rect 10672 2202 10696 2204
rect 10752 2202 10776 2204
rect 10832 2202 10856 2204
rect 10912 2202 10918 2204
rect 10672 2150 10674 2202
rect 10854 2150 10856 2202
rect 10610 2148 10616 2150
rect 10672 2148 10696 2150
rect 10752 2148 10776 2150
rect 10832 2148 10856 2150
rect 10912 2148 10918 2150
rect 10610 2139 10918 2148
rect 18610 2204 18918 2213
rect 18610 2202 18616 2204
rect 18672 2202 18696 2204
rect 18752 2202 18776 2204
rect 18832 2202 18856 2204
rect 18912 2202 18918 2204
rect 18672 2150 18674 2202
rect 18854 2150 18856 2202
rect 18610 2148 18616 2150
rect 18672 2148 18696 2150
rect 18752 2148 18776 2150
rect 18832 2148 18856 2150
rect 18912 2148 18918 2150
rect 18610 2139 18918 2148
rect 26610 2204 26918 2213
rect 26610 2202 26616 2204
rect 26672 2202 26696 2204
rect 26752 2202 26776 2204
rect 26832 2202 26856 2204
rect 26912 2202 26918 2204
rect 26672 2150 26674 2202
rect 26854 2150 26856 2202
rect 26610 2148 26616 2150
rect 26672 2148 26696 2150
rect 26752 2148 26776 2150
rect 26832 2148 26856 2150
rect 26912 2148 26918 2150
rect 26610 2139 26918 2148
<< via2 >>
rect 1956 27770 2012 27772
rect 2036 27770 2092 27772
rect 2116 27770 2172 27772
rect 2196 27770 2252 27772
rect 1956 27718 2002 27770
rect 2002 27718 2012 27770
rect 2036 27718 2066 27770
rect 2066 27718 2078 27770
rect 2078 27718 2092 27770
rect 2116 27718 2130 27770
rect 2130 27718 2142 27770
rect 2142 27718 2172 27770
rect 2196 27718 2206 27770
rect 2206 27718 2252 27770
rect 1956 27716 2012 27718
rect 2036 27716 2092 27718
rect 2116 27716 2172 27718
rect 2196 27716 2252 27718
rect 9956 27770 10012 27772
rect 10036 27770 10092 27772
rect 10116 27770 10172 27772
rect 10196 27770 10252 27772
rect 9956 27718 10002 27770
rect 10002 27718 10012 27770
rect 10036 27718 10066 27770
rect 10066 27718 10078 27770
rect 10078 27718 10092 27770
rect 10116 27718 10130 27770
rect 10130 27718 10142 27770
rect 10142 27718 10172 27770
rect 10196 27718 10206 27770
rect 10206 27718 10252 27770
rect 9956 27716 10012 27718
rect 10036 27716 10092 27718
rect 10116 27716 10172 27718
rect 10196 27716 10252 27718
rect 17956 27770 18012 27772
rect 18036 27770 18092 27772
rect 18116 27770 18172 27772
rect 18196 27770 18252 27772
rect 17956 27718 18002 27770
rect 18002 27718 18012 27770
rect 18036 27718 18066 27770
rect 18066 27718 18078 27770
rect 18078 27718 18092 27770
rect 18116 27718 18130 27770
rect 18130 27718 18142 27770
rect 18142 27718 18172 27770
rect 18196 27718 18206 27770
rect 18206 27718 18252 27770
rect 17956 27716 18012 27718
rect 18036 27716 18092 27718
rect 18116 27716 18172 27718
rect 18196 27716 18252 27718
rect 25956 27770 26012 27772
rect 26036 27770 26092 27772
rect 26116 27770 26172 27772
rect 26196 27770 26252 27772
rect 25956 27718 26002 27770
rect 26002 27718 26012 27770
rect 26036 27718 26066 27770
rect 26066 27718 26078 27770
rect 26078 27718 26092 27770
rect 26116 27718 26130 27770
rect 26130 27718 26142 27770
rect 26142 27718 26172 27770
rect 26196 27718 26206 27770
rect 26206 27718 26252 27770
rect 25956 27716 26012 27718
rect 26036 27716 26092 27718
rect 26116 27716 26172 27718
rect 26196 27716 26252 27718
rect 2616 27226 2672 27228
rect 2696 27226 2752 27228
rect 2776 27226 2832 27228
rect 2856 27226 2912 27228
rect 2616 27174 2662 27226
rect 2662 27174 2672 27226
rect 2696 27174 2726 27226
rect 2726 27174 2738 27226
rect 2738 27174 2752 27226
rect 2776 27174 2790 27226
rect 2790 27174 2802 27226
rect 2802 27174 2832 27226
rect 2856 27174 2866 27226
rect 2866 27174 2912 27226
rect 2616 27172 2672 27174
rect 2696 27172 2752 27174
rect 2776 27172 2832 27174
rect 2856 27172 2912 27174
rect 10616 27226 10672 27228
rect 10696 27226 10752 27228
rect 10776 27226 10832 27228
rect 10856 27226 10912 27228
rect 10616 27174 10662 27226
rect 10662 27174 10672 27226
rect 10696 27174 10726 27226
rect 10726 27174 10738 27226
rect 10738 27174 10752 27226
rect 10776 27174 10790 27226
rect 10790 27174 10802 27226
rect 10802 27174 10832 27226
rect 10856 27174 10866 27226
rect 10866 27174 10912 27226
rect 10616 27172 10672 27174
rect 10696 27172 10752 27174
rect 10776 27172 10832 27174
rect 10856 27172 10912 27174
rect 18616 27226 18672 27228
rect 18696 27226 18752 27228
rect 18776 27226 18832 27228
rect 18856 27226 18912 27228
rect 18616 27174 18662 27226
rect 18662 27174 18672 27226
rect 18696 27174 18726 27226
rect 18726 27174 18738 27226
rect 18738 27174 18752 27226
rect 18776 27174 18790 27226
rect 18790 27174 18802 27226
rect 18802 27174 18832 27226
rect 18856 27174 18866 27226
rect 18866 27174 18912 27226
rect 18616 27172 18672 27174
rect 18696 27172 18752 27174
rect 18776 27172 18832 27174
rect 18856 27172 18912 27174
rect 26616 27226 26672 27228
rect 26696 27226 26752 27228
rect 26776 27226 26832 27228
rect 26856 27226 26912 27228
rect 26616 27174 26662 27226
rect 26662 27174 26672 27226
rect 26696 27174 26726 27226
rect 26726 27174 26738 27226
rect 26738 27174 26752 27226
rect 26776 27174 26790 27226
rect 26790 27174 26802 27226
rect 26802 27174 26832 27226
rect 26856 27174 26866 27226
rect 26866 27174 26912 27226
rect 26616 27172 26672 27174
rect 26696 27172 26752 27174
rect 26776 27172 26832 27174
rect 26856 27172 26912 27174
rect 1956 26682 2012 26684
rect 2036 26682 2092 26684
rect 2116 26682 2172 26684
rect 2196 26682 2252 26684
rect 1956 26630 2002 26682
rect 2002 26630 2012 26682
rect 2036 26630 2066 26682
rect 2066 26630 2078 26682
rect 2078 26630 2092 26682
rect 2116 26630 2130 26682
rect 2130 26630 2142 26682
rect 2142 26630 2172 26682
rect 2196 26630 2206 26682
rect 2206 26630 2252 26682
rect 1956 26628 2012 26630
rect 2036 26628 2092 26630
rect 2116 26628 2172 26630
rect 2196 26628 2252 26630
rect 9956 26682 10012 26684
rect 10036 26682 10092 26684
rect 10116 26682 10172 26684
rect 10196 26682 10252 26684
rect 9956 26630 10002 26682
rect 10002 26630 10012 26682
rect 10036 26630 10066 26682
rect 10066 26630 10078 26682
rect 10078 26630 10092 26682
rect 10116 26630 10130 26682
rect 10130 26630 10142 26682
rect 10142 26630 10172 26682
rect 10196 26630 10206 26682
rect 10206 26630 10252 26682
rect 9956 26628 10012 26630
rect 10036 26628 10092 26630
rect 10116 26628 10172 26630
rect 10196 26628 10252 26630
rect 17956 26682 18012 26684
rect 18036 26682 18092 26684
rect 18116 26682 18172 26684
rect 18196 26682 18252 26684
rect 17956 26630 18002 26682
rect 18002 26630 18012 26682
rect 18036 26630 18066 26682
rect 18066 26630 18078 26682
rect 18078 26630 18092 26682
rect 18116 26630 18130 26682
rect 18130 26630 18142 26682
rect 18142 26630 18172 26682
rect 18196 26630 18206 26682
rect 18206 26630 18252 26682
rect 17956 26628 18012 26630
rect 18036 26628 18092 26630
rect 18116 26628 18172 26630
rect 18196 26628 18252 26630
rect 25956 26682 26012 26684
rect 26036 26682 26092 26684
rect 26116 26682 26172 26684
rect 26196 26682 26252 26684
rect 25956 26630 26002 26682
rect 26002 26630 26012 26682
rect 26036 26630 26066 26682
rect 26066 26630 26078 26682
rect 26078 26630 26092 26682
rect 26116 26630 26130 26682
rect 26130 26630 26142 26682
rect 26142 26630 26172 26682
rect 26196 26630 26206 26682
rect 26206 26630 26252 26682
rect 25956 26628 26012 26630
rect 26036 26628 26092 26630
rect 26116 26628 26172 26630
rect 26196 26628 26252 26630
rect 2616 26138 2672 26140
rect 2696 26138 2752 26140
rect 2776 26138 2832 26140
rect 2856 26138 2912 26140
rect 2616 26086 2662 26138
rect 2662 26086 2672 26138
rect 2696 26086 2726 26138
rect 2726 26086 2738 26138
rect 2738 26086 2752 26138
rect 2776 26086 2790 26138
rect 2790 26086 2802 26138
rect 2802 26086 2832 26138
rect 2856 26086 2866 26138
rect 2866 26086 2912 26138
rect 2616 26084 2672 26086
rect 2696 26084 2752 26086
rect 2776 26084 2832 26086
rect 2856 26084 2912 26086
rect 10616 26138 10672 26140
rect 10696 26138 10752 26140
rect 10776 26138 10832 26140
rect 10856 26138 10912 26140
rect 10616 26086 10662 26138
rect 10662 26086 10672 26138
rect 10696 26086 10726 26138
rect 10726 26086 10738 26138
rect 10738 26086 10752 26138
rect 10776 26086 10790 26138
rect 10790 26086 10802 26138
rect 10802 26086 10832 26138
rect 10856 26086 10866 26138
rect 10866 26086 10912 26138
rect 10616 26084 10672 26086
rect 10696 26084 10752 26086
rect 10776 26084 10832 26086
rect 10856 26084 10912 26086
rect 18616 26138 18672 26140
rect 18696 26138 18752 26140
rect 18776 26138 18832 26140
rect 18856 26138 18912 26140
rect 18616 26086 18662 26138
rect 18662 26086 18672 26138
rect 18696 26086 18726 26138
rect 18726 26086 18738 26138
rect 18738 26086 18752 26138
rect 18776 26086 18790 26138
rect 18790 26086 18802 26138
rect 18802 26086 18832 26138
rect 18856 26086 18866 26138
rect 18866 26086 18912 26138
rect 18616 26084 18672 26086
rect 18696 26084 18752 26086
rect 18776 26084 18832 26086
rect 18856 26084 18912 26086
rect 26616 26138 26672 26140
rect 26696 26138 26752 26140
rect 26776 26138 26832 26140
rect 26856 26138 26912 26140
rect 26616 26086 26662 26138
rect 26662 26086 26672 26138
rect 26696 26086 26726 26138
rect 26726 26086 26738 26138
rect 26738 26086 26752 26138
rect 26776 26086 26790 26138
rect 26790 26086 26802 26138
rect 26802 26086 26832 26138
rect 26856 26086 26866 26138
rect 26866 26086 26912 26138
rect 26616 26084 26672 26086
rect 26696 26084 26752 26086
rect 26776 26084 26832 26086
rect 26856 26084 26912 26086
rect 1956 25594 2012 25596
rect 2036 25594 2092 25596
rect 2116 25594 2172 25596
rect 2196 25594 2252 25596
rect 1956 25542 2002 25594
rect 2002 25542 2012 25594
rect 2036 25542 2066 25594
rect 2066 25542 2078 25594
rect 2078 25542 2092 25594
rect 2116 25542 2130 25594
rect 2130 25542 2142 25594
rect 2142 25542 2172 25594
rect 2196 25542 2206 25594
rect 2206 25542 2252 25594
rect 1956 25540 2012 25542
rect 2036 25540 2092 25542
rect 2116 25540 2172 25542
rect 2196 25540 2252 25542
rect 9956 25594 10012 25596
rect 10036 25594 10092 25596
rect 10116 25594 10172 25596
rect 10196 25594 10252 25596
rect 9956 25542 10002 25594
rect 10002 25542 10012 25594
rect 10036 25542 10066 25594
rect 10066 25542 10078 25594
rect 10078 25542 10092 25594
rect 10116 25542 10130 25594
rect 10130 25542 10142 25594
rect 10142 25542 10172 25594
rect 10196 25542 10206 25594
rect 10206 25542 10252 25594
rect 9956 25540 10012 25542
rect 10036 25540 10092 25542
rect 10116 25540 10172 25542
rect 10196 25540 10252 25542
rect 17956 25594 18012 25596
rect 18036 25594 18092 25596
rect 18116 25594 18172 25596
rect 18196 25594 18252 25596
rect 17956 25542 18002 25594
rect 18002 25542 18012 25594
rect 18036 25542 18066 25594
rect 18066 25542 18078 25594
rect 18078 25542 18092 25594
rect 18116 25542 18130 25594
rect 18130 25542 18142 25594
rect 18142 25542 18172 25594
rect 18196 25542 18206 25594
rect 18206 25542 18252 25594
rect 17956 25540 18012 25542
rect 18036 25540 18092 25542
rect 18116 25540 18172 25542
rect 18196 25540 18252 25542
rect 25956 25594 26012 25596
rect 26036 25594 26092 25596
rect 26116 25594 26172 25596
rect 26196 25594 26252 25596
rect 25956 25542 26002 25594
rect 26002 25542 26012 25594
rect 26036 25542 26066 25594
rect 26066 25542 26078 25594
rect 26078 25542 26092 25594
rect 26116 25542 26130 25594
rect 26130 25542 26142 25594
rect 26142 25542 26172 25594
rect 26196 25542 26206 25594
rect 26206 25542 26252 25594
rect 25956 25540 26012 25542
rect 26036 25540 26092 25542
rect 26116 25540 26172 25542
rect 26196 25540 26252 25542
rect 2616 25050 2672 25052
rect 2696 25050 2752 25052
rect 2776 25050 2832 25052
rect 2856 25050 2912 25052
rect 2616 24998 2662 25050
rect 2662 24998 2672 25050
rect 2696 24998 2726 25050
rect 2726 24998 2738 25050
rect 2738 24998 2752 25050
rect 2776 24998 2790 25050
rect 2790 24998 2802 25050
rect 2802 24998 2832 25050
rect 2856 24998 2866 25050
rect 2866 24998 2912 25050
rect 2616 24996 2672 24998
rect 2696 24996 2752 24998
rect 2776 24996 2832 24998
rect 2856 24996 2912 24998
rect 10616 25050 10672 25052
rect 10696 25050 10752 25052
rect 10776 25050 10832 25052
rect 10856 25050 10912 25052
rect 10616 24998 10662 25050
rect 10662 24998 10672 25050
rect 10696 24998 10726 25050
rect 10726 24998 10738 25050
rect 10738 24998 10752 25050
rect 10776 24998 10790 25050
rect 10790 24998 10802 25050
rect 10802 24998 10832 25050
rect 10856 24998 10866 25050
rect 10866 24998 10912 25050
rect 10616 24996 10672 24998
rect 10696 24996 10752 24998
rect 10776 24996 10832 24998
rect 10856 24996 10912 24998
rect 18616 25050 18672 25052
rect 18696 25050 18752 25052
rect 18776 25050 18832 25052
rect 18856 25050 18912 25052
rect 18616 24998 18662 25050
rect 18662 24998 18672 25050
rect 18696 24998 18726 25050
rect 18726 24998 18738 25050
rect 18738 24998 18752 25050
rect 18776 24998 18790 25050
rect 18790 24998 18802 25050
rect 18802 24998 18832 25050
rect 18856 24998 18866 25050
rect 18866 24998 18912 25050
rect 18616 24996 18672 24998
rect 18696 24996 18752 24998
rect 18776 24996 18832 24998
rect 18856 24996 18912 24998
rect 26616 25050 26672 25052
rect 26696 25050 26752 25052
rect 26776 25050 26832 25052
rect 26856 25050 26912 25052
rect 26616 24998 26662 25050
rect 26662 24998 26672 25050
rect 26696 24998 26726 25050
rect 26726 24998 26738 25050
rect 26738 24998 26752 25050
rect 26776 24998 26790 25050
rect 26790 24998 26802 25050
rect 26802 24998 26832 25050
rect 26856 24998 26866 25050
rect 26866 24998 26912 25050
rect 26616 24996 26672 24998
rect 26696 24996 26752 24998
rect 26776 24996 26832 24998
rect 26856 24996 26912 24998
rect 1956 24506 2012 24508
rect 2036 24506 2092 24508
rect 2116 24506 2172 24508
rect 2196 24506 2252 24508
rect 1956 24454 2002 24506
rect 2002 24454 2012 24506
rect 2036 24454 2066 24506
rect 2066 24454 2078 24506
rect 2078 24454 2092 24506
rect 2116 24454 2130 24506
rect 2130 24454 2142 24506
rect 2142 24454 2172 24506
rect 2196 24454 2206 24506
rect 2206 24454 2252 24506
rect 1956 24452 2012 24454
rect 2036 24452 2092 24454
rect 2116 24452 2172 24454
rect 2196 24452 2252 24454
rect 9956 24506 10012 24508
rect 10036 24506 10092 24508
rect 10116 24506 10172 24508
rect 10196 24506 10252 24508
rect 9956 24454 10002 24506
rect 10002 24454 10012 24506
rect 10036 24454 10066 24506
rect 10066 24454 10078 24506
rect 10078 24454 10092 24506
rect 10116 24454 10130 24506
rect 10130 24454 10142 24506
rect 10142 24454 10172 24506
rect 10196 24454 10206 24506
rect 10206 24454 10252 24506
rect 9956 24452 10012 24454
rect 10036 24452 10092 24454
rect 10116 24452 10172 24454
rect 10196 24452 10252 24454
rect 17956 24506 18012 24508
rect 18036 24506 18092 24508
rect 18116 24506 18172 24508
rect 18196 24506 18252 24508
rect 17956 24454 18002 24506
rect 18002 24454 18012 24506
rect 18036 24454 18066 24506
rect 18066 24454 18078 24506
rect 18078 24454 18092 24506
rect 18116 24454 18130 24506
rect 18130 24454 18142 24506
rect 18142 24454 18172 24506
rect 18196 24454 18206 24506
rect 18206 24454 18252 24506
rect 17956 24452 18012 24454
rect 18036 24452 18092 24454
rect 18116 24452 18172 24454
rect 18196 24452 18252 24454
rect 25956 24506 26012 24508
rect 26036 24506 26092 24508
rect 26116 24506 26172 24508
rect 26196 24506 26252 24508
rect 25956 24454 26002 24506
rect 26002 24454 26012 24506
rect 26036 24454 26066 24506
rect 26066 24454 26078 24506
rect 26078 24454 26092 24506
rect 26116 24454 26130 24506
rect 26130 24454 26142 24506
rect 26142 24454 26172 24506
rect 26196 24454 26206 24506
rect 26206 24454 26252 24506
rect 25956 24452 26012 24454
rect 26036 24452 26092 24454
rect 26116 24452 26172 24454
rect 26196 24452 26252 24454
rect 2616 23962 2672 23964
rect 2696 23962 2752 23964
rect 2776 23962 2832 23964
rect 2856 23962 2912 23964
rect 2616 23910 2662 23962
rect 2662 23910 2672 23962
rect 2696 23910 2726 23962
rect 2726 23910 2738 23962
rect 2738 23910 2752 23962
rect 2776 23910 2790 23962
rect 2790 23910 2802 23962
rect 2802 23910 2832 23962
rect 2856 23910 2866 23962
rect 2866 23910 2912 23962
rect 2616 23908 2672 23910
rect 2696 23908 2752 23910
rect 2776 23908 2832 23910
rect 2856 23908 2912 23910
rect 10616 23962 10672 23964
rect 10696 23962 10752 23964
rect 10776 23962 10832 23964
rect 10856 23962 10912 23964
rect 10616 23910 10662 23962
rect 10662 23910 10672 23962
rect 10696 23910 10726 23962
rect 10726 23910 10738 23962
rect 10738 23910 10752 23962
rect 10776 23910 10790 23962
rect 10790 23910 10802 23962
rect 10802 23910 10832 23962
rect 10856 23910 10866 23962
rect 10866 23910 10912 23962
rect 10616 23908 10672 23910
rect 10696 23908 10752 23910
rect 10776 23908 10832 23910
rect 10856 23908 10912 23910
rect 18616 23962 18672 23964
rect 18696 23962 18752 23964
rect 18776 23962 18832 23964
rect 18856 23962 18912 23964
rect 18616 23910 18662 23962
rect 18662 23910 18672 23962
rect 18696 23910 18726 23962
rect 18726 23910 18738 23962
rect 18738 23910 18752 23962
rect 18776 23910 18790 23962
rect 18790 23910 18802 23962
rect 18802 23910 18832 23962
rect 18856 23910 18866 23962
rect 18866 23910 18912 23962
rect 18616 23908 18672 23910
rect 18696 23908 18752 23910
rect 18776 23908 18832 23910
rect 18856 23908 18912 23910
rect 26616 23962 26672 23964
rect 26696 23962 26752 23964
rect 26776 23962 26832 23964
rect 26856 23962 26912 23964
rect 26616 23910 26662 23962
rect 26662 23910 26672 23962
rect 26696 23910 26726 23962
rect 26726 23910 26738 23962
rect 26738 23910 26752 23962
rect 26776 23910 26790 23962
rect 26790 23910 26802 23962
rect 26802 23910 26832 23962
rect 26856 23910 26866 23962
rect 26866 23910 26912 23962
rect 26616 23908 26672 23910
rect 26696 23908 26752 23910
rect 26776 23908 26832 23910
rect 26856 23908 26912 23910
rect 1956 23418 2012 23420
rect 2036 23418 2092 23420
rect 2116 23418 2172 23420
rect 2196 23418 2252 23420
rect 1956 23366 2002 23418
rect 2002 23366 2012 23418
rect 2036 23366 2066 23418
rect 2066 23366 2078 23418
rect 2078 23366 2092 23418
rect 2116 23366 2130 23418
rect 2130 23366 2142 23418
rect 2142 23366 2172 23418
rect 2196 23366 2206 23418
rect 2206 23366 2252 23418
rect 1956 23364 2012 23366
rect 2036 23364 2092 23366
rect 2116 23364 2172 23366
rect 2196 23364 2252 23366
rect 9956 23418 10012 23420
rect 10036 23418 10092 23420
rect 10116 23418 10172 23420
rect 10196 23418 10252 23420
rect 9956 23366 10002 23418
rect 10002 23366 10012 23418
rect 10036 23366 10066 23418
rect 10066 23366 10078 23418
rect 10078 23366 10092 23418
rect 10116 23366 10130 23418
rect 10130 23366 10142 23418
rect 10142 23366 10172 23418
rect 10196 23366 10206 23418
rect 10206 23366 10252 23418
rect 9956 23364 10012 23366
rect 10036 23364 10092 23366
rect 10116 23364 10172 23366
rect 10196 23364 10252 23366
rect 17956 23418 18012 23420
rect 18036 23418 18092 23420
rect 18116 23418 18172 23420
rect 18196 23418 18252 23420
rect 17956 23366 18002 23418
rect 18002 23366 18012 23418
rect 18036 23366 18066 23418
rect 18066 23366 18078 23418
rect 18078 23366 18092 23418
rect 18116 23366 18130 23418
rect 18130 23366 18142 23418
rect 18142 23366 18172 23418
rect 18196 23366 18206 23418
rect 18206 23366 18252 23418
rect 17956 23364 18012 23366
rect 18036 23364 18092 23366
rect 18116 23364 18172 23366
rect 18196 23364 18252 23366
rect 25956 23418 26012 23420
rect 26036 23418 26092 23420
rect 26116 23418 26172 23420
rect 26196 23418 26252 23420
rect 25956 23366 26002 23418
rect 26002 23366 26012 23418
rect 26036 23366 26066 23418
rect 26066 23366 26078 23418
rect 26078 23366 26092 23418
rect 26116 23366 26130 23418
rect 26130 23366 26142 23418
rect 26142 23366 26172 23418
rect 26196 23366 26206 23418
rect 26206 23366 26252 23418
rect 25956 23364 26012 23366
rect 26036 23364 26092 23366
rect 26116 23364 26172 23366
rect 26196 23364 26252 23366
rect 2616 22874 2672 22876
rect 2696 22874 2752 22876
rect 2776 22874 2832 22876
rect 2856 22874 2912 22876
rect 2616 22822 2662 22874
rect 2662 22822 2672 22874
rect 2696 22822 2726 22874
rect 2726 22822 2738 22874
rect 2738 22822 2752 22874
rect 2776 22822 2790 22874
rect 2790 22822 2802 22874
rect 2802 22822 2832 22874
rect 2856 22822 2866 22874
rect 2866 22822 2912 22874
rect 2616 22820 2672 22822
rect 2696 22820 2752 22822
rect 2776 22820 2832 22822
rect 2856 22820 2912 22822
rect 10616 22874 10672 22876
rect 10696 22874 10752 22876
rect 10776 22874 10832 22876
rect 10856 22874 10912 22876
rect 10616 22822 10662 22874
rect 10662 22822 10672 22874
rect 10696 22822 10726 22874
rect 10726 22822 10738 22874
rect 10738 22822 10752 22874
rect 10776 22822 10790 22874
rect 10790 22822 10802 22874
rect 10802 22822 10832 22874
rect 10856 22822 10866 22874
rect 10866 22822 10912 22874
rect 10616 22820 10672 22822
rect 10696 22820 10752 22822
rect 10776 22820 10832 22822
rect 10856 22820 10912 22822
rect 18616 22874 18672 22876
rect 18696 22874 18752 22876
rect 18776 22874 18832 22876
rect 18856 22874 18912 22876
rect 18616 22822 18662 22874
rect 18662 22822 18672 22874
rect 18696 22822 18726 22874
rect 18726 22822 18738 22874
rect 18738 22822 18752 22874
rect 18776 22822 18790 22874
rect 18790 22822 18802 22874
rect 18802 22822 18832 22874
rect 18856 22822 18866 22874
rect 18866 22822 18912 22874
rect 18616 22820 18672 22822
rect 18696 22820 18752 22822
rect 18776 22820 18832 22822
rect 18856 22820 18912 22822
rect 26616 22874 26672 22876
rect 26696 22874 26752 22876
rect 26776 22874 26832 22876
rect 26856 22874 26912 22876
rect 26616 22822 26662 22874
rect 26662 22822 26672 22874
rect 26696 22822 26726 22874
rect 26726 22822 26738 22874
rect 26738 22822 26752 22874
rect 26776 22822 26790 22874
rect 26790 22822 26802 22874
rect 26802 22822 26832 22874
rect 26856 22822 26866 22874
rect 26866 22822 26912 22874
rect 26616 22820 26672 22822
rect 26696 22820 26752 22822
rect 26776 22820 26832 22822
rect 26856 22820 26912 22822
rect 846 22480 902 22536
rect 1956 22330 2012 22332
rect 2036 22330 2092 22332
rect 2116 22330 2172 22332
rect 2196 22330 2252 22332
rect 1956 22278 2002 22330
rect 2002 22278 2012 22330
rect 2036 22278 2066 22330
rect 2066 22278 2078 22330
rect 2078 22278 2092 22330
rect 2116 22278 2130 22330
rect 2130 22278 2142 22330
rect 2142 22278 2172 22330
rect 2196 22278 2206 22330
rect 2206 22278 2252 22330
rect 1956 22276 2012 22278
rect 2036 22276 2092 22278
rect 2116 22276 2172 22278
rect 2196 22276 2252 22278
rect 9956 22330 10012 22332
rect 10036 22330 10092 22332
rect 10116 22330 10172 22332
rect 10196 22330 10252 22332
rect 9956 22278 10002 22330
rect 10002 22278 10012 22330
rect 10036 22278 10066 22330
rect 10066 22278 10078 22330
rect 10078 22278 10092 22330
rect 10116 22278 10130 22330
rect 10130 22278 10142 22330
rect 10142 22278 10172 22330
rect 10196 22278 10206 22330
rect 10206 22278 10252 22330
rect 9956 22276 10012 22278
rect 10036 22276 10092 22278
rect 10116 22276 10172 22278
rect 10196 22276 10252 22278
rect 17956 22330 18012 22332
rect 18036 22330 18092 22332
rect 18116 22330 18172 22332
rect 18196 22330 18252 22332
rect 17956 22278 18002 22330
rect 18002 22278 18012 22330
rect 18036 22278 18066 22330
rect 18066 22278 18078 22330
rect 18078 22278 18092 22330
rect 18116 22278 18130 22330
rect 18130 22278 18142 22330
rect 18142 22278 18172 22330
rect 18196 22278 18206 22330
rect 18206 22278 18252 22330
rect 17956 22276 18012 22278
rect 18036 22276 18092 22278
rect 18116 22276 18172 22278
rect 18196 22276 18252 22278
rect 25956 22330 26012 22332
rect 26036 22330 26092 22332
rect 26116 22330 26172 22332
rect 26196 22330 26252 22332
rect 25956 22278 26002 22330
rect 26002 22278 26012 22330
rect 26036 22278 26066 22330
rect 26066 22278 26078 22330
rect 26078 22278 26092 22330
rect 26116 22278 26130 22330
rect 26130 22278 26142 22330
rect 26142 22278 26172 22330
rect 26196 22278 26206 22330
rect 26206 22278 26252 22330
rect 25956 22276 26012 22278
rect 26036 22276 26092 22278
rect 26116 22276 26172 22278
rect 26196 22276 26252 22278
rect 2616 21786 2672 21788
rect 2696 21786 2752 21788
rect 2776 21786 2832 21788
rect 2856 21786 2912 21788
rect 2616 21734 2662 21786
rect 2662 21734 2672 21786
rect 2696 21734 2726 21786
rect 2726 21734 2738 21786
rect 2738 21734 2752 21786
rect 2776 21734 2790 21786
rect 2790 21734 2802 21786
rect 2802 21734 2832 21786
rect 2856 21734 2866 21786
rect 2866 21734 2912 21786
rect 2616 21732 2672 21734
rect 2696 21732 2752 21734
rect 2776 21732 2832 21734
rect 2856 21732 2912 21734
rect 10616 21786 10672 21788
rect 10696 21786 10752 21788
rect 10776 21786 10832 21788
rect 10856 21786 10912 21788
rect 10616 21734 10662 21786
rect 10662 21734 10672 21786
rect 10696 21734 10726 21786
rect 10726 21734 10738 21786
rect 10738 21734 10752 21786
rect 10776 21734 10790 21786
rect 10790 21734 10802 21786
rect 10802 21734 10832 21786
rect 10856 21734 10866 21786
rect 10866 21734 10912 21786
rect 10616 21732 10672 21734
rect 10696 21732 10752 21734
rect 10776 21732 10832 21734
rect 10856 21732 10912 21734
rect 18616 21786 18672 21788
rect 18696 21786 18752 21788
rect 18776 21786 18832 21788
rect 18856 21786 18912 21788
rect 18616 21734 18662 21786
rect 18662 21734 18672 21786
rect 18696 21734 18726 21786
rect 18726 21734 18738 21786
rect 18738 21734 18752 21786
rect 18776 21734 18790 21786
rect 18790 21734 18802 21786
rect 18802 21734 18832 21786
rect 18856 21734 18866 21786
rect 18866 21734 18912 21786
rect 18616 21732 18672 21734
rect 18696 21732 18752 21734
rect 18776 21732 18832 21734
rect 18856 21732 18912 21734
rect 26616 21786 26672 21788
rect 26696 21786 26752 21788
rect 26776 21786 26832 21788
rect 26856 21786 26912 21788
rect 26616 21734 26662 21786
rect 26662 21734 26672 21786
rect 26696 21734 26726 21786
rect 26726 21734 26738 21786
rect 26738 21734 26752 21786
rect 26776 21734 26790 21786
rect 26790 21734 26802 21786
rect 26802 21734 26832 21786
rect 26856 21734 26866 21786
rect 26866 21734 26912 21786
rect 26616 21732 26672 21734
rect 26696 21732 26752 21734
rect 26776 21732 26832 21734
rect 26856 21732 26912 21734
rect 1956 21242 2012 21244
rect 2036 21242 2092 21244
rect 2116 21242 2172 21244
rect 2196 21242 2252 21244
rect 1956 21190 2002 21242
rect 2002 21190 2012 21242
rect 2036 21190 2066 21242
rect 2066 21190 2078 21242
rect 2078 21190 2092 21242
rect 2116 21190 2130 21242
rect 2130 21190 2142 21242
rect 2142 21190 2172 21242
rect 2196 21190 2206 21242
rect 2206 21190 2252 21242
rect 1956 21188 2012 21190
rect 2036 21188 2092 21190
rect 2116 21188 2172 21190
rect 2196 21188 2252 21190
rect 9956 21242 10012 21244
rect 10036 21242 10092 21244
rect 10116 21242 10172 21244
rect 10196 21242 10252 21244
rect 9956 21190 10002 21242
rect 10002 21190 10012 21242
rect 10036 21190 10066 21242
rect 10066 21190 10078 21242
rect 10078 21190 10092 21242
rect 10116 21190 10130 21242
rect 10130 21190 10142 21242
rect 10142 21190 10172 21242
rect 10196 21190 10206 21242
rect 10206 21190 10252 21242
rect 9956 21188 10012 21190
rect 10036 21188 10092 21190
rect 10116 21188 10172 21190
rect 10196 21188 10252 21190
rect 17956 21242 18012 21244
rect 18036 21242 18092 21244
rect 18116 21242 18172 21244
rect 18196 21242 18252 21244
rect 17956 21190 18002 21242
rect 18002 21190 18012 21242
rect 18036 21190 18066 21242
rect 18066 21190 18078 21242
rect 18078 21190 18092 21242
rect 18116 21190 18130 21242
rect 18130 21190 18142 21242
rect 18142 21190 18172 21242
rect 18196 21190 18206 21242
rect 18206 21190 18252 21242
rect 17956 21188 18012 21190
rect 18036 21188 18092 21190
rect 18116 21188 18172 21190
rect 18196 21188 18252 21190
rect 25956 21242 26012 21244
rect 26036 21242 26092 21244
rect 26116 21242 26172 21244
rect 26196 21242 26252 21244
rect 25956 21190 26002 21242
rect 26002 21190 26012 21242
rect 26036 21190 26066 21242
rect 26066 21190 26078 21242
rect 26078 21190 26092 21242
rect 26116 21190 26130 21242
rect 26130 21190 26142 21242
rect 26142 21190 26172 21242
rect 26196 21190 26206 21242
rect 26206 21190 26252 21242
rect 25956 21188 26012 21190
rect 26036 21188 26092 21190
rect 26116 21188 26172 21190
rect 26196 21188 26252 21190
rect 2616 20698 2672 20700
rect 2696 20698 2752 20700
rect 2776 20698 2832 20700
rect 2856 20698 2912 20700
rect 2616 20646 2662 20698
rect 2662 20646 2672 20698
rect 2696 20646 2726 20698
rect 2726 20646 2738 20698
rect 2738 20646 2752 20698
rect 2776 20646 2790 20698
rect 2790 20646 2802 20698
rect 2802 20646 2832 20698
rect 2856 20646 2866 20698
rect 2866 20646 2912 20698
rect 2616 20644 2672 20646
rect 2696 20644 2752 20646
rect 2776 20644 2832 20646
rect 2856 20644 2912 20646
rect 10616 20698 10672 20700
rect 10696 20698 10752 20700
rect 10776 20698 10832 20700
rect 10856 20698 10912 20700
rect 10616 20646 10662 20698
rect 10662 20646 10672 20698
rect 10696 20646 10726 20698
rect 10726 20646 10738 20698
rect 10738 20646 10752 20698
rect 10776 20646 10790 20698
rect 10790 20646 10802 20698
rect 10802 20646 10832 20698
rect 10856 20646 10866 20698
rect 10866 20646 10912 20698
rect 10616 20644 10672 20646
rect 10696 20644 10752 20646
rect 10776 20644 10832 20646
rect 10856 20644 10912 20646
rect 18616 20698 18672 20700
rect 18696 20698 18752 20700
rect 18776 20698 18832 20700
rect 18856 20698 18912 20700
rect 18616 20646 18662 20698
rect 18662 20646 18672 20698
rect 18696 20646 18726 20698
rect 18726 20646 18738 20698
rect 18738 20646 18752 20698
rect 18776 20646 18790 20698
rect 18790 20646 18802 20698
rect 18802 20646 18832 20698
rect 18856 20646 18866 20698
rect 18866 20646 18912 20698
rect 18616 20644 18672 20646
rect 18696 20644 18752 20646
rect 18776 20644 18832 20646
rect 18856 20644 18912 20646
rect 26616 20698 26672 20700
rect 26696 20698 26752 20700
rect 26776 20698 26832 20700
rect 26856 20698 26912 20700
rect 26616 20646 26662 20698
rect 26662 20646 26672 20698
rect 26696 20646 26726 20698
rect 26726 20646 26738 20698
rect 26738 20646 26752 20698
rect 26776 20646 26790 20698
rect 26790 20646 26802 20698
rect 26802 20646 26832 20698
rect 26856 20646 26866 20698
rect 26866 20646 26912 20698
rect 26616 20644 26672 20646
rect 26696 20644 26752 20646
rect 26776 20644 26832 20646
rect 26856 20644 26912 20646
rect 1956 20154 2012 20156
rect 2036 20154 2092 20156
rect 2116 20154 2172 20156
rect 2196 20154 2252 20156
rect 1956 20102 2002 20154
rect 2002 20102 2012 20154
rect 2036 20102 2066 20154
rect 2066 20102 2078 20154
rect 2078 20102 2092 20154
rect 2116 20102 2130 20154
rect 2130 20102 2142 20154
rect 2142 20102 2172 20154
rect 2196 20102 2206 20154
rect 2206 20102 2252 20154
rect 1956 20100 2012 20102
rect 2036 20100 2092 20102
rect 2116 20100 2172 20102
rect 2196 20100 2252 20102
rect 9956 20154 10012 20156
rect 10036 20154 10092 20156
rect 10116 20154 10172 20156
rect 10196 20154 10252 20156
rect 9956 20102 10002 20154
rect 10002 20102 10012 20154
rect 10036 20102 10066 20154
rect 10066 20102 10078 20154
rect 10078 20102 10092 20154
rect 10116 20102 10130 20154
rect 10130 20102 10142 20154
rect 10142 20102 10172 20154
rect 10196 20102 10206 20154
rect 10206 20102 10252 20154
rect 9956 20100 10012 20102
rect 10036 20100 10092 20102
rect 10116 20100 10172 20102
rect 10196 20100 10252 20102
rect 17956 20154 18012 20156
rect 18036 20154 18092 20156
rect 18116 20154 18172 20156
rect 18196 20154 18252 20156
rect 17956 20102 18002 20154
rect 18002 20102 18012 20154
rect 18036 20102 18066 20154
rect 18066 20102 18078 20154
rect 18078 20102 18092 20154
rect 18116 20102 18130 20154
rect 18130 20102 18142 20154
rect 18142 20102 18172 20154
rect 18196 20102 18206 20154
rect 18206 20102 18252 20154
rect 17956 20100 18012 20102
rect 18036 20100 18092 20102
rect 18116 20100 18172 20102
rect 18196 20100 18252 20102
rect 25956 20154 26012 20156
rect 26036 20154 26092 20156
rect 26116 20154 26172 20156
rect 26196 20154 26252 20156
rect 25956 20102 26002 20154
rect 26002 20102 26012 20154
rect 26036 20102 26066 20154
rect 26066 20102 26078 20154
rect 26078 20102 26092 20154
rect 26116 20102 26130 20154
rect 26130 20102 26142 20154
rect 26142 20102 26172 20154
rect 26196 20102 26206 20154
rect 26206 20102 26252 20154
rect 25956 20100 26012 20102
rect 26036 20100 26092 20102
rect 26116 20100 26172 20102
rect 26196 20100 26252 20102
rect 2616 19610 2672 19612
rect 2696 19610 2752 19612
rect 2776 19610 2832 19612
rect 2856 19610 2912 19612
rect 2616 19558 2662 19610
rect 2662 19558 2672 19610
rect 2696 19558 2726 19610
rect 2726 19558 2738 19610
rect 2738 19558 2752 19610
rect 2776 19558 2790 19610
rect 2790 19558 2802 19610
rect 2802 19558 2832 19610
rect 2856 19558 2866 19610
rect 2866 19558 2912 19610
rect 2616 19556 2672 19558
rect 2696 19556 2752 19558
rect 2776 19556 2832 19558
rect 2856 19556 2912 19558
rect 10616 19610 10672 19612
rect 10696 19610 10752 19612
rect 10776 19610 10832 19612
rect 10856 19610 10912 19612
rect 10616 19558 10662 19610
rect 10662 19558 10672 19610
rect 10696 19558 10726 19610
rect 10726 19558 10738 19610
rect 10738 19558 10752 19610
rect 10776 19558 10790 19610
rect 10790 19558 10802 19610
rect 10802 19558 10832 19610
rect 10856 19558 10866 19610
rect 10866 19558 10912 19610
rect 10616 19556 10672 19558
rect 10696 19556 10752 19558
rect 10776 19556 10832 19558
rect 10856 19556 10912 19558
rect 18616 19610 18672 19612
rect 18696 19610 18752 19612
rect 18776 19610 18832 19612
rect 18856 19610 18912 19612
rect 18616 19558 18662 19610
rect 18662 19558 18672 19610
rect 18696 19558 18726 19610
rect 18726 19558 18738 19610
rect 18738 19558 18752 19610
rect 18776 19558 18790 19610
rect 18790 19558 18802 19610
rect 18802 19558 18832 19610
rect 18856 19558 18866 19610
rect 18866 19558 18912 19610
rect 18616 19556 18672 19558
rect 18696 19556 18752 19558
rect 18776 19556 18832 19558
rect 18856 19556 18912 19558
rect 26616 19610 26672 19612
rect 26696 19610 26752 19612
rect 26776 19610 26832 19612
rect 26856 19610 26912 19612
rect 26616 19558 26662 19610
rect 26662 19558 26672 19610
rect 26696 19558 26726 19610
rect 26726 19558 26738 19610
rect 26738 19558 26752 19610
rect 26776 19558 26790 19610
rect 26790 19558 26802 19610
rect 26802 19558 26832 19610
rect 26856 19558 26866 19610
rect 26866 19558 26912 19610
rect 26616 19556 26672 19558
rect 26696 19556 26752 19558
rect 26776 19556 26832 19558
rect 26856 19556 26912 19558
rect 1956 19066 2012 19068
rect 2036 19066 2092 19068
rect 2116 19066 2172 19068
rect 2196 19066 2252 19068
rect 1956 19014 2002 19066
rect 2002 19014 2012 19066
rect 2036 19014 2066 19066
rect 2066 19014 2078 19066
rect 2078 19014 2092 19066
rect 2116 19014 2130 19066
rect 2130 19014 2142 19066
rect 2142 19014 2172 19066
rect 2196 19014 2206 19066
rect 2206 19014 2252 19066
rect 1956 19012 2012 19014
rect 2036 19012 2092 19014
rect 2116 19012 2172 19014
rect 2196 19012 2252 19014
rect 9956 19066 10012 19068
rect 10036 19066 10092 19068
rect 10116 19066 10172 19068
rect 10196 19066 10252 19068
rect 9956 19014 10002 19066
rect 10002 19014 10012 19066
rect 10036 19014 10066 19066
rect 10066 19014 10078 19066
rect 10078 19014 10092 19066
rect 10116 19014 10130 19066
rect 10130 19014 10142 19066
rect 10142 19014 10172 19066
rect 10196 19014 10206 19066
rect 10206 19014 10252 19066
rect 9956 19012 10012 19014
rect 10036 19012 10092 19014
rect 10116 19012 10172 19014
rect 10196 19012 10252 19014
rect 17956 19066 18012 19068
rect 18036 19066 18092 19068
rect 18116 19066 18172 19068
rect 18196 19066 18252 19068
rect 17956 19014 18002 19066
rect 18002 19014 18012 19066
rect 18036 19014 18066 19066
rect 18066 19014 18078 19066
rect 18078 19014 18092 19066
rect 18116 19014 18130 19066
rect 18130 19014 18142 19066
rect 18142 19014 18172 19066
rect 18196 19014 18206 19066
rect 18206 19014 18252 19066
rect 17956 19012 18012 19014
rect 18036 19012 18092 19014
rect 18116 19012 18172 19014
rect 18196 19012 18252 19014
rect 25956 19066 26012 19068
rect 26036 19066 26092 19068
rect 26116 19066 26172 19068
rect 26196 19066 26252 19068
rect 25956 19014 26002 19066
rect 26002 19014 26012 19066
rect 26036 19014 26066 19066
rect 26066 19014 26078 19066
rect 26078 19014 26092 19066
rect 26116 19014 26130 19066
rect 26130 19014 26142 19066
rect 26142 19014 26172 19066
rect 26196 19014 26206 19066
rect 26206 19014 26252 19066
rect 25956 19012 26012 19014
rect 26036 19012 26092 19014
rect 26116 19012 26172 19014
rect 26196 19012 26252 19014
rect 2616 18522 2672 18524
rect 2696 18522 2752 18524
rect 2776 18522 2832 18524
rect 2856 18522 2912 18524
rect 2616 18470 2662 18522
rect 2662 18470 2672 18522
rect 2696 18470 2726 18522
rect 2726 18470 2738 18522
rect 2738 18470 2752 18522
rect 2776 18470 2790 18522
rect 2790 18470 2802 18522
rect 2802 18470 2832 18522
rect 2856 18470 2866 18522
rect 2866 18470 2912 18522
rect 2616 18468 2672 18470
rect 2696 18468 2752 18470
rect 2776 18468 2832 18470
rect 2856 18468 2912 18470
rect 10616 18522 10672 18524
rect 10696 18522 10752 18524
rect 10776 18522 10832 18524
rect 10856 18522 10912 18524
rect 10616 18470 10662 18522
rect 10662 18470 10672 18522
rect 10696 18470 10726 18522
rect 10726 18470 10738 18522
rect 10738 18470 10752 18522
rect 10776 18470 10790 18522
rect 10790 18470 10802 18522
rect 10802 18470 10832 18522
rect 10856 18470 10866 18522
rect 10866 18470 10912 18522
rect 10616 18468 10672 18470
rect 10696 18468 10752 18470
rect 10776 18468 10832 18470
rect 10856 18468 10912 18470
rect 18616 18522 18672 18524
rect 18696 18522 18752 18524
rect 18776 18522 18832 18524
rect 18856 18522 18912 18524
rect 18616 18470 18662 18522
rect 18662 18470 18672 18522
rect 18696 18470 18726 18522
rect 18726 18470 18738 18522
rect 18738 18470 18752 18522
rect 18776 18470 18790 18522
rect 18790 18470 18802 18522
rect 18802 18470 18832 18522
rect 18856 18470 18866 18522
rect 18866 18470 18912 18522
rect 18616 18468 18672 18470
rect 18696 18468 18752 18470
rect 18776 18468 18832 18470
rect 18856 18468 18912 18470
rect 26616 18522 26672 18524
rect 26696 18522 26752 18524
rect 26776 18522 26832 18524
rect 26856 18522 26912 18524
rect 26616 18470 26662 18522
rect 26662 18470 26672 18522
rect 26696 18470 26726 18522
rect 26726 18470 26738 18522
rect 26738 18470 26752 18522
rect 26776 18470 26790 18522
rect 26790 18470 26802 18522
rect 26802 18470 26832 18522
rect 26856 18470 26866 18522
rect 26866 18470 26912 18522
rect 26616 18468 26672 18470
rect 26696 18468 26752 18470
rect 26776 18468 26832 18470
rect 26856 18468 26912 18470
rect 1956 17978 2012 17980
rect 2036 17978 2092 17980
rect 2116 17978 2172 17980
rect 2196 17978 2252 17980
rect 1956 17926 2002 17978
rect 2002 17926 2012 17978
rect 2036 17926 2066 17978
rect 2066 17926 2078 17978
rect 2078 17926 2092 17978
rect 2116 17926 2130 17978
rect 2130 17926 2142 17978
rect 2142 17926 2172 17978
rect 2196 17926 2206 17978
rect 2206 17926 2252 17978
rect 1956 17924 2012 17926
rect 2036 17924 2092 17926
rect 2116 17924 2172 17926
rect 2196 17924 2252 17926
rect 9956 17978 10012 17980
rect 10036 17978 10092 17980
rect 10116 17978 10172 17980
rect 10196 17978 10252 17980
rect 9956 17926 10002 17978
rect 10002 17926 10012 17978
rect 10036 17926 10066 17978
rect 10066 17926 10078 17978
rect 10078 17926 10092 17978
rect 10116 17926 10130 17978
rect 10130 17926 10142 17978
rect 10142 17926 10172 17978
rect 10196 17926 10206 17978
rect 10206 17926 10252 17978
rect 9956 17924 10012 17926
rect 10036 17924 10092 17926
rect 10116 17924 10172 17926
rect 10196 17924 10252 17926
rect 17956 17978 18012 17980
rect 18036 17978 18092 17980
rect 18116 17978 18172 17980
rect 18196 17978 18252 17980
rect 17956 17926 18002 17978
rect 18002 17926 18012 17978
rect 18036 17926 18066 17978
rect 18066 17926 18078 17978
rect 18078 17926 18092 17978
rect 18116 17926 18130 17978
rect 18130 17926 18142 17978
rect 18142 17926 18172 17978
rect 18196 17926 18206 17978
rect 18206 17926 18252 17978
rect 17956 17924 18012 17926
rect 18036 17924 18092 17926
rect 18116 17924 18172 17926
rect 18196 17924 18252 17926
rect 25956 17978 26012 17980
rect 26036 17978 26092 17980
rect 26116 17978 26172 17980
rect 26196 17978 26252 17980
rect 25956 17926 26002 17978
rect 26002 17926 26012 17978
rect 26036 17926 26066 17978
rect 26066 17926 26078 17978
rect 26078 17926 26092 17978
rect 26116 17926 26130 17978
rect 26130 17926 26142 17978
rect 26142 17926 26172 17978
rect 26196 17926 26206 17978
rect 26206 17926 26252 17978
rect 25956 17924 26012 17926
rect 26036 17924 26092 17926
rect 26116 17924 26172 17926
rect 26196 17924 26252 17926
rect 2616 17434 2672 17436
rect 2696 17434 2752 17436
rect 2776 17434 2832 17436
rect 2856 17434 2912 17436
rect 2616 17382 2662 17434
rect 2662 17382 2672 17434
rect 2696 17382 2726 17434
rect 2726 17382 2738 17434
rect 2738 17382 2752 17434
rect 2776 17382 2790 17434
rect 2790 17382 2802 17434
rect 2802 17382 2832 17434
rect 2856 17382 2866 17434
rect 2866 17382 2912 17434
rect 2616 17380 2672 17382
rect 2696 17380 2752 17382
rect 2776 17380 2832 17382
rect 2856 17380 2912 17382
rect 10616 17434 10672 17436
rect 10696 17434 10752 17436
rect 10776 17434 10832 17436
rect 10856 17434 10912 17436
rect 10616 17382 10662 17434
rect 10662 17382 10672 17434
rect 10696 17382 10726 17434
rect 10726 17382 10738 17434
rect 10738 17382 10752 17434
rect 10776 17382 10790 17434
rect 10790 17382 10802 17434
rect 10802 17382 10832 17434
rect 10856 17382 10866 17434
rect 10866 17382 10912 17434
rect 10616 17380 10672 17382
rect 10696 17380 10752 17382
rect 10776 17380 10832 17382
rect 10856 17380 10912 17382
rect 18616 17434 18672 17436
rect 18696 17434 18752 17436
rect 18776 17434 18832 17436
rect 18856 17434 18912 17436
rect 18616 17382 18662 17434
rect 18662 17382 18672 17434
rect 18696 17382 18726 17434
rect 18726 17382 18738 17434
rect 18738 17382 18752 17434
rect 18776 17382 18790 17434
rect 18790 17382 18802 17434
rect 18802 17382 18832 17434
rect 18856 17382 18866 17434
rect 18866 17382 18912 17434
rect 18616 17380 18672 17382
rect 18696 17380 18752 17382
rect 18776 17380 18832 17382
rect 18856 17380 18912 17382
rect 26616 17434 26672 17436
rect 26696 17434 26752 17436
rect 26776 17434 26832 17436
rect 26856 17434 26912 17436
rect 26616 17382 26662 17434
rect 26662 17382 26672 17434
rect 26696 17382 26726 17434
rect 26726 17382 26738 17434
rect 26738 17382 26752 17434
rect 26776 17382 26790 17434
rect 26790 17382 26802 17434
rect 26802 17382 26832 17434
rect 26856 17382 26866 17434
rect 26866 17382 26912 17434
rect 26616 17380 26672 17382
rect 26696 17380 26752 17382
rect 26776 17380 26832 17382
rect 26856 17380 26912 17382
rect 1956 16890 2012 16892
rect 2036 16890 2092 16892
rect 2116 16890 2172 16892
rect 2196 16890 2252 16892
rect 1956 16838 2002 16890
rect 2002 16838 2012 16890
rect 2036 16838 2066 16890
rect 2066 16838 2078 16890
rect 2078 16838 2092 16890
rect 2116 16838 2130 16890
rect 2130 16838 2142 16890
rect 2142 16838 2172 16890
rect 2196 16838 2206 16890
rect 2206 16838 2252 16890
rect 1956 16836 2012 16838
rect 2036 16836 2092 16838
rect 2116 16836 2172 16838
rect 2196 16836 2252 16838
rect 9956 16890 10012 16892
rect 10036 16890 10092 16892
rect 10116 16890 10172 16892
rect 10196 16890 10252 16892
rect 9956 16838 10002 16890
rect 10002 16838 10012 16890
rect 10036 16838 10066 16890
rect 10066 16838 10078 16890
rect 10078 16838 10092 16890
rect 10116 16838 10130 16890
rect 10130 16838 10142 16890
rect 10142 16838 10172 16890
rect 10196 16838 10206 16890
rect 10206 16838 10252 16890
rect 9956 16836 10012 16838
rect 10036 16836 10092 16838
rect 10116 16836 10172 16838
rect 10196 16836 10252 16838
rect 17956 16890 18012 16892
rect 18036 16890 18092 16892
rect 18116 16890 18172 16892
rect 18196 16890 18252 16892
rect 17956 16838 18002 16890
rect 18002 16838 18012 16890
rect 18036 16838 18066 16890
rect 18066 16838 18078 16890
rect 18078 16838 18092 16890
rect 18116 16838 18130 16890
rect 18130 16838 18142 16890
rect 18142 16838 18172 16890
rect 18196 16838 18206 16890
rect 18206 16838 18252 16890
rect 17956 16836 18012 16838
rect 18036 16836 18092 16838
rect 18116 16836 18172 16838
rect 18196 16836 18252 16838
rect 25956 16890 26012 16892
rect 26036 16890 26092 16892
rect 26116 16890 26172 16892
rect 26196 16890 26252 16892
rect 25956 16838 26002 16890
rect 26002 16838 26012 16890
rect 26036 16838 26066 16890
rect 26066 16838 26078 16890
rect 26078 16838 26092 16890
rect 26116 16838 26130 16890
rect 26130 16838 26142 16890
rect 26142 16838 26172 16890
rect 26196 16838 26206 16890
rect 26206 16838 26252 16890
rect 25956 16836 26012 16838
rect 26036 16836 26092 16838
rect 26116 16836 26172 16838
rect 26196 16836 26252 16838
rect 2616 16346 2672 16348
rect 2696 16346 2752 16348
rect 2776 16346 2832 16348
rect 2856 16346 2912 16348
rect 2616 16294 2662 16346
rect 2662 16294 2672 16346
rect 2696 16294 2726 16346
rect 2726 16294 2738 16346
rect 2738 16294 2752 16346
rect 2776 16294 2790 16346
rect 2790 16294 2802 16346
rect 2802 16294 2832 16346
rect 2856 16294 2866 16346
rect 2866 16294 2912 16346
rect 2616 16292 2672 16294
rect 2696 16292 2752 16294
rect 2776 16292 2832 16294
rect 2856 16292 2912 16294
rect 10616 16346 10672 16348
rect 10696 16346 10752 16348
rect 10776 16346 10832 16348
rect 10856 16346 10912 16348
rect 10616 16294 10662 16346
rect 10662 16294 10672 16346
rect 10696 16294 10726 16346
rect 10726 16294 10738 16346
rect 10738 16294 10752 16346
rect 10776 16294 10790 16346
rect 10790 16294 10802 16346
rect 10802 16294 10832 16346
rect 10856 16294 10866 16346
rect 10866 16294 10912 16346
rect 10616 16292 10672 16294
rect 10696 16292 10752 16294
rect 10776 16292 10832 16294
rect 10856 16292 10912 16294
rect 18616 16346 18672 16348
rect 18696 16346 18752 16348
rect 18776 16346 18832 16348
rect 18856 16346 18912 16348
rect 18616 16294 18662 16346
rect 18662 16294 18672 16346
rect 18696 16294 18726 16346
rect 18726 16294 18738 16346
rect 18738 16294 18752 16346
rect 18776 16294 18790 16346
rect 18790 16294 18802 16346
rect 18802 16294 18832 16346
rect 18856 16294 18866 16346
rect 18866 16294 18912 16346
rect 18616 16292 18672 16294
rect 18696 16292 18752 16294
rect 18776 16292 18832 16294
rect 18856 16292 18912 16294
rect 26616 16346 26672 16348
rect 26696 16346 26752 16348
rect 26776 16346 26832 16348
rect 26856 16346 26912 16348
rect 26616 16294 26662 16346
rect 26662 16294 26672 16346
rect 26696 16294 26726 16346
rect 26726 16294 26738 16346
rect 26738 16294 26752 16346
rect 26776 16294 26790 16346
rect 26790 16294 26802 16346
rect 26802 16294 26832 16346
rect 26856 16294 26866 16346
rect 26866 16294 26912 16346
rect 26616 16292 26672 16294
rect 26696 16292 26752 16294
rect 26776 16292 26832 16294
rect 26856 16292 26912 16294
rect 28354 26968 28410 27024
rect 28354 25336 28410 25392
rect 28354 23704 28410 23760
rect 28354 22072 28410 22128
rect 28354 20440 28410 20496
rect 28354 18808 28410 18864
rect 28354 17176 28410 17232
rect 1956 15802 2012 15804
rect 2036 15802 2092 15804
rect 2116 15802 2172 15804
rect 2196 15802 2252 15804
rect 1956 15750 2002 15802
rect 2002 15750 2012 15802
rect 2036 15750 2066 15802
rect 2066 15750 2078 15802
rect 2078 15750 2092 15802
rect 2116 15750 2130 15802
rect 2130 15750 2142 15802
rect 2142 15750 2172 15802
rect 2196 15750 2206 15802
rect 2206 15750 2252 15802
rect 1956 15748 2012 15750
rect 2036 15748 2092 15750
rect 2116 15748 2172 15750
rect 2196 15748 2252 15750
rect 9956 15802 10012 15804
rect 10036 15802 10092 15804
rect 10116 15802 10172 15804
rect 10196 15802 10252 15804
rect 9956 15750 10002 15802
rect 10002 15750 10012 15802
rect 10036 15750 10066 15802
rect 10066 15750 10078 15802
rect 10078 15750 10092 15802
rect 10116 15750 10130 15802
rect 10130 15750 10142 15802
rect 10142 15750 10172 15802
rect 10196 15750 10206 15802
rect 10206 15750 10252 15802
rect 9956 15748 10012 15750
rect 10036 15748 10092 15750
rect 10116 15748 10172 15750
rect 10196 15748 10252 15750
rect 17956 15802 18012 15804
rect 18036 15802 18092 15804
rect 18116 15802 18172 15804
rect 18196 15802 18252 15804
rect 17956 15750 18002 15802
rect 18002 15750 18012 15802
rect 18036 15750 18066 15802
rect 18066 15750 18078 15802
rect 18078 15750 18092 15802
rect 18116 15750 18130 15802
rect 18130 15750 18142 15802
rect 18142 15750 18172 15802
rect 18196 15750 18206 15802
rect 18206 15750 18252 15802
rect 17956 15748 18012 15750
rect 18036 15748 18092 15750
rect 18116 15748 18172 15750
rect 18196 15748 18252 15750
rect 25956 15802 26012 15804
rect 26036 15802 26092 15804
rect 26116 15802 26172 15804
rect 26196 15802 26252 15804
rect 25956 15750 26002 15802
rect 26002 15750 26012 15802
rect 26036 15750 26066 15802
rect 26066 15750 26078 15802
rect 26078 15750 26092 15802
rect 26116 15750 26130 15802
rect 26130 15750 26142 15802
rect 26142 15750 26172 15802
rect 26196 15750 26206 15802
rect 26206 15750 26252 15802
rect 25956 15748 26012 15750
rect 26036 15748 26092 15750
rect 26116 15748 26172 15750
rect 26196 15748 26252 15750
rect 2616 15258 2672 15260
rect 2696 15258 2752 15260
rect 2776 15258 2832 15260
rect 2856 15258 2912 15260
rect 2616 15206 2662 15258
rect 2662 15206 2672 15258
rect 2696 15206 2726 15258
rect 2726 15206 2738 15258
rect 2738 15206 2752 15258
rect 2776 15206 2790 15258
rect 2790 15206 2802 15258
rect 2802 15206 2832 15258
rect 2856 15206 2866 15258
rect 2866 15206 2912 15258
rect 2616 15204 2672 15206
rect 2696 15204 2752 15206
rect 2776 15204 2832 15206
rect 2856 15204 2912 15206
rect 10616 15258 10672 15260
rect 10696 15258 10752 15260
rect 10776 15258 10832 15260
rect 10856 15258 10912 15260
rect 10616 15206 10662 15258
rect 10662 15206 10672 15258
rect 10696 15206 10726 15258
rect 10726 15206 10738 15258
rect 10738 15206 10752 15258
rect 10776 15206 10790 15258
rect 10790 15206 10802 15258
rect 10802 15206 10832 15258
rect 10856 15206 10866 15258
rect 10866 15206 10912 15258
rect 10616 15204 10672 15206
rect 10696 15204 10752 15206
rect 10776 15204 10832 15206
rect 10856 15204 10912 15206
rect 18616 15258 18672 15260
rect 18696 15258 18752 15260
rect 18776 15258 18832 15260
rect 18856 15258 18912 15260
rect 18616 15206 18662 15258
rect 18662 15206 18672 15258
rect 18696 15206 18726 15258
rect 18726 15206 18738 15258
rect 18738 15206 18752 15258
rect 18776 15206 18790 15258
rect 18790 15206 18802 15258
rect 18802 15206 18832 15258
rect 18856 15206 18866 15258
rect 18866 15206 18912 15258
rect 18616 15204 18672 15206
rect 18696 15204 18752 15206
rect 18776 15204 18832 15206
rect 18856 15204 18912 15206
rect 26616 15258 26672 15260
rect 26696 15258 26752 15260
rect 26776 15258 26832 15260
rect 26856 15258 26912 15260
rect 26616 15206 26662 15258
rect 26662 15206 26672 15258
rect 26696 15206 26726 15258
rect 26726 15206 26738 15258
rect 26738 15206 26752 15258
rect 26776 15206 26790 15258
rect 26790 15206 26802 15258
rect 26802 15206 26832 15258
rect 26856 15206 26866 15258
rect 26866 15206 26912 15258
rect 26616 15204 26672 15206
rect 26696 15204 26752 15206
rect 26776 15204 26832 15206
rect 26856 15204 26912 15206
rect 1956 14714 2012 14716
rect 2036 14714 2092 14716
rect 2116 14714 2172 14716
rect 2196 14714 2252 14716
rect 1956 14662 2002 14714
rect 2002 14662 2012 14714
rect 2036 14662 2066 14714
rect 2066 14662 2078 14714
rect 2078 14662 2092 14714
rect 2116 14662 2130 14714
rect 2130 14662 2142 14714
rect 2142 14662 2172 14714
rect 2196 14662 2206 14714
rect 2206 14662 2252 14714
rect 1956 14660 2012 14662
rect 2036 14660 2092 14662
rect 2116 14660 2172 14662
rect 2196 14660 2252 14662
rect 9956 14714 10012 14716
rect 10036 14714 10092 14716
rect 10116 14714 10172 14716
rect 10196 14714 10252 14716
rect 9956 14662 10002 14714
rect 10002 14662 10012 14714
rect 10036 14662 10066 14714
rect 10066 14662 10078 14714
rect 10078 14662 10092 14714
rect 10116 14662 10130 14714
rect 10130 14662 10142 14714
rect 10142 14662 10172 14714
rect 10196 14662 10206 14714
rect 10206 14662 10252 14714
rect 9956 14660 10012 14662
rect 10036 14660 10092 14662
rect 10116 14660 10172 14662
rect 10196 14660 10252 14662
rect 17956 14714 18012 14716
rect 18036 14714 18092 14716
rect 18116 14714 18172 14716
rect 18196 14714 18252 14716
rect 17956 14662 18002 14714
rect 18002 14662 18012 14714
rect 18036 14662 18066 14714
rect 18066 14662 18078 14714
rect 18078 14662 18092 14714
rect 18116 14662 18130 14714
rect 18130 14662 18142 14714
rect 18142 14662 18172 14714
rect 18196 14662 18206 14714
rect 18206 14662 18252 14714
rect 17956 14660 18012 14662
rect 18036 14660 18092 14662
rect 18116 14660 18172 14662
rect 18196 14660 18252 14662
rect 25956 14714 26012 14716
rect 26036 14714 26092 14716
rect 26116 14714 26172 14716
rect 26196 14714 26252 14716
rect 25956 14662 26002 14714
rect 26002 14662 26012 14714
rect 26036 14662 26066 14714
rect 26066 14662 26078 14714
rect 26078 14662 26092 14714
rect 26116 14662 26130 14714
rect 26130 14662 26142 14714
rect 26142 14662 26172 14714
rect 26196 14662 26206 14714
rect 26206 14662 26252 14714
rect 25956 14660 26012 14662
rect 26036 14660 26092 14662
rect 26116 14660 26172 14662
rect 26196 14660 26252 14662
rect 2616 14170 2672 14172
rect 2696 14170 2752 14172
rect 2776 14170 2832 14172
rect 2856 14170 2912 14172
rect 2616 14118 2662 14170
rect 2662 14118 2672 14170
rect 2696 14118 2726 14170
rect 2726 14118 2738 14170
rect 2738 14118 2752 14170
rect 2776 14118 2790 14170
rect 2790 14118 2802 14170
rect 2802 14118 2832 14170
rect 2856 14118 2866 14170
rect 2866 14118 2912 14170
rect 2616 14116 2672 14118
rect 2696 14116 2752 14118
rect 2776 14116 2832 14118
rect 2856 14116 2912 14118
rect 10616 14170 10672 14172
rect 10696 14170 10752 14172
rect 10776 14170 10832 14172
rect 10856 14170 10912 14172
rect 10616 14118 10662 14170
rect 10662 14118 10672 14170
rect 10696 14118 10726 14170
rect 10726 14118 10738 14170
rect 10738 14118 10752 14170
rect 10776 14118 10790 14170
rect 10790 14118 10802 14170
rect 10802 14118 10832 14170
rect 10856 14118 10866 14170
rect 10866 14118 10912 14170
rect 10616 14116 10672 14118
rect 10696 14116 10752 14118
rect 10776 14116 10832 14118
rect 10856 14116 10912 14118
rect 18616 14170 18672 14172
rect 18696 14170 18752 14172
rect 18776 14170 18832 14172
rect 18856 14170 18912 14172
rect 18616 14118 18662 14170
rect 18662 14118 18672 14170
rect 18696 14118 18726 14170
rect 18726 14118 18738 14170
rect 18738 14118 18752 14170
rect 18776 14118 18790 14170
rect 18790 14118 18802 14170
rect 18802 14118 18832 14170
rect 18856 14118 18866 14170
rect 18866 14118 18912 14170
rect 18616 14116 18672 14118
rect 18696 14116 18752 14118
rect 18776 14116 18832 14118
rect 18856 14116 18912 14118
rect 26616 14170 26672 14172
rect 26696 14170 26752 14172
rect 26776 14170 26832 14172
rect 26856 14170 26912 14172
rect 26616 14118 26662 14170
rect 26662 14118 26672 14170
rect 26696 14118 26726 14170
rect 26726 14118 26738 14170
rect 26738 14118 26752 14170
rect 26776 14118 26790 14170
rect 26790 14118 26802 14170
rect 26802 14118 26832 14170
rect 26856 14118 26866 14170
rect 26866 14118 26912 14170
rect 26616 14116 26672 14118
rect 26696 14116 26752 14118
rect 26776 14116 26832 14118
rect 26856 14116 26912 14118
rect 1956 13626 2012 13628
rect 2036 13626 2092 13628
rect 2116 13626 2172 13628
rect 2196 13626 2252 13628
rect 1956 13574 2002 13626
rect 2002 13574 2012 13626
rect 2036 13574 2066 13626
rect 2066 13574 2078 13626
rect 2078 13574 2092 13626
rect 2116 13574 2130 13626
rect 2130 13574 2142 13626
rect 2142 13574 2172 13626
rect 2196 13574 2206 13626
rect 2206 13574 2252 13626
rect 1956 13572 2012 13574
rect 2036 13572 2092 13574
rect 2116 13572 2172 13574
rect 2196 13572 2252 13574
rect 9956 13626 10012 13628
rect 10036 13626 10092 13628
rect 10116 13626 10172 13628
rect 10196 13626 10252 13628
rect 9956 13574 10002 13626
rect 10002 13574 10012 13626
rect 10036 13574 10066 13626
rect 10066 13574 10078 13626
rect 10078 13574 10092 13626
rect 10116 13574 10130 13626
rect 10130 13574 10142 13626
rect 10142 13574 10172 13626
rect 10196 13574 10206 13626
rect 10206 13574 10252 13626
rect 9956 13572 10012 13574
rect 10036 13572 10092 13574
rect 10116 13572 10172 13574
rect 10196 13572 10252 13574
rect 17956 13626 18012 13628
rect 18036 13626 18092 13628
rect 18116 13626 18172 13628
rect 18196 13626 18252 13628
rect 17956 13574 18002 13626
rect 18002 13574 18012 13626
rect 18036 13574 18066 13626
rect 18066 13574 18078 13626
rect 18078 13574 18092 13626
rect 18116 13574 18130 13626
rect 18130 13574 18142 13626
rect 18142 13574 18172 13626
rect 18196 13574 18206 13626
rect 18206 13574 18252 13626
rect 17956 13572 18012 13574
rect 18036 13572 18092 13574
rect 18116 13572 18172 13574
rect 18196 13572 18252 13574
rect 25956 13626 26012 13628
rect 26036 13626 26092 13628
rect 26116 13626 26172 13628
rect 26196 13626 26252 13628
rect 25956 13574 26002 13626
rect 26002 13574 26012 13626
rect 26036 13574 26066 13626
rect 26066 13574 26078 13626
rect 26078 13574 26092 13626
rect 26116 13574 26130 13626
rect 26130 13574 26142 13626
rect 26142 13574 26172 13626
rect 26196 13574 26206 13626
rect 26206 13574 26252 13626
rect 25956 13572 26012 13574
rect 26036 13572 26092 13574
rect 26116 13572 26172 13574
rect 26196 13572 26252 13574
rect 2616 13082 2672 13084
rect 2696 13082 2752 13084
rect 2776 13082 2832 13084
rect 2856 13082 2912 13084
rect 2616 13030 2662 13082
rect 2662 13030 2672 13082
rect 2696 13030 2726 13082
rect 2726 13030 2738 13082
rect 2738 13030 2752 13082
rect 2776 13030 2790 13082
rect 2790 13030 2802 13082
rect 2802 13030 2832 13082
rect 2856 13030 2866 13082
rect 2866 13030 2912 13082
rect 2616 13028 2672 13030
rect 2696 13028 2752 13030
rect 2776 13028 2832 13030
rect 2856 13028 2912 13030
rect 10616 13082 10672 13084
rect 10696 13082 10752 13084
rect 10776 13082 10832 13084
rect 10856 13082 10912 13084
rect 10616 13030 10662 13082
rect 10662 13030 10672 13082
rect 10696 13030 10726 13082
rect 10726 13030 10738 13082
rect 10738 13030 10752 13082
rect 10776 13030 10790 13082
rect 10790 13030 10802 13082
rect 10802 13030 10832 13082
rect 10856 13030 10866 13082
rect 10866 13030 10912 13082
rect 10616 13028 10672 13030
rect 10696 13028 10752 13030
rect 10776 13028 10832 13030
rect 10856 13028 10912 13030
rect 18616 13082 18672 13084
rect 18696 13082 18752 13084
rect 18776 13082 18832 13084
rect 18856 13082 18912 13084
rect 18616 13030 18662 13082
rect 18662 13030 18672 13082
rect 18696 13030 18726 13082
rect 18726 13030 18738 13082
rect 18738 13030 18752 13082
rect 18776 13030 18790 13082
rect 18790 13030 18802 13082
rect 18802 13030 18832 13082
rect 18856 13030 18866 13082
rect 18866 13030 18912 13082
rect 18616 13028 18672 13030
rect 18696 13028 18752 13030
rect 18776 13028 18832 13030
rect 18856 13028 18912 13030
rect 26616 13082 26672 13084
rect 26696 13082 26752 13084
rect 26776 13082 26832 13084
rect 26856 13082 26912 13084
rect 26616 13030 26662 13082
rect 26662 13030 26672 13082
rect 26696 13030 26726 13082
rect 26726 13030 26738 13082
rect 26738 13030 26752 13082
rect 26776 13030 26790 13082
rect 26790 13030 26802 13082
rect 26802 13030 26832 13082
rect 26856 13030 26866 13082
rect 26866 13030 26912 13082
rect 26616 13028 26672 13030
rect 26696 13028 26752 13030
rect 26776 13028 26832 13030
rect 26856 13028 26912 13030
rect 28354 15564 28410 15600
rect 28354 15544 28356 15564
rect 28356 15544 28408 15564
rect 28408 15544 28410 15564
rect 28354 13912 28410 13968
rect 1956 12538 2012 12540
rect 2036 12538 2092 12540
rect 2116 12538 2172 12540
rect 2196 12538 2252 12540
rect 1956 12486 2002 12538
rect 2002 12486 2012 12538
rect 2036 12486 2066 12538
rect 2066 12486 2078 12538
rect 2078 12486 2092 12538
rect 2116 12486 2130 12538
rect 2130 12486 2142 12538
rect 2142 12486 2172 12538
rect 2196 12486 2206 12538
rect 2206 12486 2252 12538
rect 1956 12484 2012 12486
rect 2036 12484 2092 12486
rect 2116 12484 2172 12486
rect 2196 12484 2252 12486
rect 9956 12538 10012 12540
rect 10036 12538 10092 12540
rect 10116 12538 10172 12540
rect 10196 12538 10252 12540
rect 9956 12486 10002 12538
rect 10002 12486 10012 12538
rect 10036 12486 10066 12538
rect 10066 12486 10078 12538
rect 10078 12486 10092 12538
rect 10116 12486 10130 12538
rect 10130 12486 10142 12538
rect 10142 12486 10172 12538
rect 10196 12486 10206 12538
rect 10206 12486 10252 12538
rect 9956 12484 10012 12486
rect 10036 12484 10092 12486
rect 10116 12484 10172 12486
rect 10196 12484 10252 12486
rect 17956 12538 18012 12540
rect 18036 12538 18092 12540
rect 18116 12538 18172 12540
rect 18196 12538 18252 12540
rect 17956 12486 18002 12538
rect 18002 12486 18012 12538
rect 18036 12486 18066 12538
rect 18066 12486 18078 12538
rect 18078 12486 18092 12538
rect 18116 12486 18130 12538
rect 18130 12486 18142 12538
rect 18142 12486 18172 12538
rect 18196 12486 18206 12538
rect 18206 12486 18252 12538
rect 17956 12484 18012 12486
rect 18036 12484 18092 12486
rect 18116 12484 18172 12486
rect 18196 12484 18252 12486
rect 25956 12538 26012 12540
rect 26036 12538 26092 12540
rect 26116 12538 26172 12540
rect 26196 12538 26252 12540
rect 25956 12486 26002 12538
rect 26002 12486 26012 12538
rect 26036 12486 26066 12538
rect 26066 12486 26078 12538
rect 26078 12486 26092 12538
rect 26116 12486 26130 12538
rect 26130 12486 26142 12538
rect 26142 12486 26172 12538
rect 26196 12486 26206 12538
rect 26206 12486 26252 12538
rect 25956 12484 26012 12486
rect 26036 12484 26092 12486
rect 26116 12484 26172 12486
rect 26196 12484 26252 12486
rect 2616 11994 2672 11996
rect 2696 11994 2752 11996
rect 2776 11994 2832 11996
rect 2856 11994 2912 11996
rect 2616 11942 2662 11994
rect 2662 11942 2672 11994
rect 2696 11942 2726 11994
rect 2726 11942 2738 11994
rect 2738 11942 2752 11994
rect 2776 11942 2790 11994
rect 2790 11942 2802 11994
rect 2802 11942 2832 11994
rect 2856 11942 2866 11994
rect 2866 11942 2912 11994
rect 2616 11940 2672 11942
rect 2696 11940 2752 11942
rect 2776 11940 2832 11942
rect 2856 11940 2912 11942
rect 10616 11994 10672 11996
rect 10696 11994 10752 11996
rect 10776 11994 10832 11996
rect 10856 11994 10912 11996
rect 10616 11942 10662 11994
rect 10662 11942 10672 11994
rect 10696 11942 10726 11994
rect 10726 11942 10738 11994
rect 10738 11942 10752 11994
rect 10776 11942 10790 11994
rect 10790 11942 10802 11994
rect 10802 11942 10832 11994
rect 10856 11942 10866 11994
rect 10866 11942 10912 11994
rect 10616 11940 10672 11942
rect 10696 11940 10752 11942
rect 10776 11940 10832 11942
rect 10856 11940 10912 11942
rect 18616 11994 18672 11996
rect 18696 11994 18752 11996
rect 18776 11994 18832 11996
rect 18856 11994 18912 11996
rect 18616 11942 18662 11994
rect 18662 11942 18672 11994
rect 18696 11942 18726 11994
rect 18726 11942 18738 11994
rect 18738 11942 18752 11994
rect 18776 11942 18790 11994
rect 18790 11942 18802 11994
rect 18802 11942 18832 11994
rect 18856 11942 18866 11994
rect 18866 11942 18912 11994
rect 18616 11940 18672 11942
rect 18696 11940 18752 11942
rect 18776 11940 18832 11942
rect 18856 11940 18912 11942
rect 26616 11994 26672 11996
rect 26696 11994 26752 11996
rect 26776 11994 26832 11996
rect 26856 11994 26912 11996
rect 26616 11942 26662 11994
rect 26662 11942 26672 11994
rect 26696 11942 26726 11994
rect 26726 11942 26738 11994
rect 26738 11942 26752 11994
rect 26776 11942 26790 11994
rect 26790 11942 26802 11994
rect 26802 11942 26832 11994
rect 26856 11942 26866 11994
rect 26866 11942 26912 11994
rect 26616 11940 26672 11942
rect 26696 11940 26752 11942
rect 26776 11940 26832 11942
rect 26856 11940 26912 11942
rect 1956 11450 2012 11452
rect 2036 11450 2092 11452
rect 2116 11450 2172 11452
rect 2196 11450 2252 11452
rect 1956 11398 2002 11450
rect 2002 11398 2012 11450
rect 2036 11398 2066 11450
rect 2066 11398 2078 11450
rect 2078 11398 2092 11450
rect 2116 11398 2130 11450
rect 2130 11398 2142 11450
rect 2142 11398 2172 11450
rect 2196 11398 2206 11450
rect 2206 11398 2252 11450
rect 1956 11396 2012 11398
rect 2036 11396 2092 11398
rect 2116 11396 2172 11398
rect 2196 11396 2252 11398
rect 9956 11450 10012 11452
rect 10036 11450 10092 11452
rect 10116 11450 10172 11452
rect 10196 11450 10252 11452
rect 9956 11398 10002 11450
rect 10002 11398 10012 11450
rect 10036 11398 10066 11450
rect 10066 11398 10078 11450
rect 10078 11398 10092 11450
rect 10116 11398 10130 11450
rect 10130 11398 10142 11450
rect 10142 11398 10172 11450
rect 10196 11398 10206 11450
rect 10206 11398 10252 11450
rect 9956 11396 10012 11398
rect 10036 11396 10092 11398
rect 10116 11396 10172 11398
rect 10196 11396 10252 11398
rect 17956 11450 18012 11452
rect 18036 11450 18092 11452
rect 18116 11450 18172 11452
rect 18196 11450 18252 11452
rect 17956 11398 18002 11450
rect 18002 11398 18012 11450
rect 18036 11398 18066 11450
rect 18066 11398 18078 11450
rect 18078 11398 18092 11450
rect 18116 11398 18130 11450
rect 18130 11398 18142 11450
rect 18142 11398 18172 11450
rect 18196 11398 18206 11450
rect 18206 11398 18252 11450
rect 17956 11396 18012 11398
rect 18036 11396 18092 11398
rect 18116 11396 18172 11398
rect 18196 11396 18252 11398
rect 25956 11450 26012 11452
rect 26036 11450 26092 11452
rect 26116 11450 26172 11452
rect 26196 11450 26252 11452
rect 25956 11398 26002 11450
rect 26002 11398 26012 11450
rect 26036 11398 26066 11450
rect 26066 11398 26078 11450
rect 26078 11398 26092 11450
rect 26116 11398 26130 11450
rect 26130 11398 26142 11450
rect 26142 11398 26172 11450
rect 26196 11398 26206 11450
rect 26206 11398 26252 11450
rect 25956 11396 26012 11398
rect 26036 11396 26092 11398
rect 26116 11396 26172 11398
rect 26196 11396 26252 11398
rect 2616 10906 2672 10908
rect 2696 10906 2752 10908
rect 2776 10906 2832 10908
rect 2856 10906 2912 10908
rect 2616 10854 2662 10906
rect 2662 10854 2672 10906
rect 2696 10854 2726 10906
rect 2726 10854 2738 10906
rect 2738 10854 2752 10906
rect 2776 10854 2790 10906
rect 2790 10854 2802 10906
rect 2802 10854 2832 10906
rect 2856 10854 2866 10906
rect 2866 10854 2912 10906
rect 2616 10852 2672 10854
rect 2696 10852 2752 10854
rect 2776 10852 2832 10854
rect 2856 10852 2912 10854
rect 10616 10906 10672 10908
rect 10696 10906 10752 10908
rect 10776 10906 10832 10908
rect 10856 10906 10912 10908
rect 10616 10854 10662 10906
rect 10662 10854 10672 10906
rect 10696 10854 10726 10906
rect 10726 10854 10738 10906
rect 10738 10854 10752 10906
rect 10776 10854 10790 10906
rect 10790 10854 10802 10906
rect 10802 10854 10832 10906
rect 10856 10854 10866 10906
rect 10866 10854 10912 10906
rect 10616 10852 10672 10854
rect 10696 10852 10752 10854
rect 10776 10852 10832 10854
rect 10856 10852 10912 10854
rect 18616 10906 18672 10908
rect 18696 10906 18752 10908
rect 18776 10906 18832 10908
rect 18856 10906 18912 10908
rect 18616 10854 18662 10906
rect 18662 10854 18672 10906
rect 18696 10854 18726 10906
rect 18726 10854 18738 10906
rect 18738 10854 18752 10906
rect 18776 10854 18790 10906
rect 18790 10854 18802 10906
rect 18802 10854 18832 10906
rect 18856 10854 18866 10906
rect 18866 10854 18912 10906
rect 18616 10852 18672 10854
rect 18696 10852 18752 10854
rect 18776 10852 18832 10854
rect 18856 10852 18912 10854
rect 26616 10906 26672 10908
rect 26696 10906 26752 10908
rect 26776 10906 26832 10908
rect 26856 10906 26912 10908
rect 26616 10854 26662 10906
rect 26662 10854 26672 10906
rect 26696 10854 26726 10906
rect 26726 10854 26738 10906
rect 26738 10854 26752 10906
rect 26776 10854 26790 10906
rect 26790 10854 26802 10906
rect 26802 10854 26832 10906
rect 26856 10854 26866 10906
rect 26866 10854 26912 10906
rect 26616 10852 26672 10854
rect 26696 10852 26752 10854
rect 26776 10852 26832 10854
rect 26856 10852 26912 10854
rect 1956 10362 2012 10364
rect 2036 10362 2092 10364
rect 2116 10362 2172 10364
rect 2196 10362 2252 10364
rect 1956 10310 2002 10362
rect 2002 10310 2012 10362
rect 2036 10310 2066 10362
rect 2066 10310 2078 10362
rect 2078 10310 2092 10362
rect 2116 10310 2130 10362
rect 2130 10310 2142 10362
rect 2142 10310 2172 10362
rect 2196 10310 2206 10362
rect 2206 10310 2252 10362
rect 1956 10308 2012 10310
rect 2036 10308 2092 10310
rect 2116 10308 2172 10310
rect 2196 10308 2252 10310
rect 9956 10362 10012 10364
rect 10036 10362 10092 10364
rect 10116 10362 10172 10364
rect 10196 10362 10252 10364
rect 9956 10310 10002 10362
rect 10002 10310 10012 10362
rect 10036 10310 10066 10362
rect 10066 10310 10078 10362
rect 10078 10310 10092 10362
rect 10116 10310 10130 10362
rect 10130 10310 10142 10362
rect 10142 10310 10172 10362
rect 10196 10310 10206 10362
rect 10206 10310 10252 10362
rect 9956 10308 10012 10310
rect 10036 10308 10092 10310
rect 10116 10308 10172 10310
rect 10196 10308 10252 10310
rect 17956 10362 18012 10364
rect 18036 10362 18092 10364
rect 18116 10362 18172 10364
rect 18196 10362 18252 10364
rect 17956 10310 18002 10362
rect 18002 10310 18012 10362
rect 18036 10310 18066 10362
rect 18066 10310 18078 10362
rect 18078 10310 18092 10362
rect 18116 10310 18130 10362
rect 18130 10310 18142 10362
rect 18142 10310 18172 10362
rect 18196 10310 18206 10362
rect 18206 10310 18252 10362
rect 17956 10308 18012 10310
rect 18036 10308 18092 10310
rect 18116 10308 18172 10310
rect 18196 10308 18252 10310
rect 25956 10362 26012 10364
rect 26036 10362 26092 10364
rect 26116 10362 26172 10364
rect 26196 10362 26252 10364
rect 25956 10310 26002 10362
rect 26002 10310 26012 10362
rect 26036 10310 26066 10362
rect 26066 10310 26078 10362
rect 26078 10310 26092 10362
rect 26116 10310 26130 10362
rect 26130 10310 26142 10362
rect 26142 10310 26172 10362
rect 26196 10310 26206 10362
rect 26206 10310 26252 10362
rect 25956 10308 26012 10310
rect 26036 10308 26092 10310
rect 26116 10308 26172 10310
rect 26196 10308 26252 10310
rect 2616 9818 2672 9820
rect 2696 9818 2752 9820
rect 2776 9818 2832 9820
rect 2856 9818 2912 9820
rect 2616 9766 2662 9818
rect 2662 9766 2672 9818
rect 2696 9766 2726 9818
rect 2726 9766 2738 9818
rect 2738 9766 2752 9818
rect 2776 9766 2790 9818
rect 2790 9766 2802 9818
rect 2802 9766 2832 9818
rect 2856 9766 2866 9818
rect 2866 9766 2912 9818
rect 2616 9764 2672 9766
rect 2696 9764 2752 9766
rect 2776 9764 2832 9766
rect 2856 9764 2912 9766
rect 10616 9818 10672 9820
rect 10696 9818 10752 9820
rect 10776 9818 10832 9820
rect 10856 9818 10912 9820
rect 10616 9766 10662 9818
rect 10662 9766 10672 9818
rect 10696 9766 10726 9818
rect 10726 9766 10738 9818
rect 10738 9766 10752 9818
rect 10776 9766 10790 9818
rect 10790 9766 10802 9818
rect 10802 9766 10832 9818
rect 10856 9766 10866 9818
rect 10866 9766 10912 9818
rect 10616 9764 10672 9766
rect 10696 9764 10752 9766
rect 10776 9764 10832 9766
rect 10856 9764 10912 9766
rect 18616 9818 18672 9820
rect 18696 9818 18752 9820
rect 18776 9818 18832 9820
rect 18856 9818 18912 9820
rect 18616 9766 18662 9818
rect 18662 9766 18672 9818
rect 18696 9766 18726 9818
rect 18726 9766 18738 9818
rect 18738 9766 18752 9818
rect 18776 9766 18790 9818
rect 18790 9766 18802 9818
rect 18802 9766 18832 9818
rect 18856 9766 18866 9818
rect 18866 9766 18912 9818
rect 18616 9764 18672 9766
rect 18696 9764 18752 9766
rect 18776 9764 18832 9766
rect 18856 9764 18912 9766
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 9956 9274 10012 9276
rect 10036 9274 10092 9276
rect 10116 9274 10172 9276
rect 10196 9274 10252 9276
rect 9956 9222 10002 9274
rect 10002 9222 10012 9274
rect 10036 9222 10066 9274
rect 10066 9222 10078 9274
rect 10078 9222 10092 9274
rect 10116 9222 10130 9274
rect 10130 9222 10142 9274
rect 10142 9222 10172 9274
rect 10196 9222 10206 9274
rect 10206 9222 10252 9274
rect 9956 9220 10012 9222
rect 10036 9220 10092 9222
rect 10116 9220 10172 9222
rect 10196 9220 10252 9222
rect 17956 9274 18012 9276
rect 18036 9274 18092 9276
rect 18116 9274 18172 9276
rect 18196 9274 18252 9276
rect 17956 9222 18002 9274
rect 18002 9222 18012 9274
rect 18036 9222 18066 9274
rect 18066 9222 18078 9274
rect 18078 9222 18092 9274
rect 18116 9222 18130 9274
rect 18130 9222 18142 9274
rect 18142 9222 18172 9274
rect 18196 9222 18206 9274
rect 18206 9222 18252 9274
rect 17956 9220 18012 9222
rect 18036 9220 18092 9222
rect 18116 9220 18172 9222
rect 18196 9220 18252 9222
rect 25956 9274 26012 9276
rect 26036 9274 26092 9276
rect 26116 9274 26172 9276
rect 26196 9274 26252 9276
rect 25956 9222 26002 9274
rect 26002 9222 26012 9274
rect 26036 9222 26066 9274
rect 26066 9222 26078 9274
rect 26078 9222 26092 9274
rect 26116 9222 26130 9274
rect 26130 9222 26142 9274
rect 26142 9222 26172 9274
rect 26196 9222 26206 9274
rect 26206 9222 26252 9274
rect 25956 9220 26012 9222
rect 26036 9220 26092 9222
rect 26116 9220 26172 9222
rect 26196 9220 26252 9222
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 10616 8730 10672 8732
rect 10696 8730 10752 8732
rect 10776 8730 10832 8732
rect 10856 8730 10912 8732
rect 10616 8678 10662 8730
rect 10662 8678 10672 8730
rect 10696 8678 10726 8730
rect 10726 8678 10738 8730
rect 10738 8678 10752 8730
rect 10776 8678 10790 8730
rect 10790 8678 10802 8730
rect 10802 8678 10832 8730
rect 10856 8678 10866 8730
rect 10866 8678 10912 8730
rect 10616 8676 10672 8678
rect 10696 8676 10752 8678
rect 10776 8676 10832 8678
rect 10856 8676 10912 8678
rect 18616 8730 18672 8732
rect 18696 8730 18752 8732
rect 18776 8730 18832 8732
rect 18856 8730 18912 8732
rect 18616 8678 18662 8730
rect 18662 8678 18672 8730
rect 18696 8678 18726 8730
rect 18726 8678 18738 8730
rect 18738 8678 18752 8730
rect 18776 8678 18790 8730
rect 18790 8678 18802 8730
rect 18802 8678 18832 8730
rect 18856 8678 18866 8730
rect 18866 8678 18912 8730
rect 18616 8676 18672 8678
rect 18696 8676 18752 8678
rect 18776 8676 18832 8678
rect 18856 8676 18912 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 9956 8186 10012 8188
rect 10036 8186 10092 8188
rect 10116 8186 10172 8188
rect 10196 8186 10252 8188
rect 9956 8134 10002 8186
rect 10002 8134 10012 8186
rect 10036 8134 10066 8186
rect 10066 8134 10078 8186
rect 10078 8134 10092 8186
rect 10116 8134 10130 8186
rect 10130 8134 10142 8186
rect 10142 8134 10172 8186
rect 10196 8134 10206 8186
rect 10206 8134 10252 8186
rect 9956 8132 10012 8134
rect 10036 8132 10092 8134
rect 10116 8132 10172 8134
rect 10196 8132 10252 8134
rect 17956 8186 18012 8188
rect 18036 8186 18092 8188
rect 18116 8186 18172 8188
rect 18196 8186 18252 8188
rect 17956 8134 18002 8186
rect 18002 8134 18012 8186
rect 18036 8134 18066 8186
rect 18066 8134 18078 8186
rect 18078 8134 18092 8186
rect 18116 8134 18130 8186
rect 18130 8134 18142 8186
rect 18142 8134 18172 8186
rect 18196 8134 18206 8186
rect 18206 8134 18252 8186
rect 17956 8132 18012 8134
rect 18036 8132 18092 8134
rect 18116 8132 18172 8134
rect 18196 8132 18252 8134
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 26616 9818 26672 9820
rect 26696 9818 26752 9820
rect 26776 9818 26832 9820
rect 26856 9818 26912 9820
rect 26616 9766 26662 9818
rect 26662 9766 26672 9818
rect 26696 9766 26726 9818
rect 26726 9766 26738 9818
rect 26738 9766 26752 9818
rect 26776 9766 26790 9818
rect 26790 9766 26802 9818
rect 26802 9766 26832 9818
rect 26856 9766 26866 9818
rect 26866 9766 26912 9818
rect 26616 9764 26672 9766
rect 26696 9764 26752 9766
rect 26776 9764 26832 9766
rect 26856 9764 26912 9766
rect 26616 8730 26672 8732
rect 26696 8730 26752 8732
rect 26776 8730 26832 8732
rect 26856 8730 26912 8732
rect 26616 8678 26662 8730
rect 26662 8678 26672 8730
rect 26696 8678 26726 8730
rect 26726 8678 26738 8730
rect 26738 8678 26752 8730
rect 26776 8678 26790 8730
rect 26790 8678 26802 8730
rect 26802 8678 26832 8730
rect 26856 8678 26866 8730
rect 26866 8678 26912 8730
rect 26616 8676 26672 8678
rect 26696 8676 26752 8678
rect 26776 8676 26832 8678
rect 26856 8676 26912 8678
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 10616 7642 10672 7644
rect 10696 7642 10752 7644
rect 10776 7642 10832 7644
rect 10856 7642 10912 7644
rect 10616 7590 10662 7642
rect 10662 7590 10672 7642
rect 10696 7590 10726 7642
rect 10726 7590 10738 7642
rect 10738 7590 10752 7642
rect 10776 7590 10790 7642
rect 10790 7590 10802 7642
rect 10802 7590 10832 7642
rect 10856 7590 10866 7642
rect 10866 7590 10912 7642
rect 10616 7588 10672 7590
rect 10696 7588 10752 7590
rect 10776 7588 10832 7590
rect 10856 7588 10912 7590
rect 18616 7642 18672 7644
rect 18696 7642 18752 7644
rect 18776 7642 18832 7644
rect 18856 7642 18912 7644
rect 18616 7590 18662 7642
rect 18662 7590 18672 7642
rect 18696 7590 18726 7642
rect 18726 7590 18738 7642
rect 18738 7590 18752 7642
rect 18776 7590 18790 7642
rect 18790 7590 18802 7642
rect 18802 7590 18832 7642
rect 18856 7590 18866 7642
rect 18866 7590 18912 7642
rect 18616 7588 18672 7590
rect 18696 7588 18752 7590
rect 18776 7588 18832 7590
rect 18856 7588 18912 7590
rect 26616 7642 26672 7644
rect 26696 7642 26752 7644
rect 26776 7642 26832 7644
rect 26856 7642 26912 7644
rect 26616 7590 26662 7642
rect 26662 7590 26672 7642
rect 26696 7590 26726 7642
rect 26726 7590 26738 7642
rect 26738 7590 26752 7642
rect 26776 7590 26790 7642
rect 26790 7590 26802 7642
rect 26802 7590 26832 7642
rect 26856 7590 26866 7642
rect 26866 7590 26912 7642
rect 26616 7588 26672 7590
rect 26696 7588 26752 7590
rect 26776 7588 26832 7590
rect 26856 7588 26912 7590
rect 846 7520 902 7576
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 9956 7098 10012 7100
rect 10036 7098 10092 7100
rect 10116 7098 10172 7100
rect 10196 7098 10252 7100
rect 9956 7046 10002 7098
rect 10002 7046 10012 7098
rect 10036 7046 10066 7098
rect 10066 7046 10078 7098
rect 10078 7046 10092 7098
rect 10116 7046 10130 7098
rect 10130 7046 10142 7098
rect 10142 7046 10172 7098
rect 10196 7046 10206 7098
rect 10206 7046 10252 7098
rect 9956 7044 10012 7046
rect 10036 7044 10092 7046
rect 10116 7044 10172 7046
rect 10196 7044 10252 7046
rect 17956 7098 18012 7100
rect 18036 7098 18092 7100
rect 18116 7098 18172 7100
rect 18196 7098 18252 7100
rect 17956 7046 18002 7098
rect 18002 7046 18012 7098
rect 18036 7046 18066 7098
rect 18066 7046 18078 7098
rect 18078 7046 18092 7098
rect 18116 7046 18130 7098
rect 18130 7046 18142 7098
rect 18142 7046 18172 7098
rect 18196 7046 18206 7098
rect 18206 7046 18252 7098
rect 17956 7044 18012 7046
rect 18036 7044 18092 7046
rect 18116 7044 18172 7046
rect 18196 7044 18252 7046
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 10616 6554 10672 6556
rect 10696 6554 10752 6556
rect 10776 6554 10832 6556
rect 10856 6554 10912 6556
rect 10616 6502 10662 6554
rect 10662 6502 10672 6554
rect 10696 6502 10726 6554
rect 10726 6502 10738 6554
rect 10738 6502 10752 6554
rect 10776 6502 10790 6554
rect 10790 6502 10802 6554
rect 10802 6502 10832 6554
rect 10856 6502 10866 6554
rect 10866 6502 10912 6554
rect 10616 6500 10672 6502
rect 10696 6500 10752 6502
rect 10776 6500 10832 6502
rect 10856 6500 10912 6502
rect 18616 6554 18672 6556
rect 18696 6554 18752 6556
rect 18776 6554 18832 6556
rect 18856 6554 18912 6556
rect 18616 6502 18662 6554
rect 18662 6502 18672 6554
rect 18696 6502 18726 6554
rect 18726 6502 18738 6554
rect 18738 6502 18752 6554
rect 18776 6502 18790 6554
rect 18790 6502 18802 6554
rect 18802 6502 18832 6554
rect 18856 6502 18866 6554
rect 18866 6502 18912 6554
rect 18616 6500 18672 6502
rect 18696 6500 18752 6502
rect 18776 6500 18832 6502
rect 18856 6500 18912 6502
rect 26616 6554 26672 6556
rect 26696 6554 26752 6556
rect 26776 6554 26832 6556
rect 26856 6554 26912 6556
rect 26616 6502 26662 6554
rect 26662 6502 26672 6554
rect 26696 6502 26726 6554
rect 26726 6502 26738 6554
rect 26738 6502 26752 6554
rect 26776 6502 26790 6554
rect 26790 6502 26802 6554
rect 26802 6502 26832 6554
rect 26856 6502 26866 6554
rect 26866 6502 26912 6554
rect 26616 6500 26672 6502
rect 26696 6500 26752 6502
rect 26776 6500 26832 6502
rect 26856 6500 26912 6502
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 9956 6010 10012 6012
rect 10036 6010 10092 6012
rect 10116 6010 10172 6012
rect 10196 6010 10252 6012
rect 9956 5958 10002 6010
rect 10002 5958 10012 6010
rect 10036 5958 10066 6010
rect 10066 5958 10078 6010
rect 10078 5958 10092 6010
rect 10116 5958 10130 6010
rect 10130 5958 10142 6010
rect 10142 5958 10172 6010
rect 10196 5958 10206 6010
rect 10206 5958 10252 6010
rect 9956 5956 10012 5958
rect 10036 5956 10092 5958
rect 10116 5956 10172 5958
rect 10196 5956 10252 5958
rect 17956 6010 18012 6012
rect 18036 6010 18092 6012
rect 18116 6010 18172 6012
rect 18196 6010 18252 6012
rect 17956 5958 18002 6010
rect 18002 5958 18012 6010
rect 18036 5958 18066 6010
rect 18066 5958 18078 6010
rect 18078 5958 18092 6010
rect 18116 5958 18130 6010
rect 18130 5958 18142 6010
rect 18142 5958 18172 6010
rect 18196 5958 18206 6010
rect 18206 5958 18252 6010
rect 17956 5956 18012 5958
rect 18036 5956 18092 5958
rect 18116 5956 18172 5958
rect 18196 5956 18252 5958
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 10616 5466 10672 5468
rect 10696 5466 10752 5468
rect 10776 5466 10832 5468
rect 10856 5466 10912 5468
rect 10616 5414 10662 5466
rect 10662 5414 10672 5466
rect 10696 5414 10726 5466
rect 10726 5414 10738 5466
rect 10738 5414 10752 5466
rect 10776 5414 10790 5466
rect 10790 5414 10802 5466
rect 10802 5414 10832 5466
rect 10856 5414 10866 5466
rect 10866 5414 10912 5466
rect 10616 5412 10672 5414
rect 10696 5412 10752 5414
rect 10776 5412 10832 5414
rect 10856 5412 10912 5414
rect 18616 5466 18672 5468
rect 18696 5466 18752 5468
rect 18776 5466 18832 5468
rect 18856 5466 18912 5468
rect 18616 5414 18662 5466
rect 18662 5414 18672 5466
rect 18696 5414 18726 5466
rect 18726 5414 18738 5466
rect 18738 5414 18752 5466
rect 18776 5414 18790 5466
rect 18790 5414 18802 5466
rect 18802 5414 18832 5466
rect 18856 5414 18866 5466
rect 18866 5414 18912 5466
rect 18616 5412 18672 5414
rect 18696 5412 18752 5414
rect 18776 5412 18832 5414
rect 18856 5412 18912 5414
rect 26616 5466 26672 5468
rect 26696 5466 26752 5468
rect 26776 5466 26832 5468
rect 26856 5466 26912 5468
rect 26616 5414 26662 5466
rect 26662 5414 26672 5466
rect 26696 5414 26726 5466
rect 26726 5414 26738 5466
rect 26738 5414 26752 5466
rect 26776 5414 26790 5466
rect 26790 5414 26802 5466
rect 26802 5414 26832 5466
rect 26856 5414 26866 5466
rect 26866 5414 26912 5466
rect 26616 5412 26672 5414
rect 26696 5412 26752 5414
rect 26776 5412 26832 5414
rect 26856 5412 26912 5414
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 9956 4922 10012 4924
rect 10036 4922 10092 4924
rect 10116 4922 10172 4924
rect 10196 4922 10252 4924
rect 9956 4870 10002 4922
rect 10002 4870 10012 4922
rect 10036 4870 10066 4922
rect 10066 4870 10078 4922
rect 10078 4870 10092 4922
rect 10116 4870 10130 4922
rect 10130 4870 10142 4922
rect 10142 4870 10172 4922
rect 10196 4870 10206 4922
rect 10206 4870 10252 4922
rect 9956 4868 10012 4870
rect 10036 4868 10092 4870
rect 10116 4868 10172 4870
rect 10196 4868 10252 4870
rect 17956 4922 18012 4924
rect 18036 4922 18092 4924
rect 18116 4922 18172 4924
rect 18196 4922 18252 4924
rect 17956 4870 18002 4922
rect 18002 4870 18012 4922
rect 18036 4870 18066 4922
rect 18066 4870 18078 4922
rect 18078 4870 18092 4922
rect 18116 4870 18130 4922
rect 18130 4870 18142 4922
rect 18142 4870 18172 4922
rect 18196 4870 18206 4922
rect 18206 4870 18252 4922
rect 17956 4868 18012 4870
rect 18036 4868 18092 4870
rect 18116 4868 18172 4870
rect 18196 4868 18252 4870
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 10616 4378 10672 4380
rect 10696 4378 10752 4380
rect 10776 4378 10832 4380
rect 10856 4378 10912 4380
rect 10616 4326 10662 4378
rect 10662 4326 10672 4378
rect 10696 4326 10726 4378
rect 10726 4326 10738 4378
rect 10738 4326 10752 4378
rect 10776 4326 10790 4378
rect 10790 4326 10802 4378
rect 10802 4326 10832 4378
rect 10856 4326 10866 4378
rect 10866 4326 10912 4378
rect 10616 4324 10672 4326
rect 10696 4324 10752 4326
rect 10776 4324 10832 4326
rect 10856 4324 10912 4326
rect 18616 4378 18672 4380
rect 18696 4378 18752 4380
rect 18776 4378 18832 4380
rect 18856 4378 18912 4380
rect 18616 4326 18662 4378
rect 18662 4326 18672 4378
rect 18696 4326 18726 4378
rect 18726 4326 18738 4378
rect 18738 4326 18752 4378
rect 18776 4326 18790 4378
rect 18790 4326 18802 4378
rect 18802 4326 18832 4378
rect 18856 4326 18866 4378
rect 18866 4326 18912 4378
rect 18616 4324 18672 4326
rect 18696 4324 18752 4326
rect 18776 4324 18832 4326
rect 18856 4324 18912 4326
rect 26616 4378 26672 4380
rect 26696 4378 26752 4380
rect 26776 4378 26832 4380
rect 26856 4378 26912 4380
rect 26616 4326 26662 4378
rect 26662 4326 26672 4378
rect 26696 4326 26726 4378
rect 26726 4326 26738 4378
rect 26738 4326 26752 4378
rect 26776 4326 26790 4378
rect 26790 4326 26802 4378
rect 26802 4326 26832 4378
rect 26856 4326 26866 4378
rect 26866 4326 26912 4378
rect 26616 4324 26672 4326
rect 26696 4324 26752 4326
rect 26776 4324 26832 4326
rect 26856 4324 26912 4326
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 9956 3834 10012 3836
rect 10036 3834 10092 3836
rect 10116 3834 10172 3836
rect 10196 3834 10252 3836
rect 9956 3782 10002 3834
rect 10002 3782 10012 3834
rect 10036 3782 10066 3834
rect 10066 3782 10078 3834
rect 10078 3782 10092 3834
rect 10116 3782 10130 3834
rect 10130 3782 10142 3834
rect 10142 3782 10172 3834
rect 10196 3782 10206 3834
rect 10206 3782 10252 3834
rect 9956 3780 10012 3782
rect 10036 3780 10092 3782
rect 10116 3780 10172 3782
rect 10196 3780 10252 3782
rect 17956 3834 18012 3836
rect 18036 3834 18092 3836
rect 18116 3834 18172 3836
rect 18196 3834 18252 3836
rect 17956 3782 18002 3834
rect 18002 3782 18012 3834
rect 18036 3782 18066 3834
rect 18066 3782 18078 3834
rect 18078 3782 18092 3834
rect 18116 3782 18130 3834
rect 18130 3782 18142 3834
rect 18142 3782 18172 3834
rect 18196 3782 18206 3834
rect 18206 3782 18252 3834
rect 17956 3780 18012 3782
rect 18036 3780 18092 3782
rect 18116 3780 18172 3782
rect 18196 3780 18252 3782
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 10616 3290 10672 3292
rect 10696 3290 10752 3292
rect 10776 3290 10832 3292
rect 10856 3290 10912 3292
rect 10616 3238 10662 3290
rect 10662 3238 10672 3290
rect 10696 3238 10726 3290
rect 10726 3238 10738 3290
rect 10738 3238 10752 3290
rect 10776 3238 10790 3290
rect 10790 3238 10802 3290
rect 10802 3238 10832 3290
rect 10856 3238 10866 3290
rect 10866 3238 10912 3290
rect 10616 3236 10672 3238
rect 10696 3236 10752 3238
rect 10776 3236 10832 3238
rect 10856 3236 10912 3238
rect 18616 3290 18672 3292
rect 18696 3290 18752 3292
rect 18776 3290 18832 3292
rect 18856 3290 18912 3292
rect 18616 3238 18662 3290
rect 18662 3238 18672 3290
rect 18696 3238 18726 3290
rect 18726 3238 18738 3290
rect 18738 3238 18752 3290
rect 18776 3238 18790 3290
rect 18790 3238 18802 3290
rect 18802 3238 18832 3290
rect 18856 3238 18866 3290
rect 18866 3238 18912 3290
rect 18616 3236 18672 3238
rect 18696 3236 18752 3238
rect 18776 3236 18832 3238
rect 18856 3236 18912 3238
rect 26616 3290 26672 3292
rect 26696 3290 26752 3292
rect 26776 3290 26832 3292
rect 26856 3290 26912 3292
rect 26616 3238 26662 3290
rect 26662 3238 26672 3290
rect 26696 3238 26726 3290
rect 26726 3238 26738 3290
rect 26738 3238 26752 3290
rect 26776 3238 26790 3290
rect 26790 3238 26802 3290
rect 26802 3238 26832 3290
rect 26856 3238 26866 3290
rect 26866 3238 26912 3290
rect 26616 3236 26672 3238
rect 26696 3236 26752 3238
rect 26776 3236 26832 3238
rect 26856 3236 26912 3238
rect 28354 12280 28410 12336
rect 28354 10648 28410 10704
rect 28354 9016 28410 9072
rect 28354 7384 28410 7440
rect 28354 5752 28410 5808
rect 28354 4120 28410 4176
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 9956 2746 10012 2748
rect 10036 2746 10092 2748
rect 10116 2746 10172 2748
rect 10196 2746 10252 2748
rect 9956 2694 10002 2746
rect 10002 2694 10012 2746
rect 10036 2694 10066 2746
rect 10066 2694 10078 2746
rect 10078 2694 10092 2746
rect 10116 2694 10130 2746
rect 10130 2694 10142 2746
rect 10142 2694 10172 2746
rect 10196 2694 10206 2746
rect 10206 2694 10252 2746
rect 9956 2692 10012 2694
rect 10036 2692 10092 2694
rect 10116 2692 10172 2694
rect 10196 2692 10252 2694
rect 17956 2746 18012 2748
rect 18036 2746 18092 2748
rect 18116 2746 18172 2748
rect 18196 2746 18252 2748
rect 17956 2694 18002 2746
rect 18002 2694 18012 2746
rect 18036 2694 18066 2746
rect 18066 2694 18078 2746
rect 18078 2694 18092 2746
rect 18116 2694 18130 2746
rect 18130 2694 18142 2746
rect 18142 2694 18172 2746
rect 18196 2694 18206 2746
rect 18206 2694 18252 2746
rect 17956 2692 18012 2694
rect 18036 2692 18092 2694
rect 18116 2692 18172 2694
rect 18196 2692 18252 2694
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 28354 2488 28410 2544
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 10616 2202 10672 2204
rect 10696 2202 10752 2204
rect 10776 2202 10832 2204
rect 10856 2202 10912 2204
rect 10616 2150 10662 2202
rect 10662 2150 10672 2202
rect 10696 2150 10726 2202
rect 10726 2150 10738 2202
rect 10738 2150 10752 2202
rect 10776 2150 10790 2202
rect 10790 2150 10802 2202
rect 10802 2150 10832 2202
rect 10856 2150 10866 2202
rect 10866 2150 10912 2202
rect 10616 2148 10672 2150
rect 10696 2148 10752 2150
rect 10776 2148 10832 2150
rect 10856 2148 10912 2150
rect 18616 2202 18672 2204
rect 18696 2202 18752 2204
rect 18776 2202 18832 2204
rect 18856 2202 18912 2204
rect 18616 2150 18662 2202
rect 18662 2150 18672 2202
rect 18696 2150 18726 2202
rect 18726 2150 18738 2202
rect 18738 2150 18752 2202
rect 18776 2150 18790 2202
rect 18790 2150 18802 2202
rect 18802 2150 18832 2202
rect 18856 2150 18866 2202
rect 18866 2150 18912 2202
rect 18616 2148 18672 2150
rect 18696 2148 18752 2150
rect 18776 2148 18832 2150
rect 18856 2148 18912 2150
rect 26616 2202 26672 2204
rect 26696 2202 26752 2204
rect 26776 2202 26832 2204
rect 26856 2202 26912 2204
rect 26616 2150 26662 2202
rect 26662 2150 26672 2202
rect 26696 2150 26726 2202
rect 26726 2150 26738 2202
rect 26738 2150 26752 2202
rect 26776 2150 26790 2202
rect 26790 2150 26802 2202
rect 26802 2150 26832 2202
rect 26856 2150 26866 2202
rect 26866 2150 26912 2202
rect 26616 2148 26672 2150
rect 26696 2148 26752 2150
rect 26776 2148 26832 2150
rect 26856 2148 26912 2150
<< metal3 >>
rect 1946 27776 2262 27777
rect 1946 27712 1952 27776
rect 2016 27712 2032 27776
rect 2096 27712 2112 27776
rect 2176 27712 2192 27776
rect 2256 27712 2262 27776
rect 1946 27711 2262 27712
rect 9946 27776 10262 27777
rect 9946 27712 9952 27776
rect 10016 27712 10032 27776
rect 10096 27712 10112 27776
rect 10176 27712 10192 27776
rect 10256 27712 10262 27776
rect 9946 27711 10262 27712
rect 17946 27776 18262 27777
rect 17946 27712 17952 27776
rect 18016 27712 18032 27776
rect 18096 27712 18112 27776
rect 18176 27712 18192 27776
rect 18256 27712 18262 27776
rect 17946 27711 18262 27712
rect 25946 27776 26262 27777
rect 25946 27712 25952 27776
rect 26016 27712 26032 27776
rect 26096 27712 26112 27776
rect 26176 27712 26192 27776
rect 26256 27712 26262 27776
rect 25946 27711 26262 27712
rect 2606 27232 2922 27233
rect 2606 27168 2612 27232
rect 2676 27168 2692 27232
rect 2756 27168 2772 27232
rect 2836 27168 2852 27232
rect 2916 27168 2922 27232
rect 2606 27167 2922 27168
rect 10606 27232 10922 27233
rect 10606 27168 10612 27232
rect 10676 27168 10692 27232
rect 10756 27168 10772 27232
rect 10836 27168 10852 27232
rect 10916 27168 10922 27232
rect 10606 27167 10922 27168
rect 18606 27232 18922 27233
rect 18606 27168 18612 27232
rect 18676 27168 18692 27232
rect 18756 27168 18772 27232
rect 18836 27168 18852 27232
rect 18916 27168 18922 27232
rect 18606 27167 18922 27168
rect 26606 27232 26922 27233
rect 26606 27168 26612 27232
rect 26676 27168 26692 27232
rect 26756 27168 26772 27232
rect 26836 27168 26852 27232
rect 26916 27168 26922 27232
rect 26606 27167 26922 27168
rect 28349 27026 28415 27029
rect 29200 27026 30000 27056
rect 28349 27024 30000 27026
rect 28349 26968 28354 27024
rect 28410 26968 30000 27024
rect 28349 26966 30000 26968
rect 28349 26963 28415 26966
rect 29200 26936 30000 26966
rect 1946 26688 2262 26689
rect 1946 26624 1952 26688
rect 2016 26624 2032 26688
rect 2096 26624 2112 26688
rect 2176 26624 2192 26688
rect 2256 26624 2262 26688
rect 1946 26623 2262 26624
rect 9946 26688 10262 26689
rect 9946 26624 9952 26688
rect 10016 26624 10032 26688
rect 10096 26624 10112 26688
rect 10176 26624 10192 26688
rect 10256 26624 10262 26688
rect 9946 26623 10262 26624
rect 17946 26688 18262 26689
rect 17946 26624 17952 26688
rect 18016 26624 18032 26688
rect 18096 26624 18112 26688
rect 18176 26624 18192 26688
rect 18256 26624 18262 26688
rect 17946 26623 18262 26624
rect 25946 26688 26262 26689
rect 25946 26624 25952 26688
rect 26016 26624 26032 26688
rect 26096 26624 26112 26688
rect 26176 26624 26192 26688
rect 26256 26624 26262 26688
rect 25946 26623 26262 26624
rect 2606 26144 2922 26145
rect 2606 26080 2612 26144
rect 2676 26080 2692 26144
rect 2756 26080 2772 26144
rect 2836 26080 2852 26144
rect 2916 26080 2922 26144
rect 2606 26079 2922 26080
rect 10606 26144 10922 26145
rect 10606 26080 10612 26144
rect 10676 26080 10692 26144
rect 10756 26080 10772 26144
rect 10836 26080 10852 26144
rect 10916 26080 10922 26144
rect 10606 26079 10922 26080
rect 18606 26144 18922 26145
rect 18606 26080 18612 26144
rect 18676 26080 18692 26144
rect 18756 26080 18772 26144
rect 18836 26080 18852 26144
rect 18916 26080 18922 26144
rect 18606 26079 18922 26080
rect 26606 26144 26922 26145
rect 26606 26080 26612 26144
rect 26676 26080 26692 26144
rect 26756 26080 26772 26144
rect 26836 26080 26852 26144
rect 26916 26080 26922 26144
rect 26606 26079 26922 26080
rect 1946 25600 2262 25601
rect 1946 25536 1952 25600
rect 2016 25536 2032 25600
rect 2096 25536 2112 25600
rect 2176 25536 2192 25600
rect 2256 25536 2262 25600
rect 1946 25535 2262 25536
rect 9946 25600 10262 25601
rect 9946 25536 9952 25600
rect 10016 25536 10032 25600
rect 10096 25536 10112 25600
rect 10176 25536 10192 25600
rect 10256 25536 10262 25600
rect 9946 25535 10262 25536
rect 17946 25600 18262 25601
rect 17946 25536 17952 25600
rect 18016 25536 18032 25600
rect 18096 25536 18112 25600
rect 18176 25536 18192 25600
rect 18256 25536 18262 25600
rect 17946 25535 18262 25536
rect 25946 25600 26262 25601
rect 25946 25536 25952 25600
rect 26016 25536 26032 25600
rect 26096 25536 26112 25600
rect 26176 25536 26192 25600
rect 26256 25536 26262 25600
rect 25946 25535 26262 25536
rect 28349 25394 28415 25397
rect 29200 25394 30000 25424
rect 28349 25392 30000 25394
rect 28349 25336 28354 25392
rect 28410 25336 30000 25392
rect 28349 25334 30000 25336
rect 28349 25331 28415 25334
rect 29200 25304 30000 25334
rect 2606 25056 2922 25057
rect 2606 24992 2612 25056
rect 2676 24992 2692 25056
rect 2756 24992 2772 25056
rect 2836 24992 2852 25056
rect 2916 24992 2922 25056
rect 2606 24991 2922 24992
rect 10606 25056 10922 25057
rect 10606 24992 10612 25056
rect 10676 24992 10692 25056
rect 10756 24992 10772 25056
rect 10836 24992 10852 25056
rect 10916 24992 10922 25056
rect 10606 24991 10922 24992
rect 18606 25056 18922 25057
rect 18606 24992 18612 25056
rect 18676 24992 18692 25056
rect 18756 24992 18772 25056
rect 18836 24992 18852 25056
rect 18916 24992 18922 25056
rect 18606 24991 18922 24992
rect 26606 25056 26922 25057
rect 26606 24992 26612 25056
rect 26676 24992 26692 25056
rect 26756 24992 26772 25056
rect 26836 24992 26852 25056
rect 26916 24992 26922 25056
rect 26606 24991 26922 24992
rect 1946 24512 2262 24513
rect 1946 24448 1952 24512
rect 2016 24448 2032 24512
rect 2096 24448 2112 24512
rect 2176 24448 2192 24512
rect 2256 24448 2262 24512
rect 1946 24447 2262 24448
rect 9946 24512 10262 24513
rect 9946 24448 9952 24512
rect 10016 24448 10032 24512
rect 10096 24448 10112 24512
rect 10176 24448 10192 24512
rect 10256 24448 10262 24512
rect 9946 24447 10262 24448
rect 17946 24512 18262 24513
rect 17946 24448 17952 24512
rect 18016 24448 18032 24512
rect 18096 24448 18112 24512
rect 18176 24448 18192 24512
rect 18256 24448 18262 24512
rect 17946 24447 18262 24448
rect 25946 24512 26262 24513
rect 25946 24448 25952 24512
rect 26016 24448 26032 24512
rect 26096 24448 26112 24512
rect 26176 24448 26192 24512
rect 26256 24448 26262 24512
rect 25946 24447 26262 24448
rect 2606 23968 2922 23969
rect 2606 23904 2612 23968
rect 2676 23904 2692 23968
rect 2756 23904 2772 23968
rect 2836 23904 2852 23968
rect 2916 23904 2922 23968
rect 2606 23903 2922 23904
rect 10606 23968 10922 23969
rect 10606 23904 10612 23968
rect 10676 23904 10692 23968
rect 10756 23904 10772 23968
rect 10836 23904 10852 23968
rect 10916 23904 10922 23968
rect 10606 23903 10922 23904
rect 18606 23968 18922 23969
rect 18606 23904 18612 23968
rect 18676 23904 18692 23968
rect 18756 23904 18772 23968
rect 18836 23904 18852 23968
rect 18916 23904 18922 23968
rect 18606 23903 18922 23904
rect 26606 23968 26922 23969
rect 26606 23904 26612 23968
rect 26676 23904 26692 23968
rect 26756 23904 26772 23968
rect 26836 23904 26852 23968
rect 26916 23904 26922 23968
rect 26606 23903 26922 23904
rect 28349 23762 28415 23765
rect 29200 23762 30000 23792
rect 28349 23760 30000 23762
rect 28349 23704 28354 23760
rect 28410 23704 30000 23760
rect 28349 23702 30000 23704
rect 28349 23699 28415 23702
rect 29200 23672 30000 23702
rect 1946 23424 2262 23425
rect 1946 23360 1952 23424
rect 2016 23360 2032 23424
rect 2096 23360 2112 23424
rect 2176 23360 2192 23424
rect 2256 23360 2262 23424
rect 1946 23359 2262 23360
rect 9946 23424 10262 23425
rect 9946 23360 9952 23424
rect 10016 23360 10032 23424
rect 10096 23360 10112 23424
rect 10176 23360 10192 23424
rect 10256 23360 10262 23424
rect 9946 23359 10262 23360
rect 17946 23424 18262 23425
rect 17946 23360 17952 23424
rect 18016 23360 18032 23424
rect 18096 23360 18112 23424
rect 18176 23360 18192 23424
rect 18256 23360 18262 23424
rect 17946 23359 18262 23360
rect 25946 23424 26262 23425
rect 25946 23360 25952 23424
rect 26016 23360 26032 23424
rect 26096 23360 26112 23424
rect 26176 23360 26192 23424
rect 26256 23360 26262 23424
rect 25946 23359 26262 23360
rect 2606 22880 2922 22881
rect 2606 22816 2612 22880
rect 2676 22816 2692 22880
rect 2756 22816 2772 22880
rect 2836 22816 2852 22880
rect 2916 22816 2922 22880
rect 2606 22815 2922 22816
rect 10606 22880 10922 22881
rect 10606 22816 10612 22880
rect 10676 22816 10692 22880
rect 10756 22816 10772 22880
rect 10836 22816 10852 22880
rect 10916 22816 10922 22880
rect 10606 22815 10922 22816
rect 18606 22880 18922 22881
rect 18606 22816 18612 22880
rect 18676 22816 18692 22880
rect 18756 22816 18772 22880
rect 18836 22816 18852 22880
rect 18916 22816 18922 22880
rect 18606 22815 18922 22816
rect 26606 22880 26922 22881
rect 26606 22816 26612 22880
rect 26676 22816 26692 22880
rect 26756 22816 26772 22880
rect 26836 22816 26852 22880
rect 26916 22816 26922 22880
rect 26606 22815 26922 22816
rect 841 22538 907 22541
rect 798 22536 907 22538
rect 798 22480 846 22536
rect 902 22480 907 22536
rect 798 22475 907 22480
rect 798 22432 858 22475
rect 0 22342 858 22432
rect 0 22312 800 22342
rect 1946 22336 2262 22337
rect 1946 22272 1952 22336
rect 2016 22272 2032 22336
rect 2096 22272 2112 22336
rect 2176 22272 2192 22336
rect 2256 22272 2262 22336
rect 1946 22271 2262 22272
rect 9946 22336 10262 22337
rect 9946 22272 9952 22336
rect 10016 22272 10032 22336
rect 10096 22272 10112 22336
rect 10176 22272 10192 22336
rect 10256 22272 10262 22336
rect 9946 22271 10262 22272
rect 17946 22336 18262 22337
rect 17946 22272 17952 22336
rect 18016 22272 18032 22336
rect 18096 22272 18112 22336
rect 18176 22272 18192 22336
rect 18256 22272 18262 22336
rect 17946 22271 18262 22272
rect 25946 22336 26262 22337
rect 25946 22272 25952 22336
rect 26016 22272 26032 22336
rect 26096 22272 26112 22336
rect 26176 22272 26192 22336
rect 26256 22272 26262 22336
rect 25946 22271 26262 22272
rect 28349 22130 28415 22133
rect 29200 22130 30000 22160
rect 28349 22128 30000 22130
rect 28349 22072 28354 22128
rect 28410 22072 30000 22128
rect 28349 22070 30000 22072
rect 28349 22067 28415 22070
rect 29200 22040 30000 22070
rect 2606 21792 2922 21793
rect 2606 21728 2612 21792
rect 2676 21728 2692 21792
rect 2756 21728 2772 21792
rect 2836 21728 2852 21792
rect 2916 21728 2922 21792
rect 2606 21727 2922 21728
rect 10606 21792 10922 21793
rect 10606 21728 10612 21792
rect 10676 21728 10692 21792
rect 10756 21728 10772 21792
rect 10836 21728 10852 21792
rect 10916 21728 10922 21792
rect 10606 21727 10922 21728
rect 18606 21792 18922 21793
rect 18606 21728 18612 21792
rect 18676 21728 18692 21792
rect 18756 21728 18772 21792
rect 18836 21728 18852 21792
rect 18916 21728 18922 21792
rect 18606 21727 18922 21728
rect 26606 21792 26922 21793
rect 26606 21728 26612 21792
rect 26676 21728 26692 21792
rect 26756 21728 26772 21792
rect 26836 21728 26852 21792
rect 26916 21728 26922 21792
rect 26606 21727 26922 21728
rect 1946 21248 2262 21249
rect 1946 21184 1952 21248
rect 2016 21184 2032 21248
rect 2096 21184 2112 21248
rect 2176 21184 2192 21248
rect 2256 21184 2262 21248
rect 1946 21183 2262 21184
rect 9946 21248 10262 21249
rect 9946 21184 9952 21248
rect 10016 21184 10032 21248
rect 10096 21184 10112 21248
rect 10176 21184 10192 21248
rect 10256 21184 10262 21248
rect 9946 21183 10262 21184
rect 17946 21248 18262 21249
rect 17946 21184 17952 21248
rect 18016 21184 18032 21248
rect 18096 21184 18112 21248
rect 18176 21184 18192 21248
rect 18256 21184 18262 21248
rect 17946 21183 18262 21184
rect 25946 21248 26262 21249
rect 25946 21184 25952 21248
rect 26016 21184 26032 21248
rect 26096 21184 26112 21248
rect 26176 21184 26192 21248
rect 26256 21184 26262 21248
rect 25946 21183 26262 21184
rect 2606 20704 2922 20705
rect 2606 20640 2612 20704
rect 2676 20640 2692 20704
rect 2756 20640 2772 20704
rect 2836 20640 2852 20704
rect 2916 20640 2922 20704
rect 2606 20639 2922 20640
rect 10606 20704 10922 20705
rect 10606 20640 10612 20704
rect 10676 20640 10692 20704
rect 10756 20640 10772 20704
rect 10836 20640 10852 20704
rect 10916 20640 10922 20704
rect 10606 20639 10922 20640
rect 18606 20704 18922 20705
rect 18606 20640 18612 20704
rect 18676 20640 18692 20704
rect 18756 20640 18772 20704
rect 18836 20640 18852 20704
rect 18916 20640 18922 20704
rect 18606 20639 18922 20640
rect 26606 20704 26922 20705
rect 26606 20640 26612 20704
rect 26676 20640 26692 20704
rect 26756 20640 26772 20704
rect 26836 20640 26852 20704
rect 26916 20640 26922 20704
rect 26606 20639 26922 20640
rect 28349 20498 28415 20501
rect 29200 20498 30000 20528
rect 28349 20496 30000 20498
rect 28349 20440 28354 20496
rect 28410 20440 30000 20496
rect 28349 20438 30000 20440
rect 28349 20435 28415 20438
rect 29200 20408 30000 20438
rect 1946 20160 2262 20161
rect 1946 20096 1952 20160
rect 2016 20096 2032 20160
rect 2096 20096 2112 20160
rect 2176 20096 2192 20160
rect 2256 20096 2262 20160
rect 1946 20095 2262 20096
rect 9946 20160 10262 20161
rect 9946 20096 9952 20160
rect 10016 20096 10032 20160
rect 10096 20096 10112 20160
rect 10176 20096 10192 20160
rect 10256 20096 10262 20160
rect 9946 20095 10262 20096
rect 17946 20160 18262 20161
rect 17946 20096 17952 20160
rect 18016 20096 18032 20160
rect 18096 20096 18112 20160
rect 18176 20096 18192 20160
rect 18256 20096 18262 20160
rect 17946 20095 18262 20096
rect 25946 20160 26262 20161
rect 25946 20096 25952 20160
rect 26016 20096 26032 20160
rect 26096 20096 26112 20160
rect 26176 20096 26192 20160
rect 26256 20096 26262 20160
rect 25946 20095 26262 20096
rect 2606 19616 2922 19617
rect 2606 19552 2612 19616
rect 2676 19552 2692 19616
rect 2756 19552 2772 19616
rect 2836 19552 2852 19616
rect 2916 19552 2922 19616
rect 2606 19551 2922 19552
rect 10606 19616 10922 19617
rect 10606 19552 10612 19616
rect 10676 19552 10692 19616
rect 10756 19552 10772 19616
rect 10836 19552 10852 19616
rect 10916 19552 10922 19616
rect 10606 19551 10922 19552
rect 18606 19616 18922 19617
rect 18606 19552 18612 19616
rect 18676 19552 18692 19616
rect 18756 19552 18772 19616
rect 18836 19552 18852 19616
rect 18916 19552 18922 19616
rect 18606 19551 18922 19552
rect 26606 19616 26922 19617
rect 26606 19552 26612 19616
rect 26676 19552 26692 19616
rect 26756 19552 26772 19616
rect 26836 19552 26852 19616
rect 26916 19552 26922 19616
rect 26606 19551 26922 19552
rect 1946 19072 2262 19073
rect 1946 19008 1952 19072
rect 2016 19008 2032 19072
rect 2096 19008 2112 19072
rect 2176 19008 2192 19072
rect 2256 19008 2262 19072
rect 1946 19007 2262 19008
rect 9946 19072 10262 19073
rect 9946 19008 9952 19072
rect 10016 19008 10032 19072
rect 10096 19008 10112 19072
rect 10176 19008 10192 19072
rect 10256 19008 10262 19072
rect 9946 19007 10262 19008
rect 17946 19072 18262 19073
rect 17946 19008 17952 19072
rect 18016 19008 18032 19072
rect 18096 19008 18112 19072
rect 18176 19008 18192 19072
rect 18256 19008 18262 19072
rect 17946 19007 18262 19008
rect 25946 19072 26262 19073
rect 25946 19008 25952 19072
rect 26016 19008 26032 19072
rect 26096 19008 26112 19072
rect 26176 19008 26192 19072
rect 26256 19008 26262 19072
rect 25946 19007 26262 19008
rect 28349 18866 28415 18869
rect 29200 18866 30000 18896
rect 28349 18864 30000 18866
rect 28349 18808 28354 18864
rect 28410 18808 30000 18864
rect 28349 18806 30000 18808
rect 28349 18803 28415 18806
rect 29200 18776 30000 18806
rect 2606 18528 2922 18529
rect 2606 18464 2612 18528
rect 2676 18464 2692 18528
rect 2756 18464 2772 18528
rect 2836 18464 2852 18528
rect 2916 18464 2922 18528
rect 2606 18463 2922 18464
rect 10606 18528 10922 18529
rect 10606 18464 10612 18528
rect 10676 18464 10692 18528
rect 10756 18464 10772 18528
rect 10836 18464 10852 18528
rect 10916 18464 10922 18528
rect 10606 18463 10922 18464
rect 18606 18528 18922 18529
rect 18606 18464 18612 18528
rect 18676 18464 18692 18528
rect 18756 18464 18772 18528
rect 18836 18464 18852 18528
rect 18916 18464 18922 18528
rect 18606 18463 18922 18464
rect 26606 18528 26922 18529
rect 26606 18464 26612 18528
rect 26676 18464 26692 18528
rect 26756 18464 26772 18528
rect 26836 18464 26852 18528
rect 26916 18464 26922 18528
rect 26606 18463 26922 18464
rect 1946 17984 2262 17985
rect 1946 17920 1952 17984
rect 2016 17920 2032 17984
rect 2096 17920 2112 17984
rect 2176 17920 2192 17984
rect 2256 17920 2262 17984
rect 1946 17919 2262 17920
rect 9946 17984 10262 17985
rect 9946 17920 9952 17984
rect 10016 17920 10032 17984
rect 10096 17920 10112 17984
rect 10176 17920 10192 17984
rect 10256 17920 10262 17984
rect 9946 17919 10262 17920
rect 17946 17984 18262 17985
rect 17946 17920 17952 17984
rect 18016 17920 18032 17984
rect 18096 17920 18112 17984
rect 18176 17920 18192 17984
rect 18256 17920 18262 17984
rect 17946 17919 18262 17920
rect 25946 17984 26262 17985
rect 25946 17920 25952 17984
rect 26016 17920 26032 17984
rect 26096 17920 26112 17984
rect 26176 17920 26192 17984
rect 26256 17920 26262 17984
rect 25946 17919 26262 17920
rect 2606 17440 2922 17441
rect 2606 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2922 17440
rect 2606 17375 2922 17376
rect 10606 17440 10922 17441
rect 10606 17376 10612 17440
rect 10676 17376 10692 17440
rect 10756 17376 10772 17440
rect 10836 17376 10852 17440
rect 10916 17376 10922 17440
rect 10606 17375 10922 17376
rect 18606 17440 18922 17441
rect 18606 17376 18612 17440
rect 18676 17376 18692 17440
rect 18756 17376 18772 17440
rect 18836 17376 18852 17440
rect 18916 17376 18922 17440
rect 18606 17375 18922 17376
rect 26606 17440 26922 17441
rect 26606 17376 26612 17440
rect 26676 17376 26692 17440
rect 26756 17376 26772 17440
rect 26836 17376 26852 17440
rect 26916 17376 26922 17440
rect 26606 17375 26922 17376
rect 28349 17234 28415 17237
rect 29200 17234 30000 17264
rect 28349 17232 30000 17234
rect 28349 17176 28354 17232
rect 28410 17176 30000 17232
rect 28349 17174 30000 17176
rect 28349 17171 28415 17174
rect 29200 17144 30000 17174
rect 1946 16896 2262 16897
rect 1946 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2262 16896
rect 1946 16831 2262 16832
rect 9946 16896 10262 16897
rect 9946 16832 9952 16896
rect 10016 16832 10032 16896
rect 10096 16832 10112 16896
rect 10176 16832 10192 16896
rect 10256 16832 10262 16896
rect 9946 16831 10262 16832
rect 17946 16896 18262 16897
rect 17946 16832 17952 16896
rect 18016 16832 18032 16896
rect 18096 16832 18112 16896
rect 18176 16832 18192 16896
rect 18256 16832 18262 16896
rect 17946 16831 18262 16832
rect 25946 16896 26262 16897
rect 25946 16832 25952 16896
rect 26016 16832 26032 16896
rect 26096 16832 26112 16896
rect 26176 16832 26192 16896
rect 26256 16832 26262 16896
rect 25946 16831 26262 16832
rect 2606 16352 2922 16353
rect 2606 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2922 16352
rect 2606 16287 2922 16288
rect 10606 16352 10922 16353
rect 10606 16288 10612 16352
rect 10676 16288 10692 16352
rect 10756 16288 10772 16352
rect 10836 16288 10852 16352
rect 10916 16288 10922 16352
rect 10606 16287 10922 16288
rect 18606 16352 18922 16353
rect 18606 16288 18612 16352
rect 18676 16288 18692 16352
rect 18756 16288 18772 16352
rect 18836 16288 18852 16352
rect 18916 16288 18922 16352
rect 18606 16287 18922 16288
rect 26606 16352 26922 16353
rect 26606 16288 26612 16352
rect 26676 16288 26692 16352
rect 26756 16288 26772 16352
rect 26836 16288 26852 16352
rect 26916 16288 26922 16352
rect 26606 16287 26922 16288
rect 1946 15808 2262 15809
rect 1946 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2262 15808
rect 1946 15743 2262 15744
rect 9946 15808 10262 15809
rect 9946 15744 9952 15808
rect 10016 15744 10032 15808
rect 10096 15744 10112 15808
rect 10176 15744 10192 15808
rect 10256 15744 10262 15808
rect 9946 15743 10262 15744
rect 17946 15808 18262 15809
rect 17946 15744 17952 15808
rect 18016 15744 18032 15808
rect 18096 15744 18112 15808
rect 18176 15744 18192 15808
rect 18256 15744 18262 15808
rect 17946 15743 18262 15744
rect 25946 15808 26262 15809
rect 25946 15744 25952 15808
rect 26016 15744 26032 15808
rect 26096 15744 26112 15808
rect 26176 15744 26192 15808
rect 26256 15744 26262 15808
rect 25946 15743 26262 15744
rect 28349 15602 28415 15605
rect 29200 15602 30000 15632
rect 28349 15600 30000 15602
rect 28349 15544 28354 15600
rect 28410 15544 30000 15600
rect 28349 15542 30000 15544
rect 28349 15539 28415 15542
rect 29200 15512 30000 15542
rect 2606 15264 2922 15265
rect 2606 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2922 15264
rect 2606 15199 2922 15200
rect 10606 15264 10922 15265
rect 10606 15200 10612 15264
rect 10676 15200 10692 15264
rect 10756 15200 10772 15264
rect 10836 15200 10852 15264
rect 10916 15200 10922 15264
rect 10606 15199 10922 15200
rect 18606 15264 18922 15265
rect 18606 15200 18612 15264
rect 18676 15200 18692 15264
rect 18756 15200 18772 15264
rect 18836 15200 18852 15264
rect 18916 15200 18922 15264
rect 18606 15199 18922 15200
rect 26606 15264 26922 15265
rect 26606 15200 26612 15264
rect 26676 15200 26692 15264
rect 26756 15200 26772 15264
rect 26836 15200 26852 15264
rect 26916 15200 26922 15264
rect 26606 15199 26922 15200
rect 1946 14720 2262 14721
rect 1946 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2262 14720
rect 1946 14655 2262 14656
rect 9946 14720 10262 14721
rect 9946 14656 9952 14720
rect 10016 14656 10032 14720
rect 10096 14656 10112 14720
rect 10176 14656 10192 14720
rect 10256 14656 10262 14720
rect 9946 14655 10262 14656
rect 17946 14720 18262 14721
rect 17946 14656 17952 14720
rect 18016 14656 18032 14720
rect 18096 14656 18112 14720
rect 18176 14656 18192 14720
rect 18256 14656 18262 14720
rect 17946 14655 18262 14656
rect 25946 14720 26262 14721
rect 25946 14656 25952 14720
rect 26016 14656 26032 14720
rect 26096 14656 26112 14720
rect 26176 14656 26192 14720
rect 26256 14656 26262 14720
rect 25946 14655 26262 14656
rect 2606 14176 2922 14177
rect 2606 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2922 14176
rect 2606 14111 2922 14112
rect 10606 14176 10922 14177
rect 10606 14112 10612 14176
rect 10676 14112 10692 14176
rect 10756 14112 10772 14176
rect 10836 14112 10852 14176
rect 10916 14112 10922 14176
rect 10606 14111 10922 14112
rect 18606 14176 18922 14177
rect 18606 14112 18612 14176
rect 18676 14112 18692 14176
rect 18756 14112 18772 14176
rect 18836 14112 18852 14176
rect 18916 14112 18922 14176
rect 18606 14111 18922 14112
rect 26606 14176 26922 14177
rect 26606 14112 26612 14176
rect 26676 14112 26692 14176
rect 26756 14112 26772 14176
rect 26836 14112 26852 14176
rect 26916 14112 26922 14176
rect 26606 14111 26922 14112
rect 28349 13970 28415 13973
rect 29200 13970 30000 14000
rect 28349 13968 30000 13970
rect 28349 13912 28354 13968
rect 28410 13912 30000 13968
rect 28349 13910 30000 13912
rect 28349 13907 28415 13910
rect 29200 13880 30000 13910
rect 1946 13632 2262 13633
rect 1946 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2262 13632
rect 1946 13567 2262 13568
rect 9946 13632 10262 13633
rect 9946 13568 9952 13632
rect 10016 13568 10032 13632
rect 10096 13568 10112 13632
rect 10176 13568 10192 13632
rect 10256 13568 10262 13632
rect 9946 13567 10262 13568
rect 17946 13632 18262 13633
rect 17946 13568 17952 13632
rect 18016 13568 18032 13632
rect 18096 13568 18112 13632
rect 18176 13568 18192 13632
rect 18256 13568 18262 13632
rect 17946 13567 18262 13568
rect 25946 13632 26262 13633
rect 25946 13568 25952 13632
rect 26016 13568 26032 13632
rect 26096 13568 26112 13632
rect 26176 13568 26192 13632
rect 26256 13568 26262 13632
rect 25946 13567 26262 13568
rect 2606 13088 2922 13089
rect 2606 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2922 13088
rect 2606 13023 2922 13024
rect 10606 13088 10922 13089
rect 10606 13024 10612 13088
rect 10676 13024 10692 13088
rect 10756 13024 10772 13088
rect 10836 13024 10852 13088
rect 10916 13024 10922 13088
rect 10606 13023 10922 13024
rect 18606 13088 18922 13089
rect 18606 13024 18612 13088
rect 18676 13024 18692 13088
rect 18756 13024 18772 13088
rect 18836 13024 18852 13088
rect 18916 13024 18922 13088
rect 18606 13023 18922 13024
rect 26606 13088 26922 13089
rect 26606 13024 26612 13088
rect 26676 13024 26692 13088
rect 26756 13024 26772 13088
rect 26836 13024 26852 13088
rect 26916 13024 26922 13088
rect 26606 13023 26922 13024
rect 1946 12544 2262 12545
rect 1946 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2262 12544
rect 1946 12479 2262 12480
rect 9946 12544 10262 12545
rect 9946 12480 9952 12544
rect 10016 12480 10032 12544
rect 10096 12480 10112 12544
rect 10176 12480 10192 12544
rect 10256 12480 10262 12544
rect 9946 12479 10262 12480
rect 17946 12544 18262 12545
rect 17946 12480 17952 12544
rect 18016 12480 18032 12544
rect 18096 12480 18112 12544
rect 18176 12480 18192 12544
rect 18256 12480 18262 12544
rect 17946 12479 18262 12480
rect 25946 12544 26262 12545
rect 25946 12480 25952 12544
rect 26016 12480 26032 12544
rect 26096 12480 26112 12544
rect 26176 12480 26192 12544
rect 26256 12480 26262 12544
rect 25946 12479 26262 12480
rect 28349 12338 28415 12341
rect 29200 12338 30000 12368
rect 28349 12336 30000 12338
rect 28349 12280 28354 12336
rect 28410 12280 30000 12336
rect 28349 12278 30000 12280
rect 28349 12275 28415 12278
rect 29200 12248 30000 12278
rect 2606 12000 2922 12001
rect 2606 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2922 12000
rect 2606 11935 2922 11936
rect 10606 12000 10922 12001
rect 10606 11936 10612 12000
rect 10676 11936 10692 12000
rect 10756 11936 10772 12000
rect 10836 11936 10852 12000
rect 10916 11936 10922 12000
rect 10606 11935 10922 11936
rect 18606 12000 18922 12001
rect 18606 11936 18612 12000
rect 18676 11936 18692 12000
rect 18756 11936 18772 12000
rect 18836 11936 18852 12000
rect 18916 11936 18922 12000
rect 18606 11935 18922 11936
rect 26606 12000 26922 12001
rect 26606 11936 26612 12000
rect 26676 11936 26692 12000
rect 26756 11936 26772 12000
rect 26836 11936 26852 12000
rect 26916 11936 26922 12000
rect 26606 11935 26922 11936
rect 1946 11456 2262 11457
rect 1946 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2262 11456
rect 1946 11391 2262 11392
rect 9946 11456 10262 11457
rect 9946 11392 9952 11456
rect 10016 11392 10032 11456
rect 10096 11392 10112 11456
rect 10176 11392 10192 11456
rect 10256 11392 10262 11456
rect 9946 11391 10262 11392
rect 17946 11456 18262 11457
rect 17946 11392 17952 11456
rect 18016 11392 18032 11456
rect 18096 11392 18112 11456
rect 18176 11392 18192 11456
rect 18256 11392 18262 11456
rect 17946 11391 18262 11392
rect 25946 11456 26262 11457
rect 25946 11392 25952 11456
rect 26016 11392 26032 11456
rect 26096 11392 26112 11456
rect 26176 11392 26192 11456
rect 26256 11392 26262 11456
rect 25946 11391 26262 11392
rect 2606 10912 2922 10913
rect 2606 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2922 10912
rect 2606 10847 2922 10848
rect 10606 10912 10922 10913
rect 10606 10848 10612 10912
rect 10676 10848 10692 10912
rect 10756 10848 10772 10912
rect 10836 10848 10852 10912
rect 10916 10848 10922 10912
rect 10606 10847 10922 10848
rect 18606 10912 18922 10913
rect 18606 10848 18612 10912
rect 18676 10848 18692 10912
rect 18756 10848 18772 10912
rect 18836 10848 18852 10912
rect 18916 10848 18922 10912
rect 18606 10847 18922 10848
rect 26606 10912 26922 10913
rect 26606 10848 26612 10912
rect 26676 10848 26692 10912
rect 26756 10848 26772 10912
rect 26836 10848 26852 10912
rect 26916 10848 26922 10912
rect 26606 10847 26922 10848
rect 28349 10706 28415 10709
rect 29200 10706 30000 10736
rect 28349 10704 30000 10706
rect 28349 10648 28354 10704
rect 28410 10648 30000 10704
rect 28349 10646 30000 10648
rect 28349 10643 28415 10646
rect 29200 10616 30000 10646
rect 1946 10368 2262 10369
rect 1946 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2262 10368
rect 1946 10303 2262 10304
rect 9946 10368 10262 10369
rect 9946 10304 9952 10368
rect 10016 10304 10032 10368
rect 10096 10304 10112 10368
rect 10176 10304 10192 10368
rect 10256 10304 10262 10368
rect 9946 10303 10262 10304
rect 17946 10368 18262 10369
rect 17946 10304 17952 10368
rect 18016 10304 18032 10368
rect 18096 10304 18112 10368
rect 18176 10304 18192 10368
rect 18256 10304 18262 10368
rect 17946 10303 18262 10304
rect 25946 10368 26262 10369
rect 25946 10304 25952 10368
rect 26016 10304 26032 10368
rect 26096 10304 26112 10368
rect 26176 10304 26192 10368
rect 26256 10304 26262 10368
rect 25946 10303 26262 10304
rect 2606 9824 2922 9825
rect 2606 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2922 9824
rect 2606 9759 2922 9760
rect 10606 9824 10922 9825
rect 10606 9760 10612 9824
rect 10676 9760 10692 9824
rect 10756 9760 10772 9824
rect 10836 9760 10852 9824
rect 10916 9760 10922 9824
rect 10606 9759 10922 9760
rect 18606 9824 18922 9825
rect 18606 9760 18612 9824
rect 18676 9760 18692 9824
rect 18756 9760 18772 9824
rect 18836 9760 18852 9824
rect 18916 9760 18922 9824
rect 18606 9759 18922 9760
rect 26606 9824 26922 9825
rect 26606 9760 26612 9824
rect 26676 9760 26692 9824
rect 26756 9760 26772 9824
rect 26836 9760 26852 9824
rect 26916 9760 26922 9824
rect 26606 9759 26922 9760
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 9946 9280 10262 9281
rect 9946 9216 9952 9280
rect 10016 9216 10032 9280
rect 10096 9216 10112 9280
rect 10176 9216 10192 9280
rect 10256 9216 10262 9280
rect 9946 9215 10262 9216
rect 17946 9280 18262 9281
rect 17946 9216 17952 9280
rect 18016 9216 18032 9280
rect 18096 9216 18112 9280
rect 18176 9216 18192 9280
rect 18256 9216 18262 9280
rect 17946 9215 18262 9216
rect 25946 9280 26262 9281
rect 25946 9216 25952 9280
rect 26016 9216 26032 9280
rect 26096 9216 26112 9280
rect 26176 9216 26192 9280
rect 26256 9216 26262 9280
rect 25946 9215 26262 9216
rect 28349 9074 28415 9077
rect 29200 9074 30000 9104
rect 28349 9072 30000 9074
rect 28349 9016 28354 9072
rect 28410 9016 30000 9072
rect 28349 9014 30000 9016
rect 28349 9011 28415 9014
rect 29200 8984 30000 9014
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 10606 8736 10922 8737
rect 10606 8672 10612 8736
rect 10676 8672 10692 8736
rect 10756 8672 10772 8736
rect 10836 8672 10852 8736
rect 10916 8672 10922 8736
rect 10606 8671 10922 8672
rect 18606 8736 18922 8737
rect 18606 8672 18612 8736
rect 18676 8672 18692 8736
rect 18756 8672 18772 8736
rect 18836 8672 18852 8736
rect 18916 8672 18922 8736
rect 18606 8671 18922 8672
rect 26606 8736 26922 8737
rect 26606 8672 26612 8736
rect 26676 8672 26692 8736
rect 26756 8672 26772 8736
rect 26836 8672 26852 8736
rect 26916 8672 26922 8736
rect 26606 8671 26922 8672
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 9946 8192 10262 8193
rect 9946 8128 9952 8192
rect 10016 8128 10032 8192
rect 10096 8128 10112 8192
rect 10176 8128 10192 8192
rect 10256 8128 10262 8192
rect 9946 8127 10262 8128
rect 17946 8192 18262 8193
rect 17946 8128 17952 8192
rect 18016 8128 18032 8192
rect 18096 8128 18112 8192
rect 18176 8128 18192 8192
rect 18256 8128 18262 8192
rect 17946 8127 18262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 10606 7648 10922 7649
rect 10606 7584 10612 7648
rect 10676 7584 10692 7648
rect 10756 7584 10772 7648
rect 10836 7584 10852 7648
rect 10916 7584 10922 7648
rect 10606 7583 10922 7584
rect 18606 7648 18922 7649
rect 18606 7584 18612 7648
rect 18676 7584 18692 7648
rect 18756 7584 18772 7648
rect 18836 7584 18852 7648
rect 18916 7584 18922 7648
rect 18606 7583 18922 7584
rect 26606 7648 26922 7649
rect 26606 7584 26612 7648
rect 26676 7584 26692 7648
rect 26756 7584 26772 7648
rect 26836 7584 26852 7648
rect 26916 7584 26922 7648
rect 26606 7583 26922 7584
rect 841 7578 907 7581
rect 798 7576 907 7578
rect 798 7520 846 7576
rect 902 7520 907 7576
rect 798 7515 907 7520
rect 798 7472 858 7515
rect 0 7382 858 7472
rect 28349 7442 28415 7445
rect 29200 7442 30000 7472
rect 28349 7440 30000 7442
rect 28349 7384 28354 7440
rect 28410 7384 30000 7440
rect 28349 7382 30000 7384
rect 0 7352 800 7382
rect 28349 7379 28415 7382
rect 29200 7352 30000 7382
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 9946 7104 10262 7105
rect 9946 7040 9952 7104
rect 10016 7040 10032 7104
rect 10096 7040 10112 7104
rect 10176 7040 10192 7104
rect 10256 7040 10262 7104
rect 9946 7039 10262 7040
rect 17946 7104 18262 7105
rect 17946 7040 17952 7104
rect 18016 7040 18032 7104
rect 18096 7040 18112 7104
rect 18176 7040 18192 7104
rect 18256 7040 18262 7104
rect 17946 7039 18262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 10606 6560 10922 6561
rect 10606 6496 10612 6560
rect 10676 6496 10692 6560
rect 10756 6496 10772 6560
rect 10836 6496 10852 6560
rect 10916 6496 10922 6560
rect 10606 6495 10922 6496
rect 18606 6560 18922 6561
rect 18606 6496 18612 6560
rect 18676 6496 18692 6560
rect 18756 6496 18772 6560
rect 18836 6496 18852 6560
rect 18916 6496 18922 6560
rect 18606 6495 18922 6496
rect 26606 6560 26922 6561
rect 26606 6496 26612 6560
rect 26676 6496 26692 6560
rect 26756 6496 26772 6560
rect 26836 6496 26852 6560
rect 26916 6496 26922 6560
rect 26606 6495 26922 6496
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 9946 6016 10262 6017
rect 9946 5952 9952 6016
rect 10016 5952 10032 6016
rect 10096 5952 10112 6016
rect 10176 5952 10192 6016
rect 10256 5952 10262 6016
rect 9946 5951 10262 5952
rect 17946 6016 18262 6017
rect 17946 5952 17952 6016
rect 18016 5952 18032 6016
rect 18096 5952 18112 6016
rect 18176 5952 18192 6016
rect 18256 5952 18262 6016
rect 17946 5951 18262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 28349 5810 28415 5813
rect 29200 5810 30000 5840
rect 28349 5808 30000 5810
rect 28349 5752 28354 5808
rect 28410 5752 30000 5808
rect 28349 5750 30000 5752
rect 28349 5747 28415 5750
rect 29200 5720 30000 5750
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 10606 5472 10922 5473
rect 10606 5408 10612 5472
rect 10676 5408 10692 5472
rect 10756 5408 10772 5472
rect 10836 5408 10852 5472
rect 10916 5408 10922 5472
rect 10606 5407 10922 5408
rect 18606 5472 18922 5473
rect 18606 5408 18612 5472
rect 18676 5408 18692 5472
rect 18756 5408 18772 5472
rect 18836 5408 18852 5472
rect 18916 5408 18922 5472
rect 18606 5407 18922 5408
rect 26606 5472 26922 5473
rect 26606 5408 26612 5472
rect 26676 5408 26692 5472
rect 26756 5408 26772 5472
rect 26836 5408 26852 5472
rect 26916 5408 26922 5472
rect 26606 5407 26922 5408
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 9946 4928 10262 4929
rect 9946 4864 9952 4928
rect 10016 4864 10032 4928
rect 10096 4864 10112 4928
rect 10176 4864 10192 4928
rect 10256 4864 10262 4928
rect 9946 4863 10262 4864
rect 17946 4928 18262 4929
rect 17946 4864 17952 4928
rect 18016 4864 18032 4928
rect 18096 4864 18112 4928
rect 18176 4864 18192 4928
rect 18256 4864 18262 4928
rect 17946 4863 18262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 10606 4384 10922 4385
rect 10606 4320 10612 4384
rect 10676 4320 10692 4384
rect 10756 4320 10772 4384
rect 10836 4320 10852 4384
rect 10916 4320 10922 4384
rect 10606 4319 10922 4320
rect 18606 4384 18922 4385
rect 18606 4320 18612 4384
rect 18676 4320 18692 4384
rect 18756 4320 18772 4384
rect 18836 4320 18852 4384
rect 18916 4320 18922 4384
rect 18606 4319 18922 4320
rect 26606 4384 26922 4385
rect 26606 4320 26612 4384
rect 26676 4320 26692 4384
rect 26756 4320 26772 4384
rect 26836 4320 26852 4384
rect 26916 4320 26922 4384
rect 26606 4319 26922 4320
rect 28349 4178 28415 4181
rect 29200 4178 30000 4208
rect 28349 4176 30000 4178
rect 28349 4120 28354 4176
rect 28410 4120 30000 4176
rect 28349 4118 30000 4120
rect 28349 4115 28415 4118
rect 29200 4088 30000 4118
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 9946 3840 10262 3841
rect 9946 3776 9952 3840
rect 10016 3776 10032 3840
rect 10096 3776 10112 3840
rect 10176 3776 10192 3840
rect 10256 3776 10262 3840
rect 9946 3775 10262 3776
rect 17946 3840 18262 3841
rect 17946 3776 17952 3840
rect 18016 3776 18032 3840
rect 18096 3776 18112 3840
rect 18176 3776 18192 3840
rect 18256 3776 18262 3840
rect 17946 3775 18262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 10606 3296 10922 3297
rect 10606 3232 10612 3296
rect 10676 3232 10692 3296
rect 10756 3232 10772 3296
rect 10836 3232 10852 3296
rect 10916 3232 10922 3296
rect 10606 3231 10922 3232
rect 18606 3296 18922 3297
rect 18606 3232 18612 3296
rect 18676 3232 18692 3296
rect 18756 3232 18772 3296
rect 18836 3232 18852 3296
rect 18916 3232 18922 3296
rect 18606 3231 18922 3232
rect 26606 3296 26922 3297
rect 26606 3232 26612 3296
rect 26676 3232 26692 3296
rect 26756 3232 26772 3296
rect 26836 3232 26852 3296
rect 26916 3232 26922 3296
rect 26606 3231 26922 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 9946 2752 10262 2753
rect 9946 2688 9952 2752
rect 10016 2688 10032 2752
rect 10096 2688 10112 2752
rect 10176 2688 10192 2752
rect 10256 2688 10262 2752
rect 9946 2687 10262 2688
rect 17946 2752 18262 2753
rect 17946 2688 17952 2752
rect 18016 2688 18032 2752
rect 18096 2688 18112 2752
rect 18176 2688 18192 2752
rect 18256 2688 18262 2752
rect 17946 2687 18262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 28349 2546 28415 2549
rect 29200 2546 30000 2576
rect 28349 2544 30000 2546
rect 28349 2488 28354 2544
rect 28410 2488 30000 2544
rect 28349 2486 30000 2488
rect 28349 2483 28415 2486
rect 29200 2456 30000 2486
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 10606 2208 10922 2209
rect 10606 2144 10612 2208
rect 10676 2144 10692 2208
rect 10756 2144 10772 2208
rect 10836 2144 10852 2208
rect 10916 2144 10922 2208
rect 10606 2143 10922 2144
rect 18606 2208 18922 2209
rect 18606 2144 18612 2208
rect 18676 2144 18692 2208
rect 18756 2144 18772 2208
rect 18836 2144 18852 2208
rect 18916 2144 18922 2208
rect 18606 2143 18922 2144
rect 26606 2208 26922 2209
rect 26606 2144 26612 2208
rect 26676 2144 26692 2208
rect 26756 2144 26772 2208
rect 26836 2144 26852 2208
rect 26916 2144 26922 2208
rect 26606 2143 26922 2144
<< via3 >>
rect 1952 27772 2016 27776
rect 1952 27716 1956 27772
rect 1956 27716 2012 27772
rect 2012 27716 2016 27772
rect 1952 27712 2016 27716
rect 2032 27772 2096 27776
rect 2032 27716 2036 27772
rect 2036 27716 2092 27772
rect 2092 27716 2096 27772
rect 2032 27712 2096 27716
rect 2112 27772 2176 27776
rect 2112 27716 2116 27772
rect 2116 27716 2172 27772
rect 2172 27716 2176 27772
rect 2112 27712 2176 27716
rect 2192 27772 2256 27776
rect 2192 27716 2196 27772
rect 2196 27716 2252 27772
rect 2252 27716 2256 27772
rect 2192 27712 2256 27716
rect 9952 27772 10016 27776
rect 9952 27716 9956 27772
rect 9956 27716 10012 27772
rect 10012 27716 10016 27772
rect 9952 27712 10016 27716
rect 10032 27772 10096 27776
rect 10032 27716 10036 27772
rect 10036 27716 10092 27772
rect 10092 27716 10096 27772
rect 10032 27712 10096 27716
rect 10112 27772 10176 27776
rect 10112 27716 10116 27772
rect 10116 27716 10172 27772
rect 10172 27716 10176 27772
rect 10112 27712 10176 27716
rect 10192 27772 10256 27776
rect 10192 27716 10196 27772
rect 10196 27716 10252 27772
rect 10252 27716 10256 27772
rect 10192 27712 10256 27716
rect 17952 27772 18016 27776
rect 17952 27716 17956 27772
rect 17956 27716 18012 27772
rect 18012 27716 18016 27772
rect 17952 27712 18016 27716
rect 18032 27772 18096 27776
rect 18032 27716 18036 27772
rect 18036 27716 18092 27772
rect 18092 27716 18096 27772
rect 18032 27712 18096 27716
rect 18112 27772 18176 27776
rect 18112 27716 18116 27772
rect 18116 27716 18172 27772
rect 18172 27716 18176 27772
rect 18112 27712 18176 27716
rect 18192 27772 18256 27776
rect 18192 27716 18196 27772
rect 18196 27716 18252 27772
rect 18252 27716 18256 27772
rect 18192 27712 18256 27716
rect 25952 27772 26016 27776
rect 25952 27716 25956 27772
rect 25956 27716 26012 27772
rect 26012 27716 26016 27772
rect 25952 27712 26016 27716
rect 26032 27772 26096 27776
rect 26032 27716 26036 27772
rect 26036 27716 26092 27772
rect 26092 27716 26096 27772
rect 26032 27712 26096 27716
rect 26112 27772 26176 27776
rect 26112 27716 26116 27772
rect 26116 27716 26172 27772
rect 26172 27716 26176 27772
rect 26112 27712 26176 27716
rect 26192 27772 26256 27776
rect 26192 27716 26196 27772
rect 26196 27716 26252 27772
rect 26252 27716 26256 27772
rect 26192 27712 26256 27716
rect 2612 27228 2676 27232
rect 2612 27172 2616 27228
rect 2616 27172 2672 27228
rect 2672 27172 2676 27228
rect 2612 27168 2676 27172
rect 2692 27228 2756 27232
rect 2692 27172 2696 27228
rect 2696 27172 2752 27228
rect 2752 27172 2756 27228
rect 2692 27168 2756 27172
rect 2772 27228 2836 27232
rect 2772 27172 2776 27228
rect 2776 27172 2832 27228
rect 2832 27172 2836 27228
rect 2772 27168 2836 27172
rect 2852 27228 2916 27232
rect 2852 27172 2856 27228
rect 2856 27172 2912 27228
rect 2912 27172 2916 27228
rect 2852 27168 2916 27172
rect 10612 27228 10676 27232
rect 10612 27172 10616 27228
rect 10616 27172 10672 27228
rect 10672 27172 10676 27228
rect 10612 27168 10676 27172
rect 10692 27228 10756 27232
rect 10692 27172 10696 27228
rect 10696 27172 10752 27228
rect 10752 27172 10756 27228
rect 10692 27168 10756 27172
rect 10772 27228 10836 27232
rect 10772 27172 10776 27228
rect 10776 27172 10832 27228
rect 10832 27172 10836 27228
rect 10772 27168 10836 27172
rect 10852 27228 10916 27232
rect 10852 27172 10856 27228
rect 10856 27172 10912 27228
rect 10912 27172 10916 27228
rect 10852 27168 10916 27172
rect 18612 27228 18676 27232
rect 18612 27172 18616 27228
rect 18616 27172 18672 27228
rect 18672 27172 18676 27228
rect 18612 27168 18676 27172
rect 18692 27228 18756 27232
rect 18692 27172 18696 27228
rect 18696 27172 18752 27228
rect 18752 27172 18756 27228
rect 18692 27168 18756 27172
rect 18772 27228 18836 27232
rect 18772 27172 18776 27228
rect 18776 27172 18832 27228
rect 18832 27172 18836 27228
rect 18772 27168 18836 27172
rect 18852 27228 18916 27232
rect 18852 27172 18856 27228
rect 18856 27172 18912 27228
rect 18912 27172 18916 27228
rect 18852 27168 18916 27172
rect 26612 27228 26676 27232
rect 26612 27172 26616 27228
rect 26616 27172 26672 27228
rect 26672 27172 26676 27228
rect 26612 27168 26676 27172
rect 26692 27228 26756 27232
rect 26692 27172 26696 27228
rect 26696 27172 26752 27228
rect 26752 27172 26756 27228
rect 26692 27168 26756 27172
rect 26772 27228 26836 27232
rect 26772 27172 26776 27228
rect 26776 27172 26832 27228
rect 26832 27172 26836 27228
rect 26772 27168 26836 27172
rect 26852 27228 26916 27232
rect 26852 27172 26856 27228
rect 26856 27172 26912 27228
rect 26912 27172 26916 27228
rect 26852 27168 26916 27172
rect 1952 26684 2016 26688
rect 1952 26628 1956 26684
rect 1956 26628 2012 26684
rect 2012 26628 2016 26684
rect 1952 26624 2016 26628
rect 2032 26684 2096 26688
rect 2032 26628 2036 26684
rect 2036 26628 2092 26684
rect 2092 26628 2096 26684
rect 2032 26624 2096 26628
rect 2112 26684 2176 26688
rect 2112 26628 2116 26684
rect 2116 26628 2172 26684
rect 2172 26628 2176 26684
rect 2112 26624 2176 26628
rect 2192 26684 2256 26688
rect 2192 26628 2196 26684
rect 2196 26628 2252 26684
rect 2252 26628 2256 26684
rect 2192 26624 2256 26628
rect 9952 26684 10016 26688
rect 9952 26628 9956 26684
rect 9956 26628 10012 26684
rect 10012 26628 10016 26684
rect 9952 26624 10016 26628
rect 10032 26684 10096 26688
rect 10032 26628 10036 26684
rect 10036 26628 10092 26684
rect 10092 26628 10096 26684
rect 10032 26624 10096 26628
rect 10112 26684 10176 26688
rect 10112 26628 10116 26684
rect 10116 26628 10172 26684
rect 10172 26628 10176 26684
rect 10112 26624 10176 26628
rect 10192 26684 10256 26688
rect 10192 26628 10196 26684
rect 10196 26628 10252 26684
rect 10252 26628 10256 26684
rect 10192 26624 10256 26628
rect 17952 26684 18016 26688
rect 17952 26628 17956 26684
rect 17956 26628 18012 26684
rect 18012 26628 18016 26684
rect 17952 26624 18016 26628
rect 18032 26684 18096 26688
rect 18032 26628 18036 26684
rect 18036 26628 18092 26684
rect 18092 26628 18096 26684
rect 18032 26624 18096 26628
rect 18112 26684 18176 26688
rect 18112 26628 18116 26684
rect 18116 26628 18172 26684
rect 18172 26628 18176 26684
rect 18112 26624 18176 26628
rect 18192 26684 18256 26688
rect 18192 26628 18196 26684
rect 18196 26628 18252 26684
rect 18252 26628 18256 26684
rect 18192 26624 18256 26628
rect 25952 26684 26016 26688
rect 25952 26628 25956 26684
rect 25956 26628 26012 26684
rect 26012 26628 26016 26684
rect 25952 26624 26016 26628
rect 26032 26684 26096 26688
rect 26032 26628 26036 26684
rect 26036 26628 26092 26684
rect 26092 26628 26096 26684
rect 26032 26624 26096 26628
rect 26112 26684 26176 26688
rect 26112 26628 26116 26684
rect 26116 26628 26172 26684
rect 26172 26628 26176 26684
rect 26112 26624 26176 26628
rect 26192 26684 26256 26688
rect 26192 26628 26196 26684
rect 26196 26628 26252 26684
rect 26252 26628 26256 26684
rect 26192 26624 26256 26628
rect 2612 26140 2676 26144
rect 2612 26084 2616 26140
rect 2616 26084 2672 26140
rect 2672 26084 2676 26140
rect 2612 26080 2676 26084
rect 2692 26140 2756 26144
rect 2692 26084 2696 26140
rect 2696 26084 2752 26140
rect 2752 26084 2756 26140
rect 2692 26080 2756 26084
rect 2772 26140 2836 26144
rect 2772 26084 2776 26140
rect 2776 26084 2832 26140
rect 2832 26084 2836 26140
rect 2772 26080 2836 26084
rect 2852 26140 2916 26144
rect 2852 26084 2856 26140
rect 2856 26084 2912 26140
rect 2912 26084 2916 26140
rect 2852 26080 2916 26084
rect 10612 26140 10676 26144
rect 10612 26084 10616 26140
rect 10616 26084 10672 26140
rect 10672 26084 10676 26140
rect 10612 26080 10676 26084
rect 10692 26140 10756 26144
rect 10692 26084 10696 26140
rect 10696 26084 10752 26140
rect 10752 26084 10756 26140
rect 10692 26080 10756 26084
rect 10772 26140 10836 26144
rect 10772 26084 10776 26140
rect 10776 26084 10832 26140
rect 10832 26084 10836 26140
rect 10772 26080 10836 26084
rect 10852 26140 10916 26144
rect 10852 26084 10856 26140
rect 10856 26084 10912 26140
rect 10912 26084 10916 26140
rect 10852 26080 10916 26084
rect 18612 26140 18676 26144
rect 18612 26084 18616 26140
rect 18616 26084 18672 26140
rect 18672 26084 18676 26140
rect 18612 26080 18676 26084
rect 18692 26140 18756 26144
rect 18692 26084 18696 26140
rect 18696 26084 18752 26140
rect 18752 26084 18756 26140
rect 18692 26080 18756 26084
rect 18772 26140 18836 26144
rect 18772 26084 18776 26140
rect 18776 26084 18832 26140
rect 18832 26084 18836 26140
rect 18772 26080 18836 26084
rect 18852 26140 18916 26144
rect 18852 26084 18856 26140
rect 18856 26084 18912 26140
rect 18912 26084 18916 26140
rect 18852 26080 18916 26084
rect 26612 26140 26676 26144
rect 26612 26084 26616 26140
rect 26616 26084 26672 26140
rect 26672 26084 26676 26140
rect 26612 26080 26676 26084
rect 26692 26140 26756 26144
rect 26692 26084 26696 26140
rect 26696 26084 26752 26140
rect 26752 26084 26756 26140
rect 26692 26080 26756 26084
rect 26772 26140 26836 26144
rect 26772 26084 26776 26140
rect 26776 26084 26832 26140
rect 26832 26084 26836 26140
rect 26772 26080 26836 26084
rect 26852 26140 26916 26144
rect 26852 26084 26856 26140
rect 26856 26084 26912 26140
rect 26912 26084 26916 26140
rect 26852 26080 26916 26084
rect 1952 25596 2016 25600
rect 1952 25540 1956 25596
rect 1956 25540 2012 25596
rect 2012 25540 2016 25596
rect 1952 25536 2016 25540
rect 2032 25596 2096 25600
rect 2032 25540 2036 25596
rect 2036 25540 2092 25596
rect 2092 25540 2096 25596
rect 2032 25536 2096 25540
rect 2112 25596 2176 25600
rect 2112 25540 2116 25596
rect 2116 25540 2172 25596
rect 2172 25540 2176 25596
rect 2112 25536 2176 25540
rect 2192 25596 2256 25600
rect 2192 25540 2196 25596
rect 2196 25540 2252 25596
rect 2252 25540 2256 25596
rect 2192 25536 2256 25540
rect 9952 25596 10016 25600
rect 9952 25540 9956 25596
rect 9956 25540 10012 25596
rect 10012 25540 10016 25596
rect 9952 25536 10016 25540
rect 10032 25596 10096 25600
rect 10032 25540 10036 25596
rect 10036 25540 10092 25596
rect 10092 25540 10096 25596
rect 10032 25536 10096 25540
rect 10112 25596 10176 25600
rect 10112 25540 10116 25596
rect 10116 25540 10172 25596
rect 10172 25540 10176 25596
rect 10112 25536 10176 25540
rect 10192 25596 10256 25600
rect 10192 25540 10196 25596
rect 10196 25540 10252 25596
rect 10252 25540 10256 25596
rect 10192 25536 10256 25540
rect 17952 25596 18016 25600
rect 17952 25540 17956 25596
rect 17956 25540 18012 25596
rect 18012 25540 18016 25596
rect 17952 25536 18016 25540
rect 18032 25596 18096 25600
rect 18032 25540 18036 25596
rect 18036 25540 18092 25596
rect 18092 25540 18096 25596
rect 18032 25536 18096 25540
rect 18112 25596 18176 25600
rect 18112 25540 18116 25596
rect 18116 25540 18172 25596
rect 18172 25540 18176 25596
rect 18112 25536 18176 25540
rect 18192 25596 18256 25600
rect 18192 25540 18196 25596
rect 18196 25540 18252 25596
rect 18252 25540 18256 25596
rect 18192 25536 18256 25540
rect 25952 25596 26016 25600
rect 25952 25540 25956 25596
rect 25956 25540 26012 25596
rect 26012 25540 26016 25596
rect 25952 25536 26016 25540
rect 26032 25596 26096 25600
rect 26032 25540 26036 25596
rect 26036 25540 26092 25596
rect 26092 25540 26096 25596
rect 26032 25536 26096 25540
rect 26112 25596 26176 25600
rect 26112 25540 26116 25596
rect 26116 25540 26172 25596
rect 26172 25540 26176 25596
rect 26112 25536 26176 25540
rect 26192 25596 26256 25600
rect 26192 25540 26196 25596
rect 26196 25540 26252 25596
rect 26252 25540 26256 25596
rect 26192 25536 26256 25540
rect 2612 25052 2676 25056
rect 2612 24996 2616 25052
rect 2616 24996 2672 25052
rect 2672 24996 2676 25052
rect 2612 24992 2676 24996
rect 2692 25052 2756 25056
rect 2692 24996 2696 25052
rect 2696 24996 2752 25052
rect 2752 24996 2756 25052
rect 2692 24992 2756 24996
rect 2772 25052 2836 25056
rect 2772 24996 2776 25052
rect 2776 24996 2832 25052
rect 2832 24996 2836 25052
rect 2772 24992 2836 24996
rect 2852 25052 2916 25056
rect 2852 24996 2856 25052
rect 2856 24996 2912 25052
rect 2912 24996 2916 25052
rect 2852 24992 2916 24996
rect 10612 25052 10676 25056
rect 10612 24996 10616 25052
rect 10616 24996 10672 25052
rect 10672 24996 10676 25052
rect 10612 24992 10676 24996
rect 10692 25052 10756 25056
rect 10692 24996 10696 25052
rect 10696 24996 10752 25052
rect 10752 24996 10756 25052
rect 10692 24992 10756 24996
rect 10772 25052 10836 25056
rect 10772 24996 10776 25052
rect 10776 24996 10832 25052
rect 10832 24996 10836 25052
rect 10772 24992 10836 24996
rect 10852 25052 10916 25056
rect 10852 24996 10856 25052
rect 10856 24996 10912 25052
rect 10912 24996 10916 25052
rect 10852 24992 10916 24996
rect 18612 25052 18676 25056
rect 18612 24996 18616 25052
rect 18616 24996 18672 25052
rect 18672 24996 18676 25052
rect 18612 24992 18676 24996
rect 18692 25052 18756 25056
rect 18692 24996 18696 25052
rect 18696 24996 18752 25052
rect 18752 24996 18756 25052
rect 18692 24992 18756 24996
rect 18772 25052 18836 25056
rect 18772 24996 18776 25052
rect 18776 24996 18832 25052
rect 18832 24996 18836 25052
rect 18772 24992 18836 24996
rect 18852 25052 18916 25056
rect 18852 24996 18856 25052
rect 18856 24996 18912 25052
rect 18912 24996 18916 25052
rect 18852 24992 18916 24996
rect 26612 25052 26676 25056
rect 26612 24996 26616 25052
rect 26616 24996 26672 25052
rect 26672 24996 26676 25052
rect 26612 24992 26676 24996
rect 26692 25052 26756 25056
rect 26692 24996 26696 25052
rect 26696 24996 26752 25052
rect 26752 24996 26756 25052
rect 26692 24992 26756 24996
rect 26772 25052 26836 25056
rect 26772 24996 26776 25052
rect 26776 24996 26832 25052
rect 26832 24996 26836 25052
rect 26772 24992 26836 24996
rect 26852 25052 26916 25056
rect 26852 24996 26856 25052
rect 26856 24996 26912 25052
rect 26912 24996 26916 25052
rect 26852 24992 26916 24996
rect 1952 24508 2016 24512
rect 1952 24452 1956 24508
rect 1956 24452 2012 24508
rect 2012 24452 2016 24508
rect 1952 24448 2016 24452
rect 2032 24508 2096 24512
rect 2032 24452 2036 24508
rect 2036 24452 2092 24508
rect 2092 24452 2096 24508
rect 2032 24448 2096 24452
rect 2112 24508 2176 24512
rect 2112 24452 2116 24508
rect 2116 24452 2172 24508
rect 2172 24452 2176 24508
rect 2112 24448 2176 24452
rect 2192 24508 2256 24512
rect 2192 24452 2196 24508
rect 2196 24452 2252 24508
rect 2252 24452 2256 24508
rect 2192 24448 2256 24452
rect 9952 24508 10016 24512
rect 9952 24452 9956 24508
rect 9956 24452 10012 24508
rect 10012 24452 10016 24508
rect 9952 24448 10016 24452
rect 10032 24508 10096 24512
rect 10032 24452 10036 24508
rect 10036 24452 10092 24508
rect 10092 24452 10096 24508
rect 10032 24448 10096 24452
rect 10112 24508 10176 24512
rect 10112 24452 10116 24508
rect 10116 24452 10172 24508
rect 10172 24452 10176 24508
rect 10112 24448 10176 24452
rect 10192 24508 10256 24512
rect 10192 24452 10196 24508
rect 10196 24452 10252 24508
rect 10252 24452 10256 24508
rect 10192 24448 10256 24452
rect 17952 24508 18016 24512
rect 17952 24452 17956 24508
rect 17956 24452 18012 24508
rect 18012 24452 18016 24508
rect 17952 24448 18016 24452
rect 18032 24508 18096 24512
rect 18032 24452 18036 24508
rect 18036 24452 18092 24508
rect 18092 24452 18096 24508
rect 18032 24448 18096 24452
rect 18112 24508 18176 24512
rect 18112 24452 18116 24508
rect 18116 24452 18172 24508
rect 18172 24452 18176 24508
rect 18112 24448 18176 24452
rect 18192 24508 18256 24512
rect 18192 24452 18196 24508
rect 18196 24452 18252 24508
rect 18252 24452 18256 24508
rect 18192 24448 18256 24452
rect 25952 24508 26016 24512
rect 25952 24452 25956 24508
rect 25956 24452 26012 24508
rect 26012 24452 26016 24508
rect 25952 24448 26016 24452
rect 26032 24508 26096 24512
rect 26032 24452 26036 24508
rect 26036 24452 26092 24508
rect 26092 24452 26096 24508
rect 26032 24448 26096 24452
rect 26112 24508 26176 24512
rect 26112 24452 26116 24508
rect 26116 24452 26172 24508
rect 26172 24452 26176 24508
rect 26112 24448 26176 24452
rect 26192 24508 26256 24512
rect 26192 24452 26196 24508
rect 26196 24452 26252 24508
rect 26252 24452 26256 24508
rect 26192 24448 26256 24452
rect 2612 23964 2676 23968
rect 2612 23908 2616 23964
rect 2616 23908 2672 23964
rect 2672 23908 2676 23964
rect 2612 23904 2676 23908
rect 2692 23964 2756 23968
rect 2692 23908 2696 23964
rect 2696 23908 2752 23964
rect 2752 23908 2756 23964
rect 2692 23904 2756 23908
rect 2772 23964 2836 23968
rect 2772 23908 2776 23964
rect 2776 23908 2832 23964
rect 2832 23908 2836 23964
rect 2772 23904 2836 23908
rect 2852 23964 2916 23968
rect 2852 23908 2856 23964
rect 2856 23908 2912 23964
rect 2912 23908 2916 23964
rect 2852 23904 2916 23908
rect 10612 23964 10676 23968
rect 10612 23908 10616 23964
rect 10616 23908 10672 23964
rect 10672 23908 10676 23964
rect 10612 23904 10676 23908
rect 10692 23964 10756 23968
rect 10692 23908 10696 23964
rect 10696 23908 10752 23964
rect 10752 23908 10756 23964
rect 10692 23904 10756 23908
rect 10772 23964 10836 23968
rect 10772 23908 10776 23964
rect 10776 23908 10832 23964
rect 10832 23908 10836 23964
rect 10772 23904 10836 23908
rect 10852 23964 10916 23968
rect 10852 23908 10856 23964
rect 10856 23908 10912 23964
rect 10912 23908 10916 23964
rect 10852 23904 10916 23908
rect 18612 23964 18676 23968
rect 18612 23908 18616 23964
rect 18616 23908 18672 23964
rect 18672 23908 18676 23964
rect 18612 23904 18676 23908
rect 18692 23964 18756 23968
rect 18692 23908 18696 23964
rect 18696 23908 18752 23964
rect 18752 23908 18756 23964
rect 18692 23904 18756 23908
rect 18772 23964 18836 23968
rect 18772 23908 18776 23964
rect 18776 23908 18832 23964
rect 18832 23908 18836 23964
rect 18772 23904 18836 23908
rect 18852 23964 18916 23968
rect 18852 23908 18856 23964
rect 18856 23908 18912 23964
rect 18912 23908 18916 23964
rect 18852 23904 18916 23908
rect 26612 23964 26676 23968
rect 26612 23908 26616 23964
rect 26616 23908 26672 23964
rect 26672 23908 26676 23964
rect 26612 23904 26676 23908
rect 26692 23964 26756 23968
rect 26692 23908 26696 23964
rect 26696 23908 26752 23964
rect 26752 23908 26756 23964
rect 26692 23904 26756 23908
rect 26772 23964 26836 23968
rect 26772 23908 26776 23964
rect 26776 23908 26832 23964
rect 26832 23908 26836 23964
rect 26772 23904 26836 23908
rect 26852 23964 26916 23968
rect 26852 23908 26856 23964
rect 26856 23908 26912 23964
rect 26912 23908 26916 23964
rect 26852 23904 26916 23908
rect 1952 23420 2016 23424
rect 1952 23364 1956 23420
rect 1956 23364 2012 23420
rect 2012 23364 2016 23420
rect 1952 23360 2016 23364
rect 2032 23420 2096 23424
rect 2032 23364 2036 23420
rect 2036 23364 2092 23420
rect 2092 23364 2096 23420
rect 2032 23360 2096 23364
rect 2112 23420 2176 23424
rect 2112 23364 2116 23420
rect 2116 23364 2172 23420
rect 2172 23364 2176 23420
rect 2112 23360 2176 23364
rect 2192 23420 2256 23424
rect 2192 23364 2196 23420
rect 2196 23364 2252 23420
rect 2252 23364 2256 23420
rect 2192 23360 2256 23364
rect 9952 23420 10016 23424
rect 9952 23364 9956 23420
rect 9956 23364 10012 23420
rect 10012 23364 10016 23420
rect 9952 23360 10016 23364
rect 10032 23420 10096 23424
rect 10032 23364 10036 23420
rect 10036 23364 10092 23420
rect 10092 23364 10096 23420
rect 10032 23360 10096 23364
rect 10112 23420 10176 23424
rect 10112 23364 10116 23420
rect 10116 23364 10172 23420
rect 10172 23364 10176 23420
rect 10112 23360 10176 23364
rect 10192 23420 10256 23424
rect 10192 23364 10196 23420
rect 10196 23364 10252 23420
rect 10252 23364 10256 23420
rect 10192 23360 10256 23364
rect 17952 23420 18016 23424
rect 17952 23364 17956 23420
rect 17956 23364 18012 23420
rect 18012 23364 18016 23420
rect 17952 23360 18016 23364
rect 18032 23420 18096 23424
rect 18032 23364 18036 23420
rect 18036 23364 18092 23420
rect 18092 23364 18096 23420
rect 18032 23360 18096 23364
rect 18112 23420 18176 23424
rect 18112 23364 18116 23420
rect 18116 23364 18172 23420
rect 18172 23364 18176 23420
rect 18112 23360 18176 23364
rect 18192 23420 18256 23424
rect 18192 23364 18196 23420
rect 18196 23364 18252 23420
rect 18252 23364 18256 23420
rect 18192 23360 18256 23364
rect 25952 23420 26016 23424
rect 25952 23364 25956 23420
rect 25956 23364 26012 23420
rect 26012 23364 26016 23420
rect 25952 23360 26016 23364
rect 26032 23420 26096 23424
rect 26032 23364 26036 23420
rect 26036 23364 26092 23420
rect 26092 23364 26096 23420
rect 26032 23360 26096 23364
rect 26112 23420 26176 23424
rect 26112 23364 26116 23420
rect 26116 23364 26172 23420
rect 26172 23364 26176 23420
rect 26112 23360 26176 23364
rect 26192 23420 26256 23424
rect 26192 23364 26196 23420
rect 26196 23364 26252 23420
rect 26252 23364 26256 23420
rect 26192 23360 26256 23364
rect 2612 22876 2676 22880
rect 2612 22820 2616 22876
rect 2616 22820 2672 22876
rect 2672 22820 2676 22876
rect 2612 22816 2676 22820
rect 2692 22876 2756 22880
rect 2692 22820 2696 22876
rect 2696 22820 2752 22876
rect 2752 22820 2756 22876
rect 2692 22816 2756 22820
rect 2772 22876 2836 22880
rect 2772 22820 2776 22876
rect 2776 22820 2832 22876
rect 2832 22820 2836 22876
rect 2772 22816 2836 22820
rect 2852 22876 2916 22880
rect 2852 22820 2856 22876
rect 2856 22820 2912 22876
rect 2912 22820 2916 22876
rect 2852 22816 2916 22820
rect 10612 22876 10676 22880
rect 10612 22820 10616 22876
rect 10616 22820 10672 22876
rect 10672 22820 10676 22876
rect 10612 22816 10676 22820
rect 10692 22876 10756 22880
rect 10692 22820 10696 22876
rect 10696 22820 10752 22876
rect 10752 22820 10756 22876
rect 10692 22816 10756 22820
rect 10772 22876 10836 22880
rect 10772 22820 10776 22876
rect 10776 22820 10832 22876
rect 10832 22820 10836 22876
rect 10772 22816 10836 22820
rect 10852 22876 10916 22880
rect 10852 22820 10856 22876
rect 10856 22820 10912 22876
rect 10912 22820 10916 22876
rect 10852 22816 10916 22820
rect 18612 22876 18676 22880
rect 18612 22820 18616 22876
rect 18616 22820 18672 22876
rect 18672 22820 18676 22876
rect 18612 22816 18676 22820
rect 18692 22876 18756 22880
rect 18692 22820 18696 22876
rect 18696 22820 18752 22876
rect 18752 22820 18756 22876
rect 18692 22816 18756 22820
rect 18772 22876 18836 22880
rect 18772 22820 18776 22876
rect 18776 22820 18832 22876
rect 18832 22820 18836 22876
rect 18772 22816 18836 22820
rect 18852 22876 18916 22880
rect 18852 22820 18856 22876
rect 18856 22820 18912 22876
rect 18912 22820 18916 22876
rect 18852 22816 18916 22820
rect 26612 22876 26676 22880
rect 26612 22820 26616 22876
rect 26616 22820 26672 22876
rect 26672 22820 26676 22876
rect 26612 22816 26676 22820
rect 26692 22876 26756 22880
rect 26692 22820 26696 22876
rect 26696 22820 26752 22876
rect 26752 22820 26756 22876
rect 26692 22816 26756 22820
rect 26772 22876 26836 22880
rect 26772 22820 26776 22876
rect 26776 22820 26832 22876
rect 26832 22820 26836 22876
rect 26772 22816 26836 22820
rect 26852 22876 26916 22880
rect 26852 22820 26856 22876
rect 26856 22820 26912 22876
rect 26912 22820 26916 22876
rect 26852 22816 26916 22820
rect 1952 22332 2016 22336
rect 1952 22276 1956 22332
rect 1956 22276 2012 22332
rect 2012 22276 2016 22332
rect 1952 22272 2016 22276
rect 2032 22332 2096 22336
rect 2032 22276 2036 22332
rect 2036 22276 2092 22332
rect 2092 22276 2096 22332
rect 2032 22272 2096 22276
rect 2112 22332 2176 22336
rect 2112 22276 2116 22332
rect 2116 22276 2172 22332
rect 2172 22276 2176 22332
rect 2112 22272 2176 22276
rect 2192 22332 2256 22336
rect 2192 22276 2196 22332
rect 2196 22276 2252 22332
rect 2252 22276 2256 22332
rect 2192 22272 2256 22276
rect 9952 22332 10016 22336
rect 9952 22276 9956 22332
rect 9956 22276 10012 22332
rect 10012 22276 10016 22332
rect 9952 22272 10016 22276
rect 10032 22332 10096 22336
rect 10032 22276 10036 22332
rect 10036 22276 10092 22332
rect 10092 22276 10096 22332
rect 10032 22272 10096 22276
rect 10112 22332 10176 22336
rect 10112 22276 10116 22332
rect 10116 22276 10172 22332
rect 10172 22276 10176 22332
rect 10112 22272 10176 22276
rect 10192 22332 10256 22336
rect 10192 22276 10196 22332
rect 10196 22276 10252 22332
rect 10252 22276 10256 22332
rect 10192 22272 10256 22276
rect 17952 22332 18016 22336
rect 17952 22276 17956 22332
rect 17956 22276 18012 22332
rect 18012 22276 18016 22332
rect 17952 22272 18016 22276
rect 18032 22332 18096 22336
rect 18032 22276 18036 22332
rect 18036 22276 18092 22332
rect 18092 22276 18096 22332
rect 18032 22272 18096 22276
rect 18112 22332 18176 22336
rect 18112 22276 18116 22332
rect 18116 22276 18172 22332
rect 18172 22276 18176 22332
rect 18112 22272 18176 22276
rect 18192 22332 18256 22336
rect 18192 22276 18196 22332
rect 18196 22276 18252 22332
rect 18252 22276 18256 22332
rect 18192 22272 18256 22276
rect 25952 22332 26016 22336
rect 25952 22276 25956 22332
rect 25956 22276 26012 22332
rect 26012 22276 26016 22332
rect 25952 22272 26016 22276
rect 26032 22332 26096 22336
rect 26032 22276 26036 22332
rect 26036 22276 26092 22332
rect 26092 22276 26096 22332
rect 26032 22272 26096 22276
rect 26112 22332 26176 22336
rect 26112 22276 26116 22332
rect 26116 22276 26172 22332
rect 26172 22276 26176 22332
rect 26112 22272 26176 22276
rect 26192 22332 26256 22336
rect 26192 22276 26196 22332
rect 26196 22276 26252 22332
rect 26252 22276 26256 22332
rect 26192 22272 26256 22276
rect 2612 21788 2676 21792
rect 2612 21732 2616 21788
rect 2616 21732 2672 21788
rect 2672 21732 2676 21788
rect 2612 21728 2676 21732
rect 2692 21788 2756 21792
rect 2692 21732 2696 21788
rect 2696 21732 2752 21788
rect 2752 21732 2756 21788
rect 2692 21728 2756 21732
rect 2772 21788 2836 21792
rect 2772 21732 2776 21788
rect 2776 21732 2832 21788
rect 2832 21732 2836 21788
rect 2772 21728 2836 21732
rect 2852 21788 2916 21792
rect 2852 21732 2856 21788
rect 2856 21732 2912 21788
rect 2912 21732 2916 21788
rect 2852 21728 2916 21732
rect 10612 21788 10676 21792
rect 10612 21732 10616 21788
rect 10616 21732 10672 21788
rect 10672 21732 10676 21788
rect 10612 21728 10676 21732
rect 10692 21788 10756 21792
rect 10692 21732 10696 21788
rect 10696 21732 10752 21788
rect 10752 21732 10756 21788
rect 10692 21728 10756 21732
rect 10772 21788 10836 21792
rect 10772 21732 10776 21788
rect 10776 21732 10832 21788
rect 10832 21732 10836 21788
rect 10772 21728 10836 21732
rect 10852 21788 10916 21792
rect 10852 21732 10856 21788
rect 10856 21732 10912 21788
rect 10912 21732 10916 21788
rect 10852 21728 10916 21732
rect 18612 21788 18676 21792
rect 18612 21732 18616 21788
rect 18616 21732 18672 21788
rect 18672 21732 18676 21788
rect 18612 21728 18676 21732
rect 18692 21788 18756 21792
rect 18692 21732 18696 21788
rect 18696 21732 18752 21788
rect 18752 21732 18756 21788
rect 18692 21728 18756 21732
rect 18772 21788 18836 21792
rect 18772 21732 18776 21788
rect 18776 21732 18832 21788
rect 18832 21732 18836 21788
rect 18772 21728 18836 21732
rect 18852 21788 18916 21792
rect 18852 21732 18856 21788
rect 18856 21732 18912 21788
rect 18912 21732 18916 21788
rect 18852 21728 18916 21732
rect 26612 21788 26676 21792
rect 26612 21732 26616 21788
rect 26616 21732 26672 21788
rect 26672 21732 26676 21788
rect 26612 21728 26676 21732
rect 26692 21788 26756 21792
rect 26692 21732 26696 21788
rect 26696 21732 26752 21788
rect 26752 21732 26756 21788
rect 26692 21728 26756 21732
rect 26772 21788 26836 21792
rect 26772 21732 26776 21788
rect 26776 21732 26832 21788
rect 26832 21732 26836 21788
rect 26772 21728 26836 21732
rect 26852 21788 26916 21792
rect 26852 21732 26856 21788
rect 26856 21732 26912 21788
rect 26912 21732 26916 21788
rect 26852 21728 26916 21732
rect 1952 21244 2016 21248
rect 1952 21188 1956 21244
rect 1956 21188 2012 21244
rect 2012 21188 2016 21244
rect 1952 21184 2016 21188
rect 2032 21244 2096 21248
rect 2032 21188 2036 21244
rect 2036 21188 2092 21244
rect 2092 21188 2096 21244
rect 2032 21184 2096 21188
rect 2112 21244 2176 21248
rect 2112 21188 2116 21244
rect 2116 21188 2172 21244
rect 2172 21188 2176 21244
rect 2112 21184 2176 21188
rect 2192 21244 2256 21248
rect 2192 21188 2196 21244
rect 2196 21188 2252 21244
rect 2252 21188 2256 21244
rect 2192 21184 2256 21188
rect 9952 21244 10016 21248
rect 9952 21188 9956 21244
rect 9956 21188 10012 21244
rect 10012 21188 10016 21244
rect 9952 21184 10016 21188
rect 10032 21244 10096 21248
rect 10032 21188 10036 21244
rect 10036 21188 10092 21244
rect 10092 21188 10096 21244
rect 10032 21184 10096 21188
rect 10112 21244 10176 21248
rect 10112 21188 10116 21244
rect 10116 21188 10172 21244
rect 10172 21188 10176 21244
rect 10112 21184 10176 21188
rect 10192 21244 10256 21248
rect 10192 21188 10196 21244
rect 10196 21188 10252 21244
rect 10252 21188 10256 21244
rect 10192 21184 10256 21188
rect 17952 21244 18016 21248
rect 17952 21188 17956 21244
rect 17956 21188 18012 21244
rect 18012 21188 18016 21244
rect 17952 21184 18016 21188
rect 18032 21244 18096 21248
rect 18032 21188 18036 21244
rect 18036 21188 18092 21244
rect 18092 21188 18096 21244
rect 18032 21184 18096 21188
rect 18112 21244 18176 21248
rect 18112 21188 18116 21244
rect 18116 21188 18172 21244
rect 18172 21188 18176 21244
rect 18112 21184 18176 21188
rect 18192 21244 18256 21248
rect 18192 21188 18196 21244
rect 18196 21188 18252 21244
rect 18252 21188 18256 21244
rect 18192 21184 18256 21188
rect 25952 21244 26016 21248
rect 25952 21188 25956 21244
rect 25956 21188 26012 21244
rect 26012 21188 26016 21244
rect 25952 21184 26016 21188
rect 26032 21244 26096 21248
rect 26032 21188 26036 21244
rect 26036 21188 26092 21244
rect 26092 21188 26096 21244
rect 26032 21184 26096 21188
rect 26112 21244 26176 21248
rect 26112 21188 26116 21244
rect 26116 21188 26172 21244
rect 26172 21188 26176 21244
rect 26112 21184 26176 21188
rect 26192 21244 26256 21248
rect 26192 21188 26196 21244
rect 26196 21188 26252 21244
rect 26252 21188 26256 21244
rect 26192 21184 26256 21188
rect 2612 20700 2676 20704
rect 2612 20644 2616 20700
rect 2616 20644 2672 20700
rect 2672 20644 2676 20700
rect 2612 20640 2676 20644
rect 2692 20700 2756 20704
rect 2692 20644 2696 20700
rect 2696 20644 2752 20700
rect 2752 20644 2756 20700
rect 2692 20640 2756 20644
rect 2772 20700 2836 20704
rect 2772 20644 2776 20700
rect 2776 20644 2832 20700
rect 2832 20644 2836 20700
rect 2772 20640 2836 20644
rect 2852 20700 2916 20704
rect 2852 20644 2856 20700
rect 2856 20644 2912 20700
rect 2912 20644 2916 20700
rect 2852 20640 2916 20644
rect 10612 20700 10676 20704
rect 10612 20644 10616 20700
rect 10616 20644 10672 20700
rect 10672 20644 10676 20700
rect 10612 20640 10676 20644
rect 10692 20700 10756 20704
rect 10692 20644 10696 20700
rect 10696 20644 10752 20700
rect 10752 20644 10756 20700
rect 10692 20640 10756 20644
rect 10772 20700 10836 20704
rect 10772 20644 10776 20700
rect 10776 20644 10832 20700
rect 10832 20644 10836 20700
rect 10772 20640 10836 20644
rect 10852 20700 10916 20704
rect 10852 20644 10856 20700
rect 10856 20644 10912 20700
rect 10912 20644 10916 20700
rect 10852 20640 10916 20644
rect 18612 20700 18676 20704
rect 18612 20644 18616 20700
rect 18616 20644 18672 20700
rect 18672 20644 18676 20700
rect 18612 20640 18676 20644
rect 18692 20700 18756 20704
rect 18692 20644 18696 20700
rect 18696 20644 18752 20700
rect 18752 20644 18756 20700
rect 18692 20640 18756 20644
rect 18772 20700 18836 20704
rect 18772 20644 18776 20700
rect 18776 20644 18832 20700
rect 18832 20644 18836 20700
rect 18772 20640 18836 20644
rect 18852 20700 18916 20704
rect 18852 20644 18856 20700
rect 18856 20644 18912 20700
rect 18912 20644 18916 20700
rect 18852 20640 18916 20644
rect 26612 20700 26676 20704
rect 26612 20644 26616 20700
rect 26616 20644 26672 20700
rect 26672 20644 26676 20700
rect 26612 20640 26676 20644
rect 26692 20700 26756 20704
rect 26692 20644 26696 20700
rect 26696 20644 26752 20700
rect 26752 20644 26756 20700
rect 26692 20640 26756 20644
rect 26772 20700 26836 20704
rect 26772 20644 26776 20700
rect 26776 20644 26832 20700
rect 26832 20644 26836 20700
rect 26772 20640 26836 20644
rect 26852 20700 26916 20704
rect 26852 20644 26856 20700
rect 26856 20644 26912 20700
rect 26912 20644 26916 20700
rect 26852 20640 26916 20644
rect 1952 20156 2016 20160
rect 1952 20100 1956 20156
rect 1956 20100 2012 20156
rect 2012 20100 2016 20156
rect 1952 20096 2016 20100
rect 2032 20156 2096 20160
rect 2032 20100 2036 20156
rect 2036 20100 2092 20156
rect 2092 20100 2096 20156
rect 2032 20096 2096 20100
rect 2112 20156 2176 20160
rect 2112 20100 2116 20156
rect 2116 20100 2172 20156
rect 2172 20100 2176 20156
rect 2112 20096 2176 20100
rect 2192 20156 2256 20160
rect 2192 20100 2196 20156
rect 2196 20100 2252 20156
rect 2252 20100 2256 20156
rect 2192 20096 2256 20100
rect 9952 20156 10016 20160
rect 9952 20100 9956 20156
rect 9956 20100 10012 20156
rect 10012 20100 10016 20156
rect 9952 20096 10016 20100
rect 10032 20156 10096 20160
rect 10032 20100 10036 20156
rect 10036 20100 10092 20156
rect 10092 20100 10096 20156
rect 10032 20096 10096 20100
rect 10112 20156 10176 20160
rect 10112 20100 10116 20156
rect 10116 20100 10172 20156
rect 10172 20100 10176 20156
rect 10112 20096 10176 20100
rect 10192 20156 10256 20160
rect 10192 20100 10196 20156
rect 10196 20100 10252 20156
rect 10252 20100 10256 20156
rect 10192 20096 10256 20100
rect 17952 20156 18016 20160
rect 17952 20100 17956 20156
rect 17956 20100 18012 20156
rect 18012 20100 18016 20156
rect 17952 20096 18016 20100
rect 18032 20156 18096 20160
rect 18032 20100 18036 20156
rect 18036 20100 18092 20156
rect 18092 20100 18096 20156
rect 18032 20096 18096 20100
rect 18112 20156 18176 20160
rect 18112 20100 18116 20156
rect 18116 20100 18172 20156
rect 18172 20100 18176 20156
rect 18112 20096 18176 20100
rect 18192 20156 18256 20160
rect 18192 20100 18196 20156
rect 18196 20100 18252 20156
rect 18252 20100 18256 20156
rect 18192 20096 18256 20100
rect 25952 20156 26016 20160
rect 25952 20100 25956 20156
rect 25956 20100 26012 20156
rect 26012 20100 26016 20156
rect 25952 20096 26016 20100
rect 26032 20156 26096 20160
rect 26032 20100 26036 20156
rect 26036 20100 26092 20156
rect 26092 20100 26096 20156
rect 26032 20096 26096 20100
rect 26112 20156 26176 20160
rect 26112 20100 26116 20156
rect 26116 20100 26172 20156
rect 26172 20100 26176 20156
rect 26112 20096 26176 20100
rect 26192 20156 26256 20160
rect 26192 20100 26196 20156
rect 26196 20100 26252 20156
rect 26252 20100 26256 20156
rect 26192 20096 26256 20100
rect 2612 19612 2676 19616
rect 2612 19556 2616 19612
rect 2616 19556 2672 19612
rect 2672 19556 2676 19612
rect 2612 19552 2676 19556
rect 2692 19612 2756 19616
rect 2692 19556 2696 19612
rect 2696 19556 2752 19612
rect 2752 19556 2756 19612
rect 2692 19552 2756 19556
rect 2772 19612 2836 19616
rect 2772 19556 2776 19612
rect 2776 19556 2832 19612
rect 2832 19556 2836 19612
rect 2772 19552 2836 19556
rect 2852 19612 2916 19616
rect 2852 19556 2856 19612
rect 2856 19556 2912 19612
rect 2912 19556 2916 19612
rect 2852 19552 2916 19556
rect 10612 19612 10676 19616
rect 10612 19556 10616 19612
rect 10616 19556 10672 19612
rect 10672 19556 10676 19612
rect 10612 19552 10676 19556
rect 10692 19612 10756 19616
rect 10692 19556 10696 19612
rect 10696 19556 10752 19612
rect 10752 19556 10756 19612
rect 10692 19552 10756 19556
rect 10772 19612 10836 19616
rect 10772 19556 10776 19612
rect 10776 19556 10832 19612
rect 10832 19556 10836 19612
rect 10772 19552 10836 19556
rect 10852 19612 10916 19616
rect 10852 19556 10856 19612
rect 10856 19556 10912 19612
rect 10912 19556 10916 19612
rect 10852 19552 10916 19556
rect 18612 19612 18676 19616
rect 18612 19556 18616 19612
rect 18616 19556 18672 19612
rect 18672 19556 18676 19612
rect 18612 19552 18676 19556
rect 18692 19612 18756 19616
rect 18692 19556 18696 19612
rect 18696 19556 18752 19612
rect 18752 19556 18756 19612
rect 18692 19552 18756 19556
rect 18772 19612 18836 19616
rect 18772 19556 18776 19612
rect 18776 19556 18832 19612
rect 18832 19556 18836 19612
rect 18772 19552 18836 19556
rect 18852 19612 18916 19616
rect 18852 19556 18856 19612
rect 18856 19556 18912 19612
rect 18912 19556 18916 19612
rect 18852 19552 18916 19556
rect 26612 19612 26676 19616
rect 26612 19556 26616 19612
rect 26616 19556 26672 19612
rect 26672 19556 26676 19612
rect 26612 19552 26676 19556
rect 26692 19612 26756 19616
rect 26692 19556 26696 19612
rect 26696 19556 26752 19612
rect 26752 19556 26756 19612
rect 26692 19552 26756 19556
rect 26772 19612 26836 19616
rect 26772 19556 26776 19612
rect 26776 19556 26832 19612
rect 26832 19556 26836 19612
rect 26772 19552 26836 19556
rect 26852 19612 26916 19616
rect 26852 19556 26856 19612
rect 26856 19556 26912 19612
rect 26912 19556 26916 19612
rect 26852 19552 26916 19556
rect 1952 19068 2016 19072
rect 1952 19012 1956 19068
rect 1956 19012 2012 19068
rect 2012 19012 2016 19068
rect 1952 19008 2016 19012
rect 2032 19068 2096 19072
rect 2032 19012 2036 19068
rect 2036 19012 2092 19068
rect 2092 19012 2096 19068
rect 2032 19008 2096 19012
rect 2112 19068 2176 19072
rect 2112 19012 2116 19068
rect 2116 19012 2172 19068
rect 2172 19012 2176 19068
rect 2112 19008 2176 19012
rect 2192 19068 2256 19072
rect 2192 19012 2196 19068
rect 2196 19012 2252 19068
rect 2252 19012 2256 19068
rect 2192 19008 2256 19012
rect 9952 19068 10016 19072
rect 9952 19012 9956 19068
rect 9956 19012 10012 19068
rect 10012 19012 10016 19068
rect 9952 19008 10016 19012
rect 10032 19068 10096 19072
rect 10032 19012 10036 19068
rect 10036 19012 10092 19068
rect 10092 19012 10096 19068
rect 10032 19008 10096 19012
rect 10112 19068 10176 19072
rect 10112 19012 10116 19068
rect 10116 19012 10172 19068
rect 10172 19012 10176 19068
rect 10112 19008 10176 19012
rect 10192 19068 10256 19072
rect 10192 19012 10196 19068
rect 10196 19012 10252 19068
rect 10252 19012 10256 19068
rect 10192 19008 10256 19012
rect 17952 19068 18016 19072
rect 17952 19012 17956 19068
rect 17956 19012 18012 19068
rect 18012 19012 18016 19068
rect 17952 19008 18016 19012
rect 18032 19068 18096 19072
rect 18032 19012 18036 19068
rect 18036 19012 18092 19068
rect 18092 19012 18096 19068
rect 18032 19008 18096 19012
rect 18112 19068 18176 19072
rect 18112 19012 18116 19068
rect 18116 19012 18172 19068
rect 18172 19012 18176 19068
rect 18112 19008 18176 19012
rect 18192 19068 18256 19072
rect 18192 19012 18196 19068
rect 18196 19012 18252 19068
rect 18252 19012 18256 19068
rect 18192 19008 18256 19012
rect 25952 19068 26016 19072
rect 25952 19012 25956 19068
rect 25956 19012 26012 19068
rect 26012 19012 26016 19068
rect 25952 19008 26016 19012
rect 26032 19068 26096 19072
rect 26032 19012 26036 19068
rect 26036 19012 26092 19068
rect 26092 19012 26096 19068
rect 26032 19008 26096 19012
rect 26112 19068 26176 19072
rect 26112 19012 26116 19068
rect 26116 19012 26172 19068
rect 26172 19012 26176 19068
rect 26112 19008 26176 19012
rect 26192 19068 26256 19072
rect 26192 19012 26196 19068
rect 26196 19012 26252 19068
rect 26252 19012 26256 19068
rect 26192 19008 26256 19012
rect 2612 18524 2676 18528
rect 2612 18468 2616 18524
rect 2616 18468 2672 18524
rect 2672 18468 2676 18524
rect 2612 18464 2676 18468
rect 2692 18524 2756 18528
rect 2692 18468 2696 18524
rect 2696 18468 2752 18524
rect 2752 18468 2756 18524
rect 2692 18464 2756 18468
rect 2772 18524 2836 18528
rect 2772 18468 2776 18524
rect 2776 18468 2832 18524
rect 2832 18468 2836 18524
rect 2772 18464 2836 18468
rect 2852 18524 2916 18528
rect 2852 18468 2856 18524
rect 2856 18468 2912 18524
rect 2912 18468 2916 18524
rect 2852 18464 2916 18468
rect 10612 18524 10676 18528
rect 10612 18468 10616 18524
rect 10616 18468 10672 18524
rect 10672 18468 10676 18524
rect 10612 18464 10676 18468
rect 10692 18524 10756 18528
rect 10692 18468 10696 18524
rect 10696 18468 10752 18524
rect 10752 18468 10756 18524
rect 10692 18464 10756 18468
rect 10772 18524 10836 18528
rect 10772 18468 10776 18524
rect 10776 18468 10832 18524
rect 10832 18468 10836 18524
rect 10772 18464 10836 18468
rect 10852 18524 10916 18528
rect 10852 18468 10856 18524
rect 10856 18468 10912 18524
rect 10912 18468 10916 18524
rect 10852 18464 10916 18468
rect 18612 18524 18676 18528
rect 18612 18468 18616 18524
rect 18616 18468 18672 18524
rect 18672 18468 18676 18524
rect 18612 18464 18676 18468
rect 18692 18524 18756 18528
rect 18692 18468 18696 18524
rect 18696 18468 18752 18524
rect 18752 18468 18756 18524
rect 18692 18464 18756 18468
rect 18772 18524 18836 18528
rect 18772 18468 18776 18524
rect 18776 18468 18832 18524
rect 18832 18468 18836 18524
rect 18772 18464 18836 18468
rect 18852 18524 18916 18528
rect 18852 18468 18856 18524
rect 18856 18468 18912 18524
rect 18912 18468 18916 18524
rect 18852 18464 18916 18468
rect 26612 18524 26676 18528
rect 26612 18468 26616 18524
rect 26616 18468 26672 18524
rect 26672 18468 26676 18524
rect 26612 18464 26676 18468
rect 26692 18524 26756 18528
rect 26692 18468 26696 18524
rect 26696 18468 26752 18524
rect 26752 18468 26756 18524
rect 26692 18464 26756 18468
rect 26772 18524 26836 18528
rect 26772 18468 26776 18524
rect 26776 18468 26832 18524
rect 26832 18468 26836 18524
rect 26772 18464 26836 18468
rect 26852 18524 26916 18528
rect 26852 18468 26856 18524
rect 26856 18468 26912 18524
rect 26912 18468 26916 18524
rect 26852 18464 26916 18468
rect 1952 17980 2016 17984
rect 1952 17924 1956 17980
rect 1956 17924 2012 17980
rect 2012 17924 2016 17980
rect 1952 17920 2016 17924
rect 2032 17980 2096 17984
rect 2032 17924 2036 17980
rect 2036 17924 2092 17980
rect 2092 17924 2096 17980
rect 2032 17920 2096 17924
rect 2112 17980 2176 17984
rect 2112 17924 2116 17980
rect 2116 17924 2172 17980
rect 2172 17924 2176 17980
rect 2112 17920 2176 17924
rect 2192 17980 2256 17984
rect 2192 17924 2196 17980
rect 2196 17924 2252 17980
rect 2252 17924 2256 17980
rect 2192 17920 2256 17924
rect 9952 17980 10016 17984
rect 9952 17924 9956 17980
rect 9956 17924 10012 17980
rect 10012 17924 10016 17980
rect 9952 17920 10016 17924
rect 10032 17980 10096 17984
rect 10032 17924 10036 17980
rect 10036 17924 10092 17980
rect 10092 17924 10096 17980
rect 10032 17920 10096 17924
rect 10112 17980 10176 17984
rect 10112 17924 10116 17980
rect 10116 17924 10172 17980
rect 10172 17924 10176 17980
rect 10112 17920 10176 17924
rect 10192 17980 10256 17984
rect 10192 17924 10196 17980
rect 10196 17924 10252 17980
rect 10252 17924 10256 17980
rect 10192 17920 10256 17924
rect 17952 17980 18016 17984
rect 17952 17924 17956 17980
rect 17956 17924 18012 17980
rect 18012 17924 18016 17980
rect 17952 17920 18016 17924
rect 18032 17980 18096 17984
rect 18032 17924 18036 17980
rect 18036 17924 18092 17980
rect 18092 17924 18096 17980
rect 18032 17920 18096 17924
rect 18112 17980 18176 17984
rect 18112 17924 18116 17980
rect 18116 17924 18172 17980
rect 18172 17924 18176 17980
rect 18112 17920 18176 17924
rect 18192 17980 18256 17984
rect 18192 17924 18196 17980
rect 18196 17924 18252 17980
rect 18252 17924 18256 17980
rect 18192 17920 18256 17924
rect 25952 17980 26016 17984
rect 25952 17924 25956 17980
rect 25956 17924 26012 17980
rect 26012 17924 26016 17980
rect 25952 17920 26016 17924
rect 26032 17980 26096 17984
rect 26032 17924 26036 17980
rect 26036 17924 26092 17980
rect 26092 17924 26096 17980
rect 26032 17920 26096 17924
rect 26112 17980 26176 17984
rect 26112 17924 26116 17980
rect 26116 17924 26172 17980
rect 26172 17924 26176 17980
rect 26112 17920 26176 17924
rect 26192 17980 26256 17984
rect 26192 17924 26196 17980
rect 26196 17924 26252 17980
rect 26252 17924 26256 17980
rect 26192 17920 26256 17924
rect 2612 17436 2676 17440
rect 2612 17380 2616 17436
rect 2616 17380 2672 17436
rect 2672 17380 2676 17436
rect 2612 17376 2676 17380
rect 2692 17436 2756 17440
rect 2692 17380 2696 17436
rect 2696 17380 2752 17436
rect 2752 17380 2756 17436
rect 2692 17376 2756 17380
rect 2772 17436 2836 17440
rect 2772 17380 2776 17436
rect 2776 17380 2832 17436
rect 2832 17380 2836 17436
rect 2772 17376 2836 17380
rect 2852 17436 2916 17440
rect 2852 17380 2856 17436
rect 2856 17380 2912 17436
rect 2912 17380 2916 17436
rect 2852 17376 2916 17380
rect 10612 17436 10676 17440
rect 10612 17380 10616 17436
rect 10616 17380 10672 17436
rect 10672 17380 10676 17436
rect 10612 17376 10676 17380
rect 10692 17436 10756 17440
rect 10692 17380 10696 17436
rect 10696 17380 10752 17436
rect 10752 17380 10756 17436
rect 10692 17376 10756 17380
rect 10772 17436 10836 17440
rect 10772 17380 10776 17436
rect 10776 17380 10832 17436
rect 10832 17380 10836 17436
rect 10772 17376 10836 17380
rect 10852 17436 10916 17440
rect 10852 17380 10856 17436
rect 10856 17380 10912 17436
rect 10912 17380 10916 17436
rect 10852 17376 10916 17380
rect 18612 17436 18676 17440
rect 18612 17380 18616 17436
rect 18616 17380 18672 17436
rect 18672 17380 18676 17436
rect 18612 17376 18676 17380
rect 18692 17436 18756 17440
rect 18692 17380 18696 17436
rect 18696 17380 18752 17436
rect 18752 17380 18756 17436
rect 18692 17376 18756 17380
rect 18772 17436 18836 17440
rect 18772 17380 18776 17436
rect 18776 17380 18832 17436
rect 18832 17380 18836 17436
rect 18772 17376 18836 17380
rect 18852 17436 18916 17440
rect 18852 17380 18856 17436
rect 18856 17380 18912 17436
rect 18912 17380 18916 17436
rect 18852 17376 18916 17380
rect 26612 17436 26676 17440
rect 26612 17380 26616 17436
rect 26616 17380 26672 17436
rect 26672 17380 26676 17436
rect 26612 17376 26676 17380
rect 26692 17436 26756 17440
rect 26692 17380 26696 17436
rect 26696 17380 26752 17436
rect 26752 17380 26756 17436
rect 26692 17376 26756 17380
rect 26772 17436 26836 17440
rect 26772 17380 26776 17436
rect 26776 17380 26832 17436
rect 26832 17380 26836 17436
rect 26772 17376 26836 17380
rect 26852 17436 26916 17440
rect 26852 17380 26856 17436
rect 26856 17380 26912 17436
rect 26912 17380 26916 17436
rect 26852 17376 26916 17380
rect 1952 16892 2016 16896
rect 1952 16836 1956 16892
rect 1956 16836 2012 16892
rect 2012 16836 2016 16892
rect 1952 16832 2016 16836
rect 2032 16892 2096 16896
rect 2032 16836 2036 16892
rect 2036 16836 2092 16892
rect 2092 16836 2096 16892
rect 2032 16832 2096 16836
rect 2112 16892 2176 16896
rect 2112 16836 2116 16892
rect 2116 16836 2172 16892
rect 2172 16836 2176 16892
rect 2112 16832 2176 16836
rect 2192 16892 2256 16896
rect 2192 16836 2196 16892
rect 2196 16836 2252 16892
rect 2252 16836 2256 16892
rect 2192 16832 2256 16836
rect 9952 16892 10016 16896
rect 9952 16836 9956 16892
rect 9956 16836 10012 16892
rect 10012 16836 10016 16892
rect 9952 16832 10016 16836
rect 10032 16892 10096 16896
rect 10032 16836 10036 16892
rect 10036 16836 10092 16892
rect 10092 16836 10096 16892
rect 10032 16832 10096 16836
rect 10112 16892 10176 16896
rect 10112 16836 10116 16892
rect 10116 16836 10172 16892
rect 10172 16836 10176 16892
rect 10112 16832 10176 16836
rect 10192 16892 10256 16896
rect 10192 16836 10196 16892
rect 10196 16836 10252 16892
rect 10252 16836 10256 16892
rect 10192 16832 10256 16836
rect 17952 16892 18016 16896
rect 17952 16836 17956 16892
rect 17956 16836 18012 16892
rect 18012 16836 18016 16892
rect 17952 16832 18016 16836
rect 18032 16892 18096 16896
rect 18032 16836 18036 16892
rect 18036 16836 18092 16892
rect 18092 16836 18096 16892
rect 18032 16832 18096 16836
rect 18112 16892 18176 16896
rect 18112 16836 18116 16892
rect 18116 16836 18172 16892
rect 18172 16836 18176 16892
rect 18112 16832 18176 16836
rect 18192 16892 18256 16896
rect 18192 16836 18196 16892
rect 18196 16836 18252 16892
rect 18252 16836 18256 16892
rect 18192 16832 18256 16836
rect 25952 16892 26016 16896
rect 25952 16836 25956 16892
rect 25956 16836 26012 16892
rect 26012 16836 26016 16892
rect 25952 16832 26016 16836
rect 26032 16892 26096 16896
rect 26032 16836 26036 16892
rect 26036 16836 26092 16892
rect 26092 16836 26096 16892
rect 26032 16832 26096 16836
rect 26112 16892 26176 16896
rect 26112 16836 26116 16892
rect 26116 16836 26172 16892
rect 26172 16836 26176 16892
rect 26112 16832 26176 16836
rect 26192 16892 26256 16896
rect 26192 16836 26196 16892
rect 26196 16836 26252 16892
rect 26252 16836 26256 16892
rect 26192 16832 26256 16836
rect 2612 16348 2676 16352
rect 2612 16292 2616 16348
rect 2616 16292 2672 16348
rect 2672 16292 2676 16348
rect 2612 16288 2676 16292
rect 2692 16348 2756 16352
rect 2692 16292 2696 16348
rect 2696 16292 2752 16348
rect 2752 16292 2756 16348
rect 2692 16288 2756 16292
rect 2772 16348 2836 16352
rect 2772 16292 2776 16348
rect 2776 16292 2832 16348
rect 2832 16292 2836 16348
rect 2772 16288 2836 16292
rect 2852 16348 2916 16352
rect 2852 16292 2856 16348
rect 2856 16292 2912 16348
rect 2912 16292 2916 16348
rect 2852 16288 2916 16292
rect 10612 16348 10676 16352
rect 10612 16292 10616 16348
rect 10616 16292 10672 16348
rect 10672 16292 10676 16348
rect 10612 16288 10676 16292
rect 10692 16348 10756 16352
rect 10692 16292 10696 16348
rect 10696 16292 10752 16348
rect 10752 16292 10756 16348
rect 10692 16288 10756 16292
rect 10772 16348 10836 16352
rect 10772 16292 10776 16348
rect 10776 16292 10832 16348
rect 10832 16292 10836 16348
rect 10772 16288 10836 16292
rect 10852 16348 10916 16352
rect 10852 16292 10856 16348
rect 10856 16292 10912 16348
rect 10912 16292 10916 16348
rect 10852 16288 10916 16292
rect 18612 16348 18676 16352
rect 18612 16292 18616 16348
rect 18616 16292 18672 16348
rect 18672 16292 18676 16348
rect 18612 16288 18676 16292
rect 18692 16348 18756 16352
rect 18692 16292 18696 16348
rect 18696 16292 18752 16348
rect 18752 16292 18756 16348
rect 18692 16288 18756 16292
rect 18772 16348 18836 16352
rect 18772 16292 18776 16348
rect 18776 16292 18832 16348
rect 18832 16292 18836 16348
rect 18772 16288 18836 16292
rect 18852 16348 18916 16352
rect 18852 16292 18856 16348
rect 18856 16292 18912 16348
rect 18912 16292 18916 16348
rect 18852 16288 18916 16292
rect 26612 16348 26676 16352
rect 26612 16292 26616 16348
rect 26616 16292 26672 16348
rect 26672 16292 26676 16348
rect 26612 16288 26676 16292
rect 26692 16348 26756 16352
rect 26692 16292 26696 16348
rect 26696 16292 26752 16348
rect 26752 16292 26756 16348
rect 26692 16288 26756 16292
rect 26772 16348 26836 16352
rect 26772 16292 26776 16348
rect 26776 16292 26832 16348
rect 26832 16292 26836 16348
rect 26772 16288 26836 16292
rect 26852 16348 26916 16352
rect 26852 16292 26856 16348
rect 26856 16292 26912 16348
rect 26912 16292 26916 16348
rect 26852 16288 26916 16292
rect 1952 15804 2016 15808
rect 1952 15748 1956 15804
rect 1956 15748 2012 15804
rect 2012 15748 2016 15804
rect 1952 15744 2016 15748
rect 2032 15804 2096 15808
rect 2032 15748 2036 15804
rect 2036 15748 2092 15804
rect 2092 15748 2096 15804
rect 2032 15744 2096 15748
rect 2112 15804 2176 15808
rect 2112 15748 2116 15804
rect 2116 15748 2172 15804
rect 2172 15748 2176 15804
rect 2112 15744 2176 15748
rect 2192 15804 2256 15808
rect 2192 15748 2196 15804
rect 2196 15748 2252 15804
rect 2252 15748 2256 15804
rect 2192 15744 2256 15748
rect 9952 15804 10016 15808
rect 9952 15748 9956 15804
rect 9956 15748 10012 15804
rect 10012 15748 10016 15804
rect 9952 15744 10016 15748
rect 10032 15804 10096 15808
rect 10032 15748 10036 15804
rect 10036 15748 10092 15804
rect 10092 15748 10096 15804
rect 10032 15744 10096 15748
rect 10112 15804 10176 15808
rect 10112 15748 10116 15804
rect 10116 15748 10172 15804
rect 10172 15748 10176 15804
rect 10112 15744 10176 15748
rect 10192 15804 10256 15808
rect 10192 15748 10196 15804
rect 10196 15748 10252 15804
rect 10252 15748 10256 15804
rect 10192 15744 10256 15748
rect 17952 15804 18016 15808
rect 17952 15748 17956 15804
rect 17956 15748 18012 15804
rect 18012 15748 18016 15804
rect 17952 15744 18016 15748
rect 18032 15804 18096 15808
rect 18032 15748 18036 15804
rect 18036 15748 18092 15804
rect 18092 15748 18096 15804
rect 18032 15744 18096 15748
rect 18112 15804 18176 15808
rect 18112 15748 18116 15804
rect 18116 15748 18172 15804
rect 18172 15748 18176 15804
rect 18112 15744 18176 15748
rect 18192 15804 18256 15808
rect 18192 15748 18196 15804
rect 18196 15748 18252 15804
rect 18252 15748 18256 15804
rect 18192 15744 18256 15748
rect 25952 15804 26016 15808
rect 25952 15748 25956 15804
rect 25956 15748 26012 15804
rect 26012 15748 26016 15804
rect 25952 15744 26016 15748
rect 26032 15804 26096 15808
rect 26032 15748 26036 15804
rect 26036 15748 26092 15804
rect 26092 15748 26096 15804
rect 26032 15744 26096 15748
rect 26112 15804 26176 15808
rect 26112 15748 26116 15804
rect 26116 15748 26172 15804
rect 26172 15748 26176 15804
rect 26112 15744 26176 15748
rect 26192 15804 26256 15808
rect 26192 15748 26196 15804
rect 26196 15748 26252 15804
rect 26252 15748 26256 15804
rect 26192 15744 26256 15748
rect 2612 15260 2676 15264
rect 2612 15204 2616 15260
rect 2616 15204 2672 15260
rect 2672 15204 2676 15260
rect 2612 15200 2676 15204
rect 2692 15260 2756 15264
rect 2692 15204 2696 15260
rect 2696 15204 2752 15260
rect 2752 15204 2756 15260
rect 2692 15200 2756 15204
rect 2772 15260 2836 15264
rect 2772 15204 2776 15260
rect 2776 15204 2832 15260
rect 2832 15204 2836 15260
rect 2772 15200 2836 15204
rect 2852 15260 2916 15264
rect 2852 15204 2856 15260
rect 2856 15204 2912 15260
rect 2912 15204 2916 15260
rect 2852 15200 2916 15204
rect 10612 15260 10676 15264
rect 10612 15204 10616 15260
rect 10616 15204 10672 15260
rect 10672 15204 10676 15260
rect 10612 15200 10676 15204
rect 10692 15260 10756 15264
rect 10692 15204 10696 15260
rect 10696 15204 10752 15260
rect 10752 15204 10756 15260
rect 10692 15200 10756 15204
rect 10772 15260 10836 15264
rect 10772 15204 10776 15260
rect 10776 15204 10832 15260
rect 10832 15204 10836 15260
rect 10772 15200 10836 15204
rect 10852 15260 10916 15264
rect 10852 15204 10856 15260
rect 10856 15204 10912 15260
rect 10912 15204 10916 15260
rect 10852 15200 10916 15204
rect 18612 15260 18676 15264
rect 18612 15204 18616 15260
rect 18616 15204 18672 15260
rect 18672 15204 18676 15260
rect 18612 15200 18676 15204
rect 18692 15260 18756 15264
rect 18692 15204 18696 15260
rect 18696 15204 18752 15260
rect 18752 15204 18756 15260
rect 18692 15200 18756 15204
rect 18772 15260 18836 15264
rect 18772 15204 18776 15260
rect 18776 15204 18832 15260
rect 18832 15204 18836 15260
rect 18772 15200 18836 15204
rect 18852 15260 18916 15264
rect 18852 15204 18856 15260
rect 18856 15204 18912 15260
rect 18912 15204 18916 15260
rect 18852 15200 18916 15204
rect 26612 15260 26676 15264
rect 26612 15204 26616 15260
rect 26616 15204 26672 15260
rect 26672 15204 26676 15260
rect 26612 15200 26676 15204
rect 26692 15260 26756 15264
rect 26692 15204 26696 15260
rect 26696 15204 26752 15260
rect 26752 15204 26756 15260
rect 26692 15200 26756 15204
rect 26772 15260 26836 15264
rect 26772 15204 26776 15260
rect 26776 15204 26832 15260
rect 26832 15204 26836 15260
rect 26772 15200 26836 15204
rect 26852 15260 26916 15264
rect 26852 15204 26856 15260
rect 26856 15204 26912 15260
rect 26912 15204 26916 15260
rect 26852 15200 26916 15204
rect 1952 14716 2016 14720
rect 1952 14660 1956 14716
rect 1956 14660 2012 14716
rect 2012 14660 2016 14716
rect 1952 14656 2016 14660
rect 2032 14716 2096 14720
rect 2032 14660 2036 14716
rect 2036 14660 2092 14716
rect 2092 14660 2096 14716
rect 2032 14656 2096 14660
rect 2112 14716 2176 14720
rect 2112 14660 2116 14716
rect 2116 14660 2172 14716
rect 2172 14660 2176 14716
rect 2112 14656 2176 14660
rect 2192 14716 2256 14720
rect 2192 14660 2196 14716
rect 2196 14660 2252 14716
rect 2252 14660 2256 14716
rect 2192 14656 2256 14660
rect 9952 14716 10016 14720
rect 9952 14660 9956 14716
rect 9956 14660 10012 14716
rect 10012 14660 10016 14716
rect 9952 14656 10016 14660
rect 10032 14716 10096 14720
rect 10032 14660 10036 14716
rect 10036 14660 10092 14716
rect 10092 14660 10096 14716
rect 10032 14656 10096 14660
rect 10112 14716 10176 14720
rect 10112 14660 10116 14716
rect 10116 14660 10172 14716
rect 10172 14660 10176 14716
rect 10112 14656 10176 14660
rect 10192 14716 10256 14720
rect 10192 14660 10196 14716
rect 10196 14660 10252 14716
rect 10252 14660 10256 14716
rect 10192 14656 10256 14660
rect 17952 14716 18016 14720
rect 17952 14660 17956 14716
rect 17956 14660 18012 14716
rect 18012 14660 18016 14716
rect 17952 14656 18016 14660
rect 18032 14716 18096 14720
rect 18032 14660 18036 14716
rect 18036 14660 18092 14716
rect 18092 14660 18096 14716
rect 18032 14656 18096 14660
rect 18112 14716 18176 14720
rect 18112 14660 18116 14716
rect 18116 14660 18172 14716
rect 18172 14660 18176 14716
rect 18112 14656 18176 14660
rect 18192 14716 18256 14720
rect 18192 14660 18196 14716
rect 18196 14660 18252 14716
rect 18252 14660 18256 14716
rect 18192 14656 18256 14660
rect 25952 14716 26016 14720
rect 25952 14660 25956 14716
rect 25956 14660 26012 14716
rect 26012 14660 26016 14716
rect 25952 14656 26016 14660
rect 26032 14716 26096 14720
rect 26032 14660 26036 14716
rect 26036 14660 26092 14716
rect 26092 14660 26096 14716
rect 26032 14656 26096 14660
rect 26112 14716 26176 14720
rect 26112 14660 26116 14716
rect 26116 14660 26172 14716
rect 26172 14660 26176 14716
rect 26112 14656 26176 14660
rect 26192 14716 26256 14720
rect 26192 14660 26196 14716
rect 26196 14660 26252 14716
rect 26252 14660 26256 14716
rect 26192 14656 26256 14660
rect 2612 14172 2676 14176
rect 2612 14116 2616 14172
rect 2616 14116 2672 14172
rect 2672 14116 2676 14172
rect 2612 14112 2676 14116
rect 2692 14172 2756 14176
rect 2692 14116 2696 14172
rect 2696 14116 2752 14172
rect 2752 14116 2756 14172
rect 2692 14112 2756 14116
rect 2772 14172 2836 14176
rect 2772 14116 2776 14172
rect 2776 14116 2832 14172
rect 2832 14116 2836 14172
rect 2772 14112 2836 14116
rect 2852 14172 2916 14176
rect 2852 14116 2856 14172
rect 2856 14116 2912 14172
rect 2912 14116 2916 14172
rect 2852 14112 2916 14116
rect 10612 14172 10676 14176
rect 10612 14116 10616 14172
rect 10616 14116 10672 14172
rect 10672 14116 10676 14172
rect 10612 14112 10676 14116
rect 10692 14172 10756 14176
rect 10692 14116 10696 14172
rect 10696 14116 10752 14172
rect 10752 14116 10756 14172
rect 10692 14112 10756 14116
rect 10772 14172 10836 14176
rect 10772 14116 10776 14172
rect 10776 14116 10832 14172
rect 10832 14116 10836 14172
rect 10772 14112 10836 14116
rect 10852 14172 10916 14176
rect 10852 14116 10856 14172
rect 10856 14116 10912 14172
rect 10912 14116 10916 14172
rect 10852 14112 10916 14116
rect 18612 14172 18676 14176
rect 18612 14116 18616 14172
rect 18616 14116 18672 14172
rect 18672 14116 18676 14172
rect 18612 14112 18676 14116
rect 18692 14172 18756 14176
rect 18692 14116 18696 14172
rect 18696 14116 18752 14172
rect 18752 14116 18756 14172
rect 18692 14112 18756 14116
rect 18772 14172 18836 14176
rect 18772 14116 18776 14172
rect 18776 14116 18832 14172
rect 18832 14116 18836 14172
rect 18772 14112 18836 14116
rect 18852 14172 18916 14176
rect 18852 14116 18856 14172
rect 18856 14116 18912 14172
rect 18912 14116 18916 14172
rect 18852 14112 18916 14116
rect 26612 14172 26676 14176
rect 26612 14116 26616 14172
rect 26616 14116 26672 14172
rect 26672 14116 26676 14172
rect 26612 14112 26676 14116
rect 26692 14172 26756 14176
rect 26692 14116 26696 14172
rect 26696 14116 26752 14172
rect 26752 14116 26756 14172
rect 26692 14112 26756 14116
rect 26772 14172 26836 14176
rect 26772 14116 26776 14172
rect 26776 14116 26832 14172
rect 26832 14116 26836 14172
rect 26772 14112 26836 14116
rect 26852 14172 26916 14176
rect 26852 14116 26856 14172
rect 26856 14116 26912 14172
rect 26912 14116 26916 14172
rect 26852 14112 26916 14116
rect 1952 13628 2016 13632
rect 1952 13572 1956 13628
rect 1956 13572 2012 13628
rect 2012 13572 2016 13628
rect 1952 13568 2016 13572
rect 2032 13628 2096 13632
rect 2032 13572 2036 13628
rect 2036 13572 2092 13628
rect 2092 13572 2096 13628
rect 2032 13568 2096 13572
rect 2112 13628 2176 13632
rect 2112 13572 2116 13628
rect 2116 13572 2172 13628
rect 2172 13572 2176 13628
rect 2112 13568 2176 13572
rect 2192 13628 2256 13632
rect 2192 13572 2196 13628
rect 2196 13572 2252 13628
rect 2252 13572 2256 13628
rect 2192 13568 2256 13572
rect 9952 13628 10016 13632
rect 9952 13572 9956 13628
rect 9956 13572 10012 13628
rect 10012 13572 10016 13628
rect 9952 13568 10016 13572
rect 10032 13628 10096 13632
rect 10032 13572 10036 13628
rect 10036 13572 10092 13628
rect 10092 13572 10096 13628
rect 10032 13568 10096 13572
rect 10112 13628 10176 13632
rect 10112 13572 10116 13628
rect 10116 13572 10172 13628
rect 10172 13572 10176 13628
rect 10112 13568 10176 13572
rect 10192 13628 10256 13632
rect 10192 13572 10196 13628
rect 10196 13572 10252 13628
rect 10252 13572 10256 13628
rect 10192 13568 10256 13572
rect 17952 13628 18016 13632
rect 17952 13572 17956 13628
rect 17956 13572 18012 13628
rect 18012 13572 18016 13628
rect 17952 13568 18016 13572
rect 18032 13628 18096 13632
rect 18032 13572 18036 13628
rect 18036 13572 18092 13628
rect 18092 13572 18096 13628
rect 18032 13568 18096 13572
rect 18112 13628 18176 13632
rect 18112 13572 18116 13628
rect 18116 13572 18172 13628
rect 18172 13572 18176 13628
rect 18112 13568 18176 13572
rect 18192 13628 18256 13632
rect 18192 13572 18196 13628
rect 18196 13572 18252 13628
rect 18252 13572 18256 13628
rect 18192 13568 18256 13572
rect 25952 13628 26016 13632
rect 25952 13572 25956 13628
rect 25956 13572 26012 13628
rect 26012 13572 26016 13628
rect 25952 13568 26016 13572
rect 26032 13628 26096 13632
rect 26032 13572 26036 13628
rect 26036 13572 26092 13628
rect 26092 13572 26096 13628
rect 26032 13568 26096 13572
rect 26112 13628 26176 13632
rect 26112 13572 26116 13628
rect 26116 13572 26172 13628
rect 26172 13572 26176 13628
rect 26112 13568 26176 13572
rect 26192 13628 26256 13632
rect 26192 13572 26196 13628
rect 26196 13572 26252 13628
rect 26252 13572 26256 13628
rect 26192 13568 26256 13572
rect 2612 13084 2676 13088
rect 2612 13028 2616 13084
rect 2616 13028 2672 13084
rect 2672 13028 2676 13084
rect 2612 13024 2676 13028
rect 2692 13084 2756 13088
rect 2692 13028 2696 13084
rect 2696 13028 2752 13084
rect 2752 13028 2756 13084
rect 2692 13024 2756 13028
rect 2772 13084 2836 13088
rect 2772 13028 2776 13084
rect 2776 13028 2832 13084
rect 2832 13028 2836 13084
rect 2772 13024 2836 13028
rect 2852 13084 2916 13088
rect 2852 13028 2856 13084
rect 2856 13028 2912 13084
rect 2912 13028 2916 13084
rect 2852 13024 2916 13028
rect 10612 13084 10676 13088
rect 10612 13028 10616 13084
rect 10616 13028 10672 13084
rect 10672 13028 10676 13084
rect 10612 13024 10676 13028
rect 10692 13084 10756 13088
rect 10692 13028 10696 13084
rect 10696 13028 10752 13084
rect 10752 13028 10756 13084
rect 10692 13024 10756 13028
rect 10772 13084 10836 13088
rect 10772 13028 10776 13084
rect 10776 13028 10832 13084
rect 10832 13028 10836 13084
rect 10772 13024 10836 13028
rect 10852 13084 10916 13088
rect 10852 13028 10856 13084
rect 10856 13028 10912 13084
rect 10912 13028 10916 13084
rect 10852 13024 10916 13028
rect 18612 13084 18676 13088
rect 18612 13028 18616 13084
rect 18616 13028 18672 13084
rect 18672 13028 18676 13084
rect 18612 13024 18676 13028
rect 18692 13084 18756 13088
rect 18692 13028 18696 13084
rect 18696 13028 18752 13084
rect 18752 13028 18756 13084
rect 18692 13024 18756 13028
rect 18772 13084 18836 13088
rect 18772 13028 18776 13084
rect 18776 13028 18832 13084
rect 18832 13028 18836 13084
rect 18772 13024 18836 13028
rect 18852 13084 18916 13088
rect 18852 13028 18856 13084
rect 18856 13028 18912 13084
rect 18912 13028 18916 13084
rect 18852 13024 18916 13028
rect 26612 13084 26676 13088
rect 26612 13028 26616 13084
rect 26616 13028 26672 13084
rect 26672 13028 26676 13084
rect 26612 13024 26676 13028
rect 26692 13084 26756 13088
rect 26692 13028 26696 13084
rect 26696 13028 26752 13084
rect 26752 13028 26756 13084
rect 26692 13024 26756 13028
rect 26772 13084 26836 13088
rect 26772 13028 26776 13084
rect 26776 13028 26832 13084
rect 26832 13028 26836 13084
rect 26772 13024 26836 13028
rect 26852 13084 26916 13088
rect 26852 13028 26856 13084
rect 26856 13028 26912 13084
rect 26912 13028 26916 13084
rect 26852 13024 26916 13028
rect 1952 12540 2016 12544
rect 1952 12484 1956 12540
rect 1956 12484 2012 12540
rect 2012 12484 2016 12540
rect 1952 12480 2016 12484
rect 2032 12540 2096 12544
rect 2032 12484 2036 12540
rect 2036 12484 2092 12540
rect 2092 12484 2096 12540
rect 2032 12480 2096 12484
rect 2112 12540 2176 12544
rect 2112 12484 2116 12540
rect 2116 12484 2172 12540
rect 2172 12484 2176 12540
rect 2112 12480 2176 12484
rect 2192 12540 2256 12544
rect 2192 12484 2196 12540
rect 2196 12484 2252 12540
rect 2252 12484 2256 12540
rect 2192 12480 2256 12484
rect 9952 12540 10016 12544
rect 9952 12484 9956 12540
rect 9956 12484 10012 12540
rect 10012 12484 10016 12540
rect 9952 12480 10016 12484
rect 10032 12540 10096 12544
rect 10032 12484 10036 12540
rect 10036 12484 10092 12540
rect 10092 12484 10096 12540
rect 10032 12480 10096 12484
rect 10112 12540 10176 12544
rect 10112 12484 10116 12540
rect 10116 12484 10172 12540
rect 10172 12484 10176 12540
rect 10112 12480 10176 12484
rect 10192 12540 10256 12544
rect 10192 12484 10196 12540
rect 10196 12484 10252 12540
rect 10252 12484 10256 12540
rect 10192 12480 10256 12484
rect 17952 12540 18016 12544
rect 17952 12484 17956 12540
rect 17956 12484 18012 12540
rect 18012 12484 18016 12540
rect 17952 12480 18016 12484
rect 18032 12540 18096 12544
rect 18032 12484 18036 12540
rect 18036 12484 18092 12540
rect 18092 12484 18096 12540
rect 18032 12480 18096 12484
rect 18112 12540 18176 12544
rect 18112 12484 18116 12540
rect 18116 12484 18172 12540
rect 18172 12484 18176 12540
rect 18112 12480 18176 12484
rect 18192 12540 18256 12544
rect 18192 12484 18196 12540
rect 18196 12484 18252 12540
rect 18252 12484 18256 12540
rect 18192 12480 18256 12484
rect 25952 12540 26016 12544
rect 25952 12484 25956 12540
rect 25956 12484 26012 12540
rect 26012 12484 26016 12540
rect 25952 12480 26016 12484
rect 26032 12540 26096 12544
rect 26032 12484 26036 12540
rect 26036 12484 26092 12540
rect 26092 12484 26096 12540
rect 26032 12480 26096 12484
rect 26112 12540 26176 12544
rect 26112 12484 26116 12540
rect 26116 12484 26172 12540
rect 26172 12484 26176 12540
rect 26112 12480 26176 12484
rect 26192 12540 26256 12544
rect 26192 12484 26196 12540
rect 26196 12484 26252 12540
rect 26252 12484 26256 12540
rect 26192 12480 26256 12484
rect 2612 11996 2676 12000
rect 2612 11940 2616 11996
rect 2616 11940 2672 11996
rect 2672 11940 2676 11996
rect 2612 11936 2676 11940
rect 2692 11996 2756 12000
rect 2692 11940 2696 11996
rect 2696 11940 2752 11996
rect 2752 11940 2756 11996
rect 2692 11936 2756 11940
rect 2772 11996 2836 12000
rect 2772 11940 2776 11996
rect 2776 11940 2832 11996
rect 2832 11940 2836 11996
rect 2772 11936 2836 11940
rect 2852 11996 2916 12000
rect 2852 11940 2856 11996
rect 2856 11940 2912 11996
rect 2912 11940 2916 11996
rect 2852 11936 2916 11940
rect 10612 11996 10676 12000
rect 10612 11940 10616 11996
rect 10616 11940 10672 11996
rect 10672 11940 10676 11996
rect 10612 11936 10676 11940
rect 10692 11996 10756 12000
rect 10692 11940 10696 11996
rect 10696 11940 10752 11996
rect 10752 11940 10756 11996
rect 10692 11936 10756 11940
rect 10772 11996 10836 12000
rect 10772 11940 10776 11996
rect 10776 11940 10832 11996
rect 10832 11940 10836 11996
rect 10772 11936 10836 11940
rect 10852 11996 10916 12000
rect 10852 11940 10856 11996
rect 10856 11940 10912 11996
rect 10912 11940 10916 11996
rect 10852 11936 10916 11940
rect 18612 11996 18676 12000
rect 18612 11940 18616 11996
rect 18616 11940 18672 11996
rect 18672 11940 18676 11996
rect 18612 11936 18676 11940
rect 18692 11996 18756 12000
rect 18692 11940 18696 11996
rect 18696 11940 18752 11996
rect 18752 11940 18756 11996
rect 18692 11936 18756 11940
rect 18772 11996 18836 12000
rect 18772 11940 18776 11996
rect 18776 11940 18832 11996
rect 18832 11940 18836 11996
rect 18772 11936 18836 11940
rect 18852 11996 18916 12000
rect 18852 11940 18856 11996
rect 18856 11940 18912 11996
rect 18912 11940 18916 11996
rect 18852 11936 18916 11940
rect 26612 11996 26676 12000
rect 26612 11940 26616 11996
rect 26616 11940 26672 11996
rect 26672 11940 26676 11996
rect 26612 11936 26676 11940
rect 26692 11996 26756 12000
rect 26692 11940 26696 11996
rect 26696 11940 26752 11996
rect 26752 11940 26756 11996
rect 26692 11936 26756 11940
rect 26772 11996 26836 12000
rect 26772 11940 26776 11996
rect 26776 11940 26832 11996
rect 26832 11940 26836 11996
rect 26772 11936 26836 11940
rect 26852 11996 26916 12000
rect 26852 11940 26856 11996
rect 26856 11940 26912 11996
rect 26912 11940 26916 11996
rect 26852 11936 26916 11940
rect 1952 11452 2016 11456
rect 1952 11396 1956 11452
rect 1956 11396 2012 11452
rect 2012 11396 2016 11452
rect 1952 11392 2016 11396
rect 2032 11452 2096 11456
rect 2032 11396 2036 11452
rect 2036 11396 2092 11452
rect 2092 11396 2096 11452
rect 2032 11392 2096 11396
rect 2112 11452 2176 11456
rect 2112 11396 2116 11452
rect 2116 11396 2172 11452
rect 2172 11396 2176 11452
rect 2112 11392 2176 11396
rect 2192 11452 2256 11456
rect 2192 11396 2196 11452
rect 2196 11396 2252 11452
rect 2252 11396 2256 11452
rect 2192 11392 2256 11396
rect 9952 11452 10016 11456
rect 9952 11396 9956 11452
rect 9956 11396 10012 11452
rect 10012 11396 10016 11452
rect 9952 11392 10016 11396
rect 10032 11452 10096 11456
rect 10032 11396 10036 11452
rect 10036 11396 10092 11452
rect 10092 11396 10096 11452
rect 10032 11392 10096 11396
rect 10112 11452 10176 11456
rect 10112 11396 10116 11452
rect 10116 11396 10172 11452
rect 10172 11396 10176 11452
rect 10112 11392 10176 11396
rect 10192 11452 10256 11456
rect 10192 11396 10196 11452
rect 10196 11396 10252 11452
rect 10252 11396 10256 11452
rect 10192 11392 10256 11396
rect 17952 11452 18016 11456
rect 17952 11396 17956 11452
rect 17956 11396 18012 11452
rect 18012 11396 18016 11452
rect 17952 11392 18016 11396
rect 18032 11452 18096 11456
rect 18032 11396 18036 11452
rect 18036 11396 18092 11452
rect 18092 11396 18096 11452
rect 18032 11392 18096 11396
rect 18112 11452 18176 11456
rect 18112 11396 18116 11452
rect 18116 11396 18172 11452
rect 18172 11396 18176 11452
rect 18112 11392 18176 11396
rect 18192 11452 18256 11456
rect 18192 11396 18196 11452
rect 18196 11396 18252 11452
rect 18252 11396 18256 11452
rect 18192 11392 18256 11396
rect 25952 11452 26016 11456
rect 25952 11396 25956 11452
rect 25956 11396 26012 11452
rect 26012 11396 26016 11452
rect 25952 11392 26016 11396
rect 26032 11452 26096 11456
rect 26032 11396 26036 11452
rect 26036 11396 26092 11452
rect 26092 11396 26096 11452
rect 26032 11392 26096 11396
rect 26112 11452 26176 11456
rect 26112 11396 26116 11452
rect 26116 11396 26172 11452
rect 26172 11396 26176 11452
rect 26112 11392 26176 11396
rect 26192 11452 26256 11456
rect 26192 11396 26196 11452
rect 26196 11396 26252 11452
rect 26252 11396 26256 11452
rect 26192 11392 26256 11396
rect 2612 10908 2676 10912
rect 2612 10852 2616 10908
rect 2616 10852 2672 10908
rect 2672 10852 2676 10908
rect 2612 10848 2676 10852
rect 2692 10908 2756 10912
rect 2692 10852 2696 10908
rect 2696 10852 2752 10908
rect 2752 10852 2756 10908
rect 2692 10848 2756 10852
rect 2772 10908 2836 10912
rect 2772 10852 2776 10908
rect 2776 10852 2832 10908
rect 2832 10852 2836 10908
rect 2772 10848 2836 10852
rect 2852 10908 2916 10912
rect 2852 10852 2856 10908
rect 2856 10852 2912 10908
rect 2912 10852 2916 10908
rect 2852 10848 2916 10852
rect 10612 10908 10676 10912
rect 10612 10852 10616 10908
rect 10616 10852 10672 10908
rect 10672 10852 10676 10908
rect 10612 10848 10676 10852
rect 10692 10908 10756 10912
rect 10692 10852 10696 10908
rect 10696 10852 10752 10908
rect 10752 10852 10756 10908
rect 10692 10848 10756 10852
rect 10772 10908 10836 10912
rect 10772 10852 10776 10908
rect 10776 10852 10832 10908
rect 10832 10852 10836 10908
rect 10772 10848 10836 10852
rect 10852 10908 10916 10912
rect 10852 10852 10856 10908
rect 10856 10852 10912 10908
rect 10912 10852 10916 10908
rect 10852 10848 10916 10852
rect 18612 10908 18676 10912
rect 18612 10852 18616 10908
rect 18616 10852 18672 10908
rect 18672 10852 18676 10908
rect 18612 10848 18676 10852
rect 18692 10908 18756 10912
rect 18692 10852 18696 10908
rect 18696 10852 18752 10908
rect 18752 10852 18756 10908
rect 18692 10848 18756 10852
rect 18772 10908 18836 10912
rect 18772 10852 18776 10908
rect 18776 10852 18832 10908
rect 18832 10852 18836 10908
rect 18772 10848 18836 10852
rect 18852 10908 18916 10912
rect 18852 10852 18856 10908
rect 18856 10852 18912 10908
rect 18912 10852 18916 10908
rect 18852 10848 18916 10852
rect 26612 10908 26676 10912
rect 26612 10852 26616 10908
rect 26616 10852 26672 10908
rect 26672 10852 26676 10908
rect 26612 10848 26676 10852
rect 26692 10908 26756 10912
rect 26692 10852 26696 10908
rect 26696 10852 26752 10908
rect 26752 10852 26756 10908
rect 26692 10848 26756 10852
rect 26772 10908 26836 10912
rect 26772 10852 26776 10908
rect 26776 10852 26832 10908
rect 26832 10852 26836 10908
rect 26772 10848 26836 10852
rect 26852 10908 26916 10912
rect 26852 10852 26856 10908
rect 26856 10852 26912 10908
rect 26912 10852 26916 10908
rect 26852 10848 26916 10852
rect 1952 10364 2016 10368
rect 1952 10308 1956 10364
rect 1956 10308 2012 10364
rect 2012 10308 2016 10364
rect 1952 10304 2016 10308
rect 2032 10364 2096 10368
rect 2032 10308 2036 10364
rect 2036 10308 2092 10364
rect 2092 10308 2096 10364
rect 2032 10304 2096 10308
rect 2112 10364 2176 10368
rect 2112 10308 2116 10364
rect 2116 10308 2172 10364
rect 2172 10308 2176 10364
rect 2112 10304 2176 10308
rect 2192 10364 2256 10368
rect 2192 10308 2196 10364
rect 2196 10308 2252 10364
rect 2252 10308 2256 10364
rect 2192 10304 2256 10308
rect 9952 10364 10016 10368
rect 9952 10308 9956 10364
rect 9956 10308 10012 10364
rect 10012 10308 10016 10364
rect 9952 10304 10016 10308
rect 10032 10364 10096 10368
rect 10032 10308 10036 10364
rect 10036 10308 10092 10364
rect 10092 10308 10096 10364
rect 10032 10304 10096 10308
rect 10112 10364 10176 10368
rect 10112 10308 10116 10364
rect 10116 10308 10172 10364
rect 10172 10308 10176 10364
rect 10112 10304 10176 10308
rect 10192 10364 10256 10368
rect 10192 10308 10196 10364
rect 10196 10308 10252 10364
rect 10252 10308 10256 10364
rect 10192 10304 10256 10308
rect 17952 10364 18016 10368
rect 17952 10308 17956 10364
rect 17956 10308 18012 10364
rect 18012 10308 18016 10364
rect 17952 10304 18016 10308
rect 18032 10364 18096 10368
rect 18032 10308 18036 10364
rect 18036 10308 18092 10364
rect 18092 10308 18096 10364
rect 18032 10304 18096 10308
rect 18112 10364 18176 10368
rect 18112 10308 18116 10364
rect 18116 10308 18172 10364
rect 18172 10308 18176 10364
rect 18112 10304 18176 10308
rect 18192 10364 18256 10368
rect 18192 10308 18196 10364
rect 18196 10308 18252 10364
rect 18252 10308 18256 10364
rect 18192 10304 18256 10308
rect 25952 10364 26016 10368
rect 25952 10308 25956 10364
rect 25956 10308 26012 10364
rect 26012 10308 26016 10364
rect 25952 10304 26016 10308
rect 26032 10364 26096 10368
rect 26032 10308 26036 10364
rect 26036 10308 26092 10364
rect 26092 10308 26096 10364
rect 26032 10304 26096 10308
rect 26112 10364 26176 10368
rect 26112 10308 26116 10364
rect 26116 10308 26172 10364
rect 26172 10308 26176 10364
rect 26112 10304 26176 10308
rect 26192 10364 26256 10368
rect 26192 10308 26196 10364
rect 26196 10308 26252 10364
rect 26252 10308 26256 10364
rect 26192 10304 26256 10308
rect 2612 9820 2676 9824
rect 2612 9764 2616 9820
rect 2616 9764 2672 9820
rect 2672 9764 2676 9820
rect 2612 9760 2676 9764
rect 2692 9820 2756 9824
rect 2692 9764 2696 9820
rect 2696 9764 2752 9820
rect 2752 9764 2756 9820
rect 2692 9760 2756 9764
rect 2772 9820 2836 9824
rect 2772 9764 2776 9820
rect 2776 9764 2832 9820
rect 2832 9764 2836 9820
rect 2772 9760 2836 9764
rect 2852 9820 2916 9824
rect 2852 9764 2856 9820
rect 2856 9764 2912 9820
rect 2912 9764 2916 9820
rect 2852 9760 2916 9764
rect 10612 9820 10676 9824
rect 10612 9764 10616 9820
rect 10616 9764 10672 9820
rect 10672 9764 10676 9820
rect 10612 9760 10676 9764
rect 10692 9820 10756 9824
rect 10692 9764 10696 9820
rect 10696 9764 10752 9820
rect 10752 9764 10756 9820
rect 10692 9760 10756 9764
rect 10772 9820 10836 9824
rect 10772 9764 10776 9820
rect 10776 9764 10832 9820
rect 10832 9764 10836 9820
rect 10772 9760 10836 9764
rect 10852 9820 10916 9824
rect 10852 9764 10856 9820
rect 10856 9764 10912 9820
rect 10912 9764 10916 9820
rect 10852 9760 10916 9764
rect 18612 9820 18676 9824
rect 18612 9764 18616 9820
rect 18616 9764 18672 9820
rect 18672 9764 18676 9820
rect 18612 9760 18676 9764
rect 18692 9820 18756 9824
rect 18692 9764 18696 9820
rect 18696 9764 18752 9820
rect 18752 9764 18756 9820
rect 18692 9760 18756 9764
rect 18772 9820 18836 9824
rect 18772 9764 18776 9820
rect 18776 9764 18832 9820
rect 18832 9764 18836 9820
rect 18772 9760 18836 9764
rect 18852 9820 18916 9824
rect 18852 9764 18856 9820
rect 18856 9764 18912 9820
rect 18912 9764 18916 9820
rect 18852 9760 18916 9764
rect 26612 9820 26676 9824
rect 26612 9764 26616 9820
rect 26616 9764 26672 9820
rect 26672 9764 26676 9820
rect 26612 9760 26676 9764
rect 26692 9820 26756 9824
rect 26692 9764 26696 9820
rect 26696 9764 26752 9820
rect 26752 9764 26756 9820
rect 26692 9760 26756 9764
rect 26772 9820 26836 9824
rect 26772 9764 26776 9820
rect 26776 9764 26832 9820
rect 26832 9764 26836 9820
rect 26772 9760 26836 9764
rect 26852 9820 26916 9824
rect 26852 9764 26856 9820
rect 26856 9764 26912 9820
rect 26912 9764 26916 9820
rect 26852 9760 26916 9764
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 9952 9276 10016 9280
rect 9952 9220 9956 9276
rect 9956 9220 10012 9276
rect 10012 9220 10016 9276
rect 9952 9216 10016 9220
rect 10032 9276 10096 9280
rect 10032 9220 10036 9276
rect 10036 9220 10092 9276
rect 10092 9220 10096 9276
rect 10032 9216 10096 9220
rect 10112 9276 10176 9280
rect 10112 9220 10116 9276
rect 10116 9220 10172 9276
rect 10172 9220 10176 9276
rect 10112 9216 10176 9220
rect 10192 9276 10256 9280
rect 10192 9220 10196 9276
rect 10196 9220 10252 9276
rect 10252 9220 10256 9276
rect 10192 9216 10256 9220
rect 17952 9276 18016 9280
rect 17952 9220 17956 9276
rect 17956 9220 18012 9276
rect 18012 9220 18016 9276
rect 17952 9216 18016 9220
rect 18032 9276 18096 9280
rect 18032 9220 18036 9276
rect 18036 9220 18092 9276
rect 18092 9220 18096 9276
rect 18032 9216 18096 9220
rect 18112 9276 18176 9280
rect 18112 9220 18116 9276
rect 18116 9220 18172 9276
rect 18172 9220 18176 9276
rect 18112 9216 18176 9220
rect 18192 9276 18256 9280
rect 18192 9220 18196 9276
rect 18196 9220 18252 9276
rect 18252 9220 18256 9276
rect 18192 9216 18256 9220
rect 25952 9276 26016 9280
rect 25952 9220 25956 9276
rect 25956 9220 26012 9276
rect 26012 9220 26016 9276
rect 25952 9216 26016 9220
rect 26032 9276 26096 9280
rect 26032 9220 26036 9276
rect 26036 9220 26092 9276
rect 26092 9220 26096 9276
rect 26032 9216 26096 9220
rect 26112 9276 26176 9280
rect 26112 9220 26116 9276
rect 26116 9220 26172 9276
rect 26172 9220 26176 9276
rect 26112 9216 26176 9220
rect 26192 9276 26256 9280
rect 26192 9220 26196 9276
rect 26196 9220 26252 9276
rect 26252 9220 26256 9276
rect 26192 9216 26256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 10612 8732 10676 8736
rect 10612 8676 10616 8732
rect 10616 8676 10672 8732
rect 10672 8676 10676 8732
rect 10612 8672 10676 8676
rect 10692 8732 10756 8736
rect 10692 8676 10696 8732
rect 10696 8676 10752 8732
rect 10752 8676 10756 8732
rect 10692 8672 10756 8676
rect 10772 8732 10836 8736
rect 10772 8676 10776 8732
rect 10776 8676 10832 8732
rect 10832 8676 10836 8732
rect 10772 8672 10836 8676
rect 10852 8732 10916 8736
rect 10852 8676 10856 8732
rect 10856 8676 10912 8732
rect 10912 8676 10916 8732
rect 10852 8672 10916 8676
rect 18612 8732 18676 8736
rect 18612 8676 18616 8732
rect 18616 8676 18672 8732
rect 18672 8676 18676 8732
rect 18612 8672 18676 8676
rect 18692 8732 18756 8736
rect 18692 8676 18696 8732
rect 18696 8676 18752 8732
rect 18752 8676 18756 8732
rect 18692 8672 18756 8676
rect 18772 8732 18836 8736
rect 18772 8676 18776 8732
rect 18776 8676 18832 8732
rect 18832 8676 18836 8732
rect 18772 8672 18836 8676
rect 18852 8732 18916 8736
rect 18852 8676 18856 8732
rect 18856 8676 18912 8732
rect 18912 8676 18916 8732
rect 18852 8672 18916 8676
rect 26612 8732 26676 8736
rect 26612 8676 26616 8732
rect 26616 8676 26672 8732
rect 26672 8676 26676 8732
rect 26612 8672 26676 8676
rect 26692 8732 26756 8736
rect 26692 8676 26696 8732
rect 26696 8676 26752 8732
rect 26752 8676 26756 8732
rect 26692 8672 26756 8676
rect 26772 8732 26836 8736
rect 26772 8676 26776 8732
rect 26776 8676 26832 8732
rect 26832 8676 26836 8732
rect 26772 8672 26836 8676
rect 26852 8732 26916 8736
rect 26852 8676 26856 8732
rect 26856 8676 26912 8732
rect 26912 8676 26916 8732
rect 26852 8672 26916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 9952 8188 10016 8192
rect 9952 8132 9956 8188
rect 9956 8132 10012 8188
rect 10012 8132 10016 8188
rect 9952 8128 10016 8132
rect 10032 8188 10096 8192
rect 10032 8132 10036 8188
rect 10036 8132 10092 8188
rect 10092 8132 10096 8188
rect 10032 8128 10096 8132
rect 10112 8188 10176 8192
rect 10112 8132 10116 8188
rect 10116 8132 10172 8188
rect 10172 8132 10176 8188
rect 10112 8128 10176 8132
rect 10192 8188 10256 8192
rect 10192 8132 10196 8188
rect 10196 8132 10252 8188
rect 10252 8132 10256 8188
rect 10192 8128 10256 8132
rect 17952 8188 18016 8192
rect 17952 8132 17956 8188
rect 17956 8132 18012 8188
rect 18012 8132 18016 8188
rect 17952 8128 18016 8132
rect 18032 8188 18096 8192
rect 18032 8132 18036 8188
rect 18036 8132 18092 8188
rect 18092 8132 18096 8188
rect 18032 8128 18096 8132
rect 18112 8188 18176 8192
rect 18112 8132 18116 8188
rect 18116 8132 18172 8188
rect 18172 8132 18176 8188
rect 18112 8128 18176 8132
rect 18192 8188 18256 8192
rect 18192 8132 18196 8188
rect 18196 8132 18252 8188
rect 18252 8132 18256 8188
rect 18192 8128 18256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 10612 7644 10676 7648
rect 10612 7588 10616 7644
rect 10616 7588 10672 7644
rect 10672 7588 10676 7644
rect 10612 7584 10676 7588
rect 10692 7644 10756 7648
rect 10692 7588 10696 7644
rect 10696 7588 10752 7644
rect 10752 7588 10756 7644
rect 10692 7584 10756 7588
rect 10772 7644 10836 7648
rect 10772 7588 10776 7644
rect 10776 7588 10832 7644
rect 10832 7588 10836 7644
rect 10772 7584 10836 7588
rect 10852 7644 10916 7648
rect 10852 7588 10856 7644
rect 10856 7588 10912 7644
rect 10912 7588 10916 7644
rect 10852 7584 10916 7588
rect 18612 7644 18676 7648
rect 18612 7588 18616 7644
rect 18616 7588 18672 7644
rect 18672 7588 18676 7644
rect 18612 7584 18676 7588
rect 18692 7644 18756 7648
rect 18692 7588 18696 7644
rect 18696 7588 18752 7644
rect 18752 7588 18756 7644
rect 18692 7584 18756 7588
rect 18772 7644 18836 7648
rect 18772 7588 18776 7644
rect 18776 7588 18832 7644
rect 18832 7588 18836 7644
rect 18772 7584 18836 7588
rect 18852 7644 18916 7648
rect 18852 7588 18856 7644
rect 18856 7588 18912 7644
rect 18912 7588 18916 7644
rect 18852 7584 18916 7588
rect 26612 7644 26676 7648
rect 26612 7588 26616 7644
rect 26616 7588 26672 7644
rect 26672 7588 26676 7644
rect 26612 7584 26676 7588
rect 26692 7644 26756 7648
rect 26692 7588 26696 7644
rect 26696 7588 26752 7644
rect 26752 7588 26756 7644
rect 26692 7584 26756 7588
rect 26772 7644 26836 7648
rect 26772 7588 26776 7644
rect 26776 7588 26832 7644
rect 26832 7588 26836 7644
rect 26772 7584 26836 7588
rect 26852 7644 26916 7648
rect 26852 7588 26856 7644
rect 26856 7588 26912 7644
rect 26912 7588 26916 7644
rect 26852 7584 26916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 9952 7100 10016 7104
rect 9952 7044 9956 7100
rect 9956 7044 10012 7100
rect 10012 7044 10016 7100
rect 9952 7040 10016 7044
rect 10032 7100 10096 7104
rect 10032 7044 10036 7100
rect 10036 7044 10092 7100
rect 10092 7044 10096 7100
rect 10032 7040 10096 7044
rect 10112 7100 10176 7104
rect 10112 7044 10116 7100
rect 10116 7044 10172 7100
rect 10172 7044 10176 7100
rect 10112 7040 10176 7044
rect 10192 7100 10256 7104
rect 10192 7044 10196 7100
rect 10196 7044 10252 7100
rect 10252 7044 10256 7100
rect 10192 7040 10256 7044
rect 17952 7100 18016 7104
rect 17952 7044 17956 7100
rect 17956 7044 18012 7100
rect 18012 7044 18016 7100
rect 17952 7040 18016 7044
rect 18032 7100 18096 7104
rect 18032 7044 18036 7100
rect 18036 7044 18092 7100
rect 18092 7044 18096 7100
rect 18032 7040 18096 7044
rect 18112 7100 18176 7104
rect 18112 7044 18116 7100
rect 18116 7044 18172 7100
rect 18172 7044 18176 7100
rect 18112 7040 18176 7044
rect 18192 7100 18256 7104
rect 18192 7044 18196 7100
rect 18196 7044 18252 7100
rect 18252 7044 18256 7100
rect 18192 7040 18256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 10612 6556 10676 6560
rect 10612 6500 10616 6556
rect 10616 6500 10672 6556
rect 10672 6500 10676 6556
rect 10612 6496 10676 6500
rect 10692 6556 10756 6560
rect 10692 6500 10696 6556
rect 10696 6500 10752 6556
rect 10752 6500 10756 6556
rect 10692 6496 10756 6500
rect 10772 6556 10836 6560
rect 10772 6500 10776 6556
rect 10776 6500 10832 6556
rect 10832 6500 10836 6556
rect 10772 6496 10836 6500
rect 10852 6556 10916 6560
rect 10852 6500 10856 6556
rect 10856 6500 10912 6556
rect 10912 6500 10916 6556
rect 10852 6496 10916 6500
rect 18612 6556 18676 6560
rect 18612 6500 18616 6556
rect 18616 6500 18672 6556
rect 18672 6500 18676 6556
rect 18612 6496 18676 6500
rect 18692 6556 18756 6560
rect 18692 6500 18696 6556
rect 18696 6500 18752 6556
rect 18752 6500 18756 6556
rect 18692 6496 18756 6500
rect 18772 6556 18836 6560
rect 18772 6500 18776 6556
rect 18776 6500 18832 6556
rect 18832 6500 18836 6556
rect 18772 6496 18836 6500
rect 18852 6556 18916 6560
rect 18852 6500 18856 6556
rect 18856 6500 18912 6556
rect 18912 6500 18916 6556
rect 18852 6496 18916 6500
rect 26612 6556 26676 6560
rect 26612 6500 26616 6556
rect 26616 6500 26672 6556
rect 26672 6500 26676 6556
rect 26612 6496 26676 6500
rect 26692 6556 26756 6560
rect 26692 6500 26696 6556
rect 26696 6500 26752 6556
rect 26752 6500 26756 6556
rect 26692 6496 26756 6500
rect 26772 6556 26836 6560
rect 26772 6500 26776 6556
rect 26776 6500 26832 6556
rect 26832 6500 26836 6556
rect 26772 6496 26836 6500
rect 26852 6556 26916 6560
rect 26852 6500 26856 6556
rect 26856 6500 26912 6556
rect 26912 6500 26916 6556
rect 26852 6496 26916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 9952 6012 10016 6016
rect 9952 5956 9956 6012
rect 9956 5956 10012 6012
rect 10012 5956 10016 6012
rect 9952 5952 10016 5956
rect 10032 6012 10096 6016
rect 10032 5956 10036 6012
rect 10036 5956 10092 6012
rect 10092 5956 10096 6012
rect 10032 5952 10096 5956
rect 10112 6012 10176 6016
rect 10112 5956 10116 6012
rect 10116 5956 10172 6012
rect 10172 5956 10176 6012
rect 10112 5952 10176 5956
rect 10192 6012 10256 6016
rect 10192 5956 10196 6012
rect 10196 5956 10252 6012
rect 10252 5956 10256 6012
rect 10192 5952 10256 5956
rect 17952 6012 18016 6016
rect 17952 5956 17956 6012
rect 17956 5956 18012 6012
rect 18012 5956 18016 6012
rect 17952 5952 18016 5956
rect 18032 6012 18096 6016
rect 18032 5956 18036 6012
rect 18036 5956 18092 6012
rect 18092 5956 18096 6012
rect 18032 5952 18096 5956
rect 18112 6012 18176 6016
rect 18112 5956 18116 6012
rect 18116 5956 18172 6012
rect 18172 5956 18176 6012
rect 18112 5952 18176 5956
rect 18192 6012 18256 6016
rect 18192 5956 18196 6012
rect 18196 5956 18252 6012
rect 18252 5956 18256 6012
rect 18192 5952 18256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 10612 5468 10676 5472
rect 10612 5412 10616 5468
rect 10616 5412 10672 5468
rect 10672 5412 10676 5468
rect 10612 5408 10676 5412
rect 10692 5468 10756 5472
rect 10692 5412 10696 5468
rect 10696 5412 10752 5468
rect 10752 5412 10756 5468
rect 10692 5408 10756 5412
rect 10772 5468 10836 5472
rect 10772 5412 10776 5468
rect 10776 5412 10832 5468
rect 10832 5412 10836 5468
rect 10772 5408 10836 5412
rect 10852 5468 10916 5472
rect 10852 5412 10856 5468
rect 10856 5412 10912 5468
rect 10912 5412 10916 5468
rect 10852 5408 10916 5412
rect 18612 5468 18676 5472
rect 18612 5412 18616 5468
rect 18616 5412 18672 5468
rect 18672 5412 18676 5468
rect 18612 5408 18676 5412
rect 18692 5468 18756 5472
rect 18692 5412 18696 5468
rect 18696 5412 18752 5468
rect 18752 5412 18756 5468
rect 18692 5408 18756 5412
rect 18772 5468 18836 5472
rect 18772 5412 18776 5468
rect 18776 5412 18832 5468
rect 18832 5412 18836 5468
rect 18772 5408 18836 5412
rect 18852 5468 18916 5472
rect 18852 5412 18856 5468
rect 18856 5412 18912 5468
rect 18912 5412 18916 5468
rect 18852 5408 18916 5412
rect 26612 5468 26676 5472
rect 26612 5412 26616 5468
rect 26616 5412 26672 5468
rect 26672 5412 26676 5468
rect 26612 5408 26676 5412
rect 26692 5468 26756 5472
rect 26692 5412 26696 5468
rect 26696 5412 26752 5468
rect 26752 5412 26756 5468
rect 26692 5408 26756 5412
rect 26772 5468 26836 5472
rect 26772 5412 26776 5468
rect 26776 5412 26832 5468
rect 26832 5412 26836 5468
rect 26772 5408 26836 5412
rect 26852 5468 26916 5472
rect 26852 5412 26856 5468
rect 26856 5412 26912 5468
rect 26912 5412 26916 5468
rect 26852 5408 26916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 9952 4924 10016 4928
rect 9952 4868 9956 4924
rect 9956 4868 10012 4924
rect 10012 4868 10016 4924
rect 9952 4864 10016 4868
rect 10032 4924 10096 4928
rect 10032 4868 10036 4924
rect 10036 4868 10092 4924
rect 10092 4868 10096 4924
rect 10032 4864 10096 4868
rect 10112 4924 10176 4928
rect 10112 4868 10116 4924
rect 10116 4868 10172 4924
rect 10172 4868 10176 4924
rect 10112 4864 10176 4868
rect 10192 4924 10256 4928
rect 10192 4868 10196 4924
rect 10196 4868 10252 4924
rect 10252 4868 10256 4924
rect 10192 4864 10256 4868
rect 17952 4924 18016 4928
rect 17952 4868 17956 4924
rect 17956 4868 18012 4924
rect 18012 4868 18016 4924
rect 17952 4864 18016 4868
rect 18032 4924 18096 4928
rect 18032 4868 18036 4924
rect 18036 4868 18092 4924
rect 18092 4868 18096 4924
rect 18032 4864 18096 4868
rect 18112 4924 18176 4928
rect 18112 4868 18116 4924
rect 18116 4868 18172 4924
rect 18172 4868 18176 4924
rect 18112 4864 18176 4868
rect 18192 4924 18256 4928
rect 18192 4868 18196 4924
rect 18196 4868 18252 4924
rect 18252 4868 18256 4924
rect 18192 4864 18256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 10612 4380 10676 4384
rect 10612 4324 10616 4380
rect 10616 4324 10672 4380
rect 10672 4324 10676 4380
rect 10612 4320 10676 4324
rect 10692 4380 10756 4384
rect 10692 4324 10696 4380
rect 10696 4324 10752 4380
rect 10752 4324 10756 4380
rect 10692 4320 10756 4324
rect 10772 4380 10836 4384
rect 10772 4324 10776 4380
rect 10776 4324 10832 4380
rect 10832 4324 10836 4380
rect 10772 4320 10836 4324
rect 10852 4380 10916 4384
rect 10852 4324 10856 4380
rect 10856 4324 10912 4380
rect 10912 4324 10916 4380
rect 10852 4320 10916 4324
rect 18612 4380 18676 4384
rect 18612 4324 18616 4380
rect 18616 4324 18672 4380
rect 18672 4324 18676 4380
rect 18612 4320 18676 4324
rect 18692 4380 18756 4384
rect 18692 4324 18696 4380
rect 18696 4324 18752 4380
rect 18752 4324 18756 4380
rect 18692 4320 18756 4324
rect 18772 4380 18836 4384
rect 18772 4324 18776 4380
rect 18776 4324 18832 4380
rect 18832 4324 18836 4380
rect 18772 4320 18836 4324
rect 18852 4380 18916 4384
rect 18852 4324 18856 4380
rect 18856 4324 18912 4380
rect 18912 4324 18916 4380
rect 18852 4320 18916 4324
rect 26612 4380 26676 4384
rect 26612 4324 26616 4380
rect 26616 4324 26672 4380
rect 26672 4324 26676 4380
rect 26612 4320 26676 4324
rect 26692 4380 26756 4384
rect 26692 4324 26696 4380
rect 26696 4324 26752 4380
rect 26752 4324 26756 4380
rect 26692 4320 26756 4324
rect 26772 4380 26836 4384
rect 26772 4324 26776 4380
rect 26776 4324 26832 4380
rect 26832 4324 26836 4380
rect 26772 4320 26836 4324
rect 26852 4380 26916 4384
rect 26852 4324 26856 4380
rect 26856 4324 26912 4380
rect 26912 4324 26916 4380
rect 26852 4320 26916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 9952 3836 10016 3840
rect 9952 3780 9956 3836
rect 9956 3780 10012 3836
rect 10012 3780 10016 3836
rect 9952 3776 10016 3780
rect 10032 3836 10096 3840
rect 10032 3780 10036 3836
rect 10036 3780 10092 3836
rect 10092 3780 10096 3836
rect 10032 3776 10096 3780
rect 10112 3836 10176 3840
rect 10112 3780 10116 3836
rect 10116 3780 10172 3836
rect 10172 3780 10176 3836
rect 10112 3776 10176 3780
rect 10192 3836 10256 3840
rect 10192 3780 10196 3836
rect 10196 3780 10252 3836
rect 10252 3780 10256 3836
rect 10192 3776 10256 3780
rect 17952 3836 18016 3840
rect 17952 3780 17956 3836
rect 17956 3780 18012 3836
rect 18012 3780 18016 3836
rect 17952 3776 18016 3780
rect 18032 3836 18096 3840
rect 18032 3780 18036 3836
rect 18036 3780 18092 3836
rect 18092 3780 18096 3836
rect 18032 3776 18096 3780
rect 18112 3836 18176 3840
rect 18112 3780 18116 3836
rect 18116 3780 18172 3836
rect 18172 3780 18176 3836
rect 18112 3776 18176 3780
rect 18192 3836 18256 3840
rect 18192 3780 18196 3836
rect 18196 3780 18252 3836
rect 18252 3780 18256 3836
rect 18192 3776 18256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 10612 3292 10676 3296
rect 10612 3236 10616 3292
rect 10616 3236 10672 3292
rect 10672 3236 10676 3292
rect 10612 3232 10676 3236
rect 10692 3292 10756 3296
rect 10692 3236 10696 3292
rect 10696 3236 10752 3292
rect 10752 3236 10756 3292
rect 10692 3232 10756 3236
rect 10772 3292 10836 3296
rect 10772 3236 10776 3292
rect 10776 3236 10832 3292
rect 10832 3236 10836 3292
rect 10772 3232 10836 3236
rect 10852 3292 10916 3296
rect 10852 3236 10856 3292
rect 10856 3236 10912 3292
rect 10912 3236 10916 3292
rect 10852 3232 10916 3236
rect 18612 3292 18676 3296
rect 18612 3236 18616 3292
rect 18616 3236 18672 3292
rect 18672 3236 18676 3292
rect 18612 3232 18676 3236
rect 18692 3292 18756 3296
rect 18692 3236 18696 3292
rect 18696 3236 18752 3292
rect 18752 3236 18756 3292
rect 18692 3232 18756 3236
rect 18772 3292 18836 3296
rect 18772 3236 18776 3292
rect 18776 3236 18832 3292
rect 18832 3236 18836 3292
rect 18772 3232 18836 3236
rect 18852 3292 18916 3296
rect 18852 3236 18856 3292
rect 18856 3236 18912 3292
rect 18912 3236 18916 3292
rect 18852 3232 18916 3236
rect 26612 3292 26676 3296
rect 26612 3236 26616 3292
rect 26616 3236 26672 3292
rect 26672 3236 26676 3292
rect 26612 3232 26676 3236
rect 26692 3292 26756 3296
rect 26692 3236 26696 3292
rect 26696 3236 26752 3292
rect 26752 3236 26756 3292
rect 26692 3232 26756 3236
rect 26772 3292 26836 3296
rect 26772 3236 26776 3292
rect 26776 3236 26832 3292
rect 26832 3236 26836 3292
rect 26772 3232 26836 3236
rect 26852 3292 26916 3296
rect 26852 3236 26856 3292
rect 26856 3236 26912 3292
rect 26912 3236 26916 3292
rect 26852 3232 26916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 9952 2748 10016 2752
rect 9952 2692 9956 2748
rect 9956 2692 10012 2748
rect 10012 2692 10016 2748
rect 9952 2688 10016 2692
rect 10032 2748 10096 2752
rect 10032 2692 10036 2748
rect 10036 2692 10092 2748
rect 10092 2692 10096 2748
rect 10032 2688 10096 2692
rect 10112 2748 10176 2752
rect 10112 2692 10116 2748
rect 10116 2692 10172 2748
rect 10172 2692 10176 2748
rect 10112 2688 10176 2692
rect 10192 2748 10256 2752
rect 10192 2692 10196 2748
rect 10196 2692 10252 2748
rect 10252 2692 10256 2748
rect 10192 2688 10256 2692
rect 17952 2748 18016 2752
rect 17952 2692 17956 2748
rect 17956 2692 18012 2748
rect 18012 2692 18016 2748
rect 17952 2688 18016 2692
rect 18032 2748 18096 2752
rect 18032 2692 18036 2748
rect 18036 2692 18092 2748
rect 18092 2692 18096 2748
rect 18032 2688 18096 2692
rect 18112 2748 18176 2752
rect 18112 2692 18116 2748
rect 18116 2692 18172 2748
rect 18172 2692 18176 2748
rect 18112 2688 18176 2692
rect 18192 2748 18256 2752
rect 18192 2692 18196 2748
rect 18196 2692 18252 2748
rect 18252 2692 18256 2748
rect 18192 2688 18256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
rect 10612 2204 10676 2208
rect 10612 2148 10616 2204
rect 10616 2148 10672 2204
rect 10672 2148 10676 2204
rect 10612 2144 10676 2148
rect 10692 2204 10756 2208
rect 10692 2148 10696 2204
rect 10696 2148 10752 2204
rect 10752 2148 10756 2204
rect 10692 2144 10756 2148
rect 10772 2204 10836 2208
rect 10772 2148 10776 2204
rect 10776 2148 10832 2204
rect 10832 2148 10836 2204
rect 10772 2144 10836 2148
rect 10852 2204 10916 2208
rect 10852 2148 10856 2204
rect 10856 2148 10912 2204
rect 10912 2148 10916 2204
rect 10852 2144 10916 2148
rect 18612 2204 18676 2208
rect 18612 2148 18616 2204
rect 18616 2148 18672 2204
rect 18672 2148 18676 2204
rect 18612 2144 18676 2148
rect 18692 2204 18756 2208
rect 18692 2148 18696 2204
rect 18696 2148 18752 2204
rect 18752 2148 18756 2204
rect 18692 2144 18756 2148
rect 18772 2204 18836 2208
rect 18772 2148 18776 2204
rect 18776 2148 18832 2204
rect 18832 2148 18836 2204
rect 18772 2144 18836 2148
rect 18852 2204 18916 2208
rect 18852 2148 18856 2204
rect 18856 2148 18912 2204
rect 18912 2148 18916 2204
rect 18852 2144 18916 2148
rect 26612 2204 26676 2208
rect 26612 2148 26616 2204
rect 26616 2148 26672 2204
rect 26672 2148 26676 2204
rect 26612 2144 26676 2148
rect 26692 2204 26756 2208
rect 26692 2148 26696 2204
rect 26696 2148 26752 2204
rect 26752 2148 26756 2204
rect 26692 2144 26756 2148
rect 26772 2204 26836 2208
rect 26772 2148 26776 2204
rect 26776 2148 26832 2204
rect 26832 2148 26836 2204
rect 26772 2144 26836 2148
rect 26852 2204 26916 2208
rect 26852 2148 26856 2204
rect 26856 2148 26912 2204
rect 26912 2148 26916 2204
rect 26852 2144 26916 2148
<< metal4 >>
rect 1944 27776 2264 27792
rect 1944 27712 1952 27776
rect 2016 27712 2032 27776
rect 2096 27712 2112 27776
rect 2176 27712 2192 27776
rect 2256 27712 2264 27776
rect 1944 26688 2264 27712
rect 1944 26624 1952 26688
rect 2016 26624 2032 26688
rect 2096 26624 2112 26688
rect 2176 26624 2192 26688
rect 2256 26624 2264 26688
rect 1944 25600 2264 26624
rect 1944 25536 1952 25600
rect 2016 25536 2032 25600
rect 2096 25536 2112 25600
rect 2176 25536 2192 25600
rect 2256 25536 2264 25600
rect 1944 24512 2264 25536
rect 1944 24448 1952 24512
rect 2016 24448 2032 24512
rect 2096 24448 2112 24512
rect 2176 24448 2192 24512
rect 2256 24448 2264 24512
rect 1944 23424 2264 24448
rect 1944 23360 1952 23424
rect 2016 23360 2032 23424
rect 2096 23360 2112 23424
rect 2176 23360 2192 23424
rect 2256 23360 2264 23424
rect 1944 22336 2264 23360
rect 1944 22272 1952 22336
rect 2016 22272 2032 22336
rect 2096 22272 2112 22336
rect 2176 22272 2192 22336
rect 2256 22272 2264 22336
rect 1944 21248 2264 22272
rect 1944 21184 1952 21248
rect 2016 21184 2032 21248
rect 2096 21184 2112 21248
rect 2176 21184 2192 21248
rect 2256 21184 2264 21248
rect 1944 20160 2264 21184
rect 1944 20096 1952 20160
rect 2016 20096 2032 20160
rect 2096 20096 2112 20160
rect 2176 20096 2192 20160
rect 2256 20096 2264 20160
rect 1944 19072 2264 20096
rect 1944 19008 1952 19072
rect 2016 19008 2032 19072
rect 2096 19008 2112 19072
rect 2176 19008 2192 19072
rect 2256 19008 2264 19072
rect 1944 17984 2264 19008
rect 1944 17920 1952 17984
rect 2016 17920 2032 17984
rect 2096 17920 2112 17984
rect 2176 17920 2192 17984
rect 2256 17920 2264 17984
rect 1944 16896 2264 17920
rect 1944 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2264 16896
rect 1944 15808 2264 16832
rect 1944 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2264 15808
rect 1944 14720 2264 15744
rect 1944 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2264 14720
rect 1944 13632 2264 14656
rect 1944 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2264 13632
rect 1944 12544 2264 13568
rect 1944 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2264 12544
rect 1944 11456 2264 12480
rect 1944 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2264 11456
rect 1944 10368 2264 11392
rect 1944 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2264 10368
rect 1944 9280 2264 10304
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8192 2264 9216
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 27232 2924 27792
rect 2604 27168 2612 27232
rect 2676 27168 2692 27232
rect 2756 27168 2772 27232
rect 2836 27168 2852 27232
rect 2916 27168 2924 27232
rect 2604 26144 2924 27168
rect 2604 26080 2612 26144
rect 2676 26080 2692 26144
rect 2756 26080 2772 26144
rect 2836 26080 2852 26144
rect 2916 26080 2924 26144
rect 2604 25056 2924 26080
rect 2604 24992 2612 25056
rect 2676 24992 2692 25056
rect 2756 24992 2772 25056
rect 2836 24992 2852 25056
rect 2916 24992 2924 25056
rect 2604 23968 2924 24992
rect 2604 23904 2612 23968
rect 2676 23904 2692 23968
rect 2756 23904 2772 23968
rect 2836 23904 2852 23968
rect 2916 23904 2924 23968
rect 2604 22880 2924 23904
rect 2604 22816 2612 22880
rect 2676 22816 2692 22880
rect 2756 22816 2772 22880
rect 2836 22816 2852 22880
rect 2916 22816 2924 22880
rect 2604 21792 2924 22816
rect 2604 21728 2612 21792
rect 2676 21728 2692 21792
rect 2756 21728 2772 21792
rect 2836 21728 2852 21792
rect 2916 21728 2924 21792
rect 2604 20704 2924 21728
rect 2604 20640 2612 20704
rect 2676 20640 2692 20704
rect 2756 20640 2772 20704
rect 2836 20640 2852 20704
rect 2916 20640 2924 20704
rect 2604 19616 2924 20640
rect 2604 19552 2612 19616
rect 2676 19552 2692 19616
rect 2756 19552 2772 19616
rect 2836 19552 2852 19616
rect 2916 19552 2924 19616
rect 2604 18528 2924 19552
rect 2604 18464 2612 18528
rect 2676 18464 2692 18528
rect 2756 18464 2772 18528
rect 2836 18464 2852 18528
rect 2916 18464 2924 18528
rect 2604 17440 2924 18464
rect 2604 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2924 17440
rect 2604 16352 2924 17376
rect 2604 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2924 16352
rect 2604 15264 2924 16288
rect 2604 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2924 15264
rect 2604 14176 2924 15200
rect 2604 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2924 14176
rect 2604 13088 2924 14112
rect 2604 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2924 13088
rect 2604 12000 2924 13024
rect 2604 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2924 12000
rect 2604 10912 2924 11936
rect 2604 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2924 10912
rect 2604 9824 2924 10848
rect 2604 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2924 9824
rect 2604 8736 2924 9760
rect 2604 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3296 2924 4320
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
rect 9944 27776 10264 27792
rect 9944 27712 9952 27776
rect 10016 27712 10032 27776
rect 10096 27712 10112 27776
rect 10176 27712 10192 27776
rect 10256 27712 10264 27776
rect 9944 26688 10264 27712
rect 9944 26624 9952 26688
rect 10016 26624 10032 26688
rect 10096 26624 10112 26688
rect 10176 26624 10192 26688
rect 10256 26624 10264 26688
rect 9944 25600 10264 26624
rect 9944 25536 9952 25600
rect 10016 25536 10032 25600
rect 10096 25536 10112 25600
rect 10176 25536 10192 25600
rect 10256 25536 10264 25600
rect 9944 24512 10264 25536
rect 9944 24448 9952 24512
rect 10016 24448 10032 24512
rect 10096 24448 10112 24512
rect 10176 24448 10192 24512
rect 10256 24448 10264 24512
rect 9944 23424 10264 24448
rect 9944 23360 9952 23424
rect 10016 23360 10032 23424
rect 10096 23360 10112 23424
rect 10176 23360 10192 23424
rect 10256 23360 10264 23424
rect 9944 22336 10264 23360
rect 9944 22272 9952 22336
rect 10016 22272 10032 22336
rect 10096 22272 10112 22336
rect 10176 22272 10192 22336
rect 10256 22272 10264 22336
rect 9944 21248 10264 22272
rect 9944 21184 9952 21248
rect 10016 21184 10032 21248
rect 10096 21184 10112 21248
rect 10176 21184 10192 21248
rect 10256 21184 10264 21248
rect 9944 20160 10264 21184
rect 9944 20096 9952 20160
rect 10016 20096 10032 20160
rect 10096 20096 10112 20160
rect 10176 20096 10192 20160
rect 10256 20096 10264 20160
rect 9944 19072 10264 20096
rect 9944 19008 9952 19072
rect 10016 19008 10032 19072
rect 10096 19008 10112 19072
rect 10176 19008 10192 19072
rect 10256 19008 10264 19072
rect 9944 17984 10264 19008
rect 9944 17920 9952 17984
rect 10016 17920 10032 17984
rect 10096 17920 10112 17984
rect 10176 17920 10192 17984
rect 10256 17920 10264 17984
rect 9944 16896 10264 17920
rect 9944 16832 9952 16896
rect 10016 16832 10032 16896
rect 10096 16832 10112 16896
rect 10176 16832 10192 16896
rect 10256 16832 10264 16896
rect 9944 15808 10264 16832
rect 9944 15744 9952 15808
rect 10016 15744 10032 15808
rect 10096 15744 10112 15808
rect 10176 15744 10192 15808
rect 10256 15744 10264 15808
rect 9944 14720 10264 15744
rect 9944 14656 9952 14720
rect 10016 14656 10032 14720
rect 10096 14656 10112 14720
rect 10176 14656 10192 14720
rect 10256 14656 10264 14720
rect 9944 13632 10264 14656
rect 9944 13568 9952 13632
rect 10016 13568 10032 13632
rect 10096 13568 10112 13632
rect 10176 13568 10192 13632
rect 10256 13568 10264 13632
rect 9944 12544 10264 13568
rect 9944 12480 9952 12544
rect 10016 12480 10032 12544
rect 10096 12480 10112 12544
rect 10176 12480 10192 12544
rect 10256 12480 10264 12544
rect 9944 11456 10264 12480
rect 9944 11392 9952 11456
rect 10016 11392 10032 11456
rect 10096 11392 10112 11456
rect 10176 11392 10192 11456
rect 10256 11392 10264 11456
rect 9944 10368 10264 11392
rect 9944 10304 9952 10368
rect 10016 10304 10032 10368
rect 10096 10304 10112 10368
rect 10176 10304 10192 10368
rect 10256 10304 10264 10368
rect 9944 9280 10264 10304
rect 9944 9216 9952 9280
rect 10016 9216 10032 9280
rect 10096 9216 10112 9280
rect 10176 9216 10192 9280
rect 10256 9216 10264 9280
rect 9944 8192 10264 9216
rect 9944 8128 9952 8192
rect 10016 8128 10032 8192
rect 10096 8128 10112 8192
rect 10176 8128 10192 8192
rect 10256 8128 10264 8192
rect 9944 7104 10264 8128
rect 9944 7040 9952 7104
rect 10016 7040 10032 7104
rect 10096 7040 10112 7104
rect 10176 7040 10192 7104
rect 10256 7040 10264 7104
rect 9944 6016 10264 7040
rect 9944 5952 9952 6016
rect 10016 5952 10032 6016
rect 10096 5952 10112 6016
rect 10176 5952 10192 6016
rect 10256 5952 10264 6016
rect 9944 4928 10264 5952
rect 9944 4864 9952 4928
rect 10016 4864 10032 4928
rect 10096 4864 10112 4928
rect 10176 4864 10192 4928
rect 10256 4864 10264 4928
rect 9944 3840 10264 4864
rect 9944 3776 9952 3840
rect 10016 3776 10032 3840
rect 10096 3776 10112 3840
rect 10176 3776 10192 3840
rect 10256 3776 10264 3840
rect 9944 2752 10264 3776
rect 9944 2688 9952 2752
rect 10016 2688 10032 2752
rect 10096 2688 10112 2752
rect 10176 2688 10192 2752
rect 10256 2688 10264 2752
rect 9944 2128 10264 2688
rect 10604 27232 10924 27792
rect 10604 27168 10612 27232
rect 10676 27168 10692 27232
rect 10756 27168 10772 27232
rect 10836 27168 10852 27232
rect 10916 27168 10924 27232
rect 10604 26144 10924 27168
rect 10604 26080 10612 26144
rect 10676 26080 10692 26144
rect 10756 26080 10772 26144
rect 10836 26080 10852 26144
rect 10916 26080 10924 26144
rect 10604 25056 10924 26080
rect 10604 24992 10612 25056
rect 10676 24992 10692 25056
rect 10756 24992 10772 25056
rect 10836 24992 10852 25056
rect 10916 24992 10924 25056
rect 10604 23968 10924 24992
rect 10604 23904 10612 23968
rect 10676 23904 10692 23968
rect 10756 23904 10772 23968
rect 10836 23904 10852 23968
rect 10916 23904 10924 23968
rect 10604 22880 10924 23904
rect 10604 22816 10612 22880
rect 10676 22816 10692 22880
rect 10756 22816 10772 22880
rect 10836 22816 10852 22880
rect 10916 22816 10924 22880
rect 10604 21792 10924 22816
rect 10604 21728 10612 21792
rect 10676 21728 10692 21792
rect 10756 21728 10772 21792
rect 10836 21728 10852 21792
rect 10916 21728 10924 21792
rect 10604 20704 10924 21728
rect 10604 20640 10612 20704
rect 10676 20640 10692 20704
rect 10756 20640 10772 20704
rect 10836 20640 10852 20704
rect 10916 20640 10924 20704
rect 10604 19616 10924 20640
rect 10604 19552 10612 19616
rect 10676 19552 10692 19616
rect 10756 19552 10772 19616
rect 10836 19552 10852 19616
rect 10916 19552 10924 19616
rect 10604 18528 10924 19552
rect 10604 18464 10612 18528
rect 10676 18464 10692 18528
rect 10756 18464 10772 18528
rect 10836 18464 10852 18528
rect 10916 18464 10924 18528
rect 10604 17440 10924 18464
rect 10604 17376 10612 17440
rect 10676 17376 10692 17440
rect 10756 17376 10772 17440
rect 10836 17376 10852 17440
rect 10916 17376 10924 17440
rect 10604 16352 10924 17376
rect 10604 16288 10612 16352
rect 10676 16288 10692 16352
rect 10756 16288 10772 16352
rect 10836 16288 10852 16352
rect 10916 16288 10924 16352
rect 10604 15264 10924 16288
rect 10604 15200 10612 15264
rect 10676 15200 10692 15264
rect 10756 15200 10772 15264
rect 10836 15200 10852 15264
rect 10916 15200 10924 15264
rect 10604 14176 10924 15200
rect 10604 14112 10612 14176
rect 10676 14112 10692 14176
rect 10756 14112 10772 14176
rect 10836 14112 10852 14176
rect 10916 14112 10924 14176
rect 10604 13088 10924 14112
rect 10604 13024 10612 13088
rect 10676 13024 10692 13088
rect 10756 13024 10772 13088
rect 10836 13024 10852 13088
rect 10916 13024 10924 13088
rect 10604 12000 10924 13024
rect 10604 11936 10612 12000
rect 10676 11936 10692 12000
rect 10756 11936 10772 12000
rect 10836 11936 10852 12000
rect 10916 11936 10924 12000
rect 10604 10912 10924 11936
rect 10604 10848 10612 10912
rect 10676 10848 10692 10912
rect 10756 10848 10772 10912
rect 10836 10848 10852 10912
rect 10916 10848 10924 10912
rect 10604 9824 10924 10848
rect 10604 9760 10612 9824
rect 10676 9760 10692 9824
rect 10756 9760 10772 9824
rect 10836 9760 10852 9824
rect 10916 9760 10924 9824
rect 10604 8736 10924 9760
rect 10604 8672 10612 8736
rect 10676 8672 10692 8736
rect 10756 8672 10772 8736
rect 10836 8672 10852 8736
rect 10916 8672 10924 8736
rect 10604 7648 10924 8672
rect 10604 7584 10612 7648
rect 10676 7584 10692 7648
rect 10756 7584 10772 7648
rect 10836 7584 10852 7648
rect 10916 7584 10924 7648
rect 10604 6560 10924 7584
rect 10604 6496 10612 6560
rect 10676 6496 10692 6560
rect 10756 6496 10772 6560
rect 10836 6496 10852 6560
rect 10916 6496 10924 6560
rect 10604 5472 10924 6496
rect 10604 5408 10612 5472
rect 10676 5408 10692 5472
rect 10756 5408 10772 5472
rect 10836 5408 10852 5472
rect 10916 5408 10924 5472
rect 10604 4384 10924 5408
rect 10604 4320 10612 4384
rect 10676 4320 10692 4384
rect 10756 4320 10772 4384
rect 10836 4320 10852 4384
rect 10916 4320 10924 4384
rect 10604 3296 10924 4320
rect 10604 3232 10612 3296
rect 10676 3232 10692 3296
rect 10756 3232 10772 3296
rect 10836 3232 10852 3296
rect 10916 3232 10924 3296
rect 10604 2208 10924 3232
rect 10604 2144 10612 2208
rect 10676 2144 10692 2208
rect 10756 2144 10772 2208
rect 10836 2144 10852 2208
rect 10916 2144 10924 2208
rect 10604 2128 10924 2144
rect 17944 27776 18264 27792
rect 17944 27712 17952 27776
rect 18016 27712 18032 27776
rect 18096 27712 18112 27776
rect 18176 27712 18192 27776
rect 18256 27712 18264 27776
rect 17944 26688 18264 27712
rect 17944 26624 17952 26688
rect 18016 26624 18032 26688
rect 18096 26624 18112 26688
rect 18176 26624 18192 26688
rect 18256 26624 18264 26688
rect 17944 25600 18264 26624
rect 17944 25536 17952 25600
rect 18016 25536 18032 25600
rect 18096 25536 18112 25600
rect 18176 25536 18192 25600
rect 18256 25536 18264 25600
rect 17944 24512 18264 25536
rect 17944 24448 17952 24512
rect 18016 24448 18032 24512
rect 18096 24448 18112 24512
rect 18176 24448 18192 24512
rect 18256 24448 18264 24512
rect 17944 23424 18264 24448
rect 17944 23360 17952 23424
rect 18016 23360 18032 23424
rect 18096 23360 18112 23424
rect 18176 23360 18192 23424
rect 18256 23360 18264 23424
rect 17944 22336 18264 23360
rect 17944 22272 17952 22336
rect 18016 22272 18032 22336
rect 18096 22272 18112 22336
rect 18176 22272 18192 22336
rect 18256 22272 18264 22336
rect 17944 21248 18264 22272
rect 17944 21184 17952 21248
rect 18016 21184 18032 21248
rect 18096 21184 18112 21248
rect 18176 21184 18192 21248
rect 18256 21184 18264 21248
rect 17944 20160 18264 21184
rect 17944 20096 17952 20160
rect 18016 20096 18032 20160
rect 18096 20096 18112 20160
rect 18176 20096 18192 20160
rect 18256 20096 18264 20160
rect 17944 19072 18264 20096
rect 17944 19008 17952 19072
rect 18016 19008 18032 19072
rect 18096 19008 18112 19072
rect 18176 19008 18192 19072
rect 18256 19008 18264 19072
rect 17944 17984 18264 19008
rect 17944 17920 17952 17984
rect 18016 17920 18032 17984
rect 18096 17920 18112 17984
rect 18176 17920 18192 17984
rect 18256 17920 18264 17984
rect 17944 16896 18264 17920
rect 17944 16832 17952 16896
rect 18016 16832 18032 16896
rect 18096 16832 18112 16896
rect 18176 16832 18192 16896
rect 18256 16832 18264 16896
rect 17944 15808 18264 16832
rect 17944 15744 17952 15808
rect 18016 15744 18032 15808
rect 18096 15744 18112 15808
rect 18176 15744 18192 15808
rect 18256 15744 18264 15808
rect 17944 14720 18264 15744
rect 17944 14656 17952 14720
rect 18016 14656 18032 14720
rect 18096 14656 18112 14720
rect 18176 14656 18192 14720
rect 18256 14656 18264 14720
rect 17944 13632 18264 14656
rect 17944 13568 17952 13632
rect 18016 13568 18032 13632
rect 18096 13568 18112 13632
rect 18176 13568 18192 13632
rect 18256 13568 18264 13632
rect 17944 12544 18264 13568
rect 17944 12480 17952 12544
rect 18016 12480 18032 12544
rect 18096 12480 18112 12544
rect 18176 12480 18192 12544
rect 18256 12480 18264 12544
rect 17944 11456 18264 12480
rect 17944 11392 17952 11456
rect 18016 11392 18032 11456
rect 18096 11392 18112 11456
rect 18176 11392 18192 11456
rect 18256 11392 18264 11456
rect 17944 10368 18264 11392
rect 17944 10304 17952 10368
rect 18016 10304 18032 10368
rect 18096 10304 18112 10368
rect 18176 10304 18192 10368
rect 18256 10304 18264 10368
rect 17944 9280 18264 10304
rect 17944 9216 17952 9280
rect 18016 9216 18032 9280
rect 18096 9216 18112 9280
rect 18176 9216 18192 9280
rect 18256 9216 18264 9280
rect 17944 8192 18264 9216
rect 17944 8128 17952 8192
rect 18016 8128 18032 8192
rect 18096 8128 18112 8192
rect 18176 8128 18192 8192
rect 18256 8128 18264 8192
rect 17944 7104 18264 8128
rect 17944 7040 17952 7104
rect 18016 7040 18032 7104
rect 18096 7040 18112 7104
rect 18176 7040 18192 7104
rect 18256 7040 18264 7104
rect 17944 6016 18264 7040
rect 17944 5952 17952 6016
rect 18016 5952 18032 6016
rect 18096 5952 18112 6016
rect 18176 5952 18192 6016
rect 18256 5952 18264 6016
rect 17944 4928 18264 5952
rect 17944 4864 17952 4928
rect 18016 4864 18032 4928
rect 18096 4864 18112 4928
rect 18176 4864 18192 4928
rect 18256 4864 18264 4928
rect 17944 3840 18264 4864
rect 17944 3776 17952 3840
rect 18016 3776 18032 3840
rect 18096 3776 18112 3840
rect 18176 3776 18192 3840
rect 18256 3776 18264 3840
rect 17944 2752 18264 3776
rect 17944 2688 17952 2752
rect 18016 2688 18032 2752
rect 18096 2688 18112 2752
rect 18176 2688 18192 2752
rect 18256 2688 18264 2752
rect 17944 2128 18264 2688
rect 18604 27232 18924 27792
rect 18604 27168 18612 27232
rect 18676 27168 18692 27232
rect 18756 27168 18772 27232
rect 18836 27168 18852 27232
rect 18916 27168 18924 27232
rect 18604 26144 18924 27168
rect 18604 26080 18612 26144
rect 18676 26080 18692 26144
rect 18756 26080 18772 26144
rect 18836 26080 18852 26144
rect 18916 26080 18924 26144
rect 18604 25056 18924 26080
rect 18604 24992 18612 25056
rect 18676 24992 18692 25056
rect 18756 24992 18772 25056
rect 18836 24992 18852 25056
rect 18916 24992 18924 25056
rect 18604 23968 18924 24992
rect 18604 23904 18612 23968
rect 18676 23904 18692 23968
rect 18756 23904 18772 23968
rect 18836 23904 18852 23968
rect 18916 23904 18924 23968
rect 18604 22880 18924 23904
rect 18604 22816 18612 22880
rect 18676 22816 18692 22880
rect 18756 22816 18772 22880
rect 18836 22816 18852 22880
rect 18916 22816 18924 22880
rect 18604 21792 18924 22816
rect 18604 21728 18612 21792
rect 18676 21728 18692 21792
rect 18756 21728 18772 21792
rect 18836 21728 18852 21792
rect 18916 21728 18924 21792
rect 18604 20704 18924 21728
rect 18604 20640 18612 20704
rect 18676 20640 18692 20704
rect 18756 20640 18772 20704
rect 18836 20640 18852 20704
rect 18916 20640 18924 20704
rect 18604 19616 18924 20640
rect 18604 19552 18612 19616
rect 18676 19552 18692 19616
rect 18756 19552 18772 19616
rect 18836 19552 18852 19616
rect 18916 19552 18924 19616
rect 18604 18528 18924 19552
rect 18604 18464 18612 18528
rect 18676 18464 18692 18528
rect 18756 18464 18772 18528
rect 18836 18464 18852 18528
rect 18916 18464 18924 18528
rect 18604 17440 18924 18464
rect 18604 17376 18612 17440
rect 18676 17376 18692 17440
rect 18756 17376 18772 17440
rect 18836 17376 18852 17440
rect 18916 17376 18924 17440
rect 18604 16352 18924 17376
rect 18604 16288 18612 16352
rect 18676 16288 18692 16352
rect 18756 16288 18772 16352
rect 18836 16288 18852 16352
rect 18916 16288 18924 16352
rect 18604 15264 18924 16288
rect 18604 15200 18612 15264
rect 18676 15200 18692 15264
rect 18756 15200 18772 15264
rect 18836 15200 18852 15264
rect 18916 15200 18924 15264
rect 18604 14176 18924 15200
rect 18604 14112 18612 14176
rect 18676 14112 18692 14176
rect 18756 14112 18772 14176
rect 18836 14112 18852 14176
rect 18916 14112 18924 14176
rect 18604 13088 18924 14112
rect 18604 13024 18612 13088
rect 18676 13024 18692 13088
rect 18756 13024 18772 13088
rect 18836 13024 18852 13088
rect 18916 13024 18924 13088
rect 18604 12000 18924 13024
rect 18604 11936 18612 12000
rect 18676 11936 18692 12000
rect 18756 11936 18772 12000
rect 18836 11936 18852 12000
rect 18916 11936 18924 12000
rect 18604 10912 18924 11936
rect 18604 10848 18612 10912
rect 18676 10848 18692 10912
rect 18756 10848 18772 10912
rect 18836 10848 18852 10912
rect 18916 10848 18924 10912
rect 18604 9824 18924 10848
rect 18604 9760 18612 9824
rect 18676 9760 18692 9824
rect 18756 9760 18772 9824
rect 18836 9760 18852 9824
rect 18916 9760 18924 9824
rect 18604 8736 18924 9760
rect 18604 8672 18612 8736
rect 18676 8672 18692 8736
rect 18756 8672 18772 8736
rect 18836 8672 18852 8736
rect 18916 8672 18924 8736
rect 18604 7648 18924 8672
rect 18604 7584 18612 7648
rect 18676 7584 18692 7648
rect 18756 7584 18772 7648
rect 18836 7584 18852 7648
rect 18916 7584 18924 7648
rect 18604 6560 18924 7584
rect 18604 6496 18612 6560
rect 18676 6496 18692 6560
rect 18756 6496 18772 6560
rect 18836 6496 18852 6560
rect 18916 6496 18924 6560
rect 18604 5472 18924 6496
rect 18604 5408 18612 5472
rect 18676 5408 18692 5472
rect 18756 5408 18772 5472
rect 18836 5408 18852 5472
rect 18916 5408 18924 5472
rect 18604 4384 18924 5408
rect 18604 4320 18612 4384
rect 18676 4320 18692 4384
rect 18756 4320 18772 4384
rect 18836 4320 18852 4384
rect 18916 4320 18924 4384
rect 18604 3296 18924 4320
rect 18604 3232 18612 3296
rect 18676 3232 18692 3296
rect 18756 3232 18772 3296
rect 18836 3232 18852 3296
rect 18916 3232 18924 3296
rect 18604 2208 18924 3232
rect 18604 2144 18612 2208
rect 18676 2144 18692 2208
rect 18756 2144 18772 2208
rect 18836 2144 18852 2208
rect 18916 2144 18924 2208
rect 18604 2128 18924 2144
rect 25944 27776 26264 27792
rect 25944 27712 25952 27776
rect 26016 27712 26032 27776
rect 26096 27712 26112 27776
rect 26176 27712 26192 27776
rect 26256 27712 26264 27776
rect 25944 26688 26264 27712
rect 25944 26624 25952 26688
rect 26016 26624 26032 26688
rect 26096 26624 26112 26688
rect 26176 26624 26192 26688
rect 26256 26624 26264 26688
rect 25944 25600 26264 26624
rect 25944 25536 25952 25600
rect 26016 25536 26032 25600
rect 26096 25536 26112 25600
rect 26176 25536 26192 25600
rect 26256 25536 26264 25600
rect 25944 24512 26264 25536
rect 25944 24448 25952 24512
rect 26016 24448 26032 24512
rect 26096 24448 26112 24512
rect 26176 24448 26192 24512
rect 26256 24448 26264 24512
rect 25944 23424 26264 24448
rect 25944 23360 25952 23424
rect 26016 23360 26032 23424
rect 26096 23360 26112 23424
rect 26176 23360 26192 23424
rect 26256 23360 26264 23424
rect 25944 22336 26264 23360
rect 25944 22272 25952 22336
rect 26016 22272 26032 22336
rect 26096 22272 26112 22336
rect 26176 22272 26192 22336
rect 26256 22272 26264 22336
rect 25944 21248 26264 22272
rect 25944 21184 25952 21248
rect 26016 21184 26032 21248
rect 26096 21184 26112 21248
rect 26176 21184 26192 21248
rect 26256 21184 26264 21248
rect 25944 20160 26264 21184
rect 25944 20096 25952 20160
rect 26016 20096 26032 20160
rect 26096 20096 26112 20160
rect 26176 20096 26192 20160
rect 26256 20096 26264 20160
rect 25944 19072 26264 20096
rect 25944 19008 25952 19072
rect 26016 19008 26032 19072
rect 26096 19008 26112 19072
rect 26176 19008 26192 19072
rect 26256 19008 26264 19072
rect 25944 17984 26264 19008
rect 25944 17920 25952 17984
rect 26016 17920 26032 17984
rect 26096 17920 26112 17984
rect 26176 17920 26192 17984
rect 26256 17920 26264 17984
rect 25944 16896 26264 17920
rect 25944 16832 25952 16896
rect 26016 16832 26032 16896
rect 26096 16832 26112 16896
rect 26176 16832 26192 16896
rect 26256 16832 26264 16896
rect 25944 15808 26264 16832
rect 25944 15744 25952 15808
rect 26016 15744 26032 15808
rect 26096 15744 26112 15808
rect 26176 15744 26192 15808
rect 26256 15744 26264 15808
rect 25944 14720 26264 15744
rect 25944 14656 25952 14720
rect 26016 14656 26032 14720
rect 26096 14656 26112 14720
rect 26176 14656 26192 14720
rect 26256 14656 26264 14720
rect 25944 13632 26264 14656
rect 25944 13568 25952 13632
rect 26016 13568 26032 13632
rect 26096 13568 26112 13632
rect 26176 13568 26192 13632
rect 26256 13568 26264 13632
rect 25944 12544 26264 13568
rect 25944 12480 25952 12544
rect 26016 12480 26032 12544
rect 26096 12480 26112 12544
rect 26176 12480 26192 12544
rect 26256 12480 26264 12544
rect 25944 11456 26264 12480
rect 25944 11392 25952 11456
rect 26016 11392 26032 11456
rect 26096 11392 26112 11456
rect 26176 11392 26192 11456
rect 26256 11392 26264 11456
rect 25944 10368 26264 11392
rect 25944 10304 25952 10368
rect 26016 10304 26032 10368
rect 26096 10304 26112 10368
rect 26176 10304 26192 10368
rect 26256 10304 26264 10368
rect 25944 9280 26264 10304
rect 25944 9216 25952 9280
rect 26016 9216 26032 9280
rect 26096 9216 26112 9280
rect 26176 9216 26192 9280
rect 26256 9216 26264 9280
rect 25944 8192 26264 9216
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 2128 26264 2688
rect 26604 27232 26924 27792
rect 26604 27168 26612 27232
rect 26676 27168 26692 27232
rect 26756 27168 26772 27232
rect 26836 27168 26852 27232
rect 26916 27168 26924 27232
rect 26604 26144 26924 27168
rect 26604 26080 26612 26144
rect 26676 26080 26692 26144
rect 26756 26080 26772 26144
rect 26836 26080 26852 26144
rect 26916 26080 26924 26144
rect 26604 25056 26924 26080
rect 26604 24992 26612 25056
rect 26676 24992 26692 25056
rect 26756 24992 26772 25056
rect 26836 24992 26852 25056
rect 26916 24992 26924 25056
rect 26604 23968 26924 24992
rect 26604 23904 26612 23968
rect 26676 23904 26692 23968
rect 26756 23904 26772 23968
rect 26836 23904 26852 23968
rect 26916 23904 26924 23968
rect 26604 22880 26924 23904
rect 26604 22816 26612 22880
rect 26676 22816 26692 22880
rect 26756 22816 26772 22880
rect 26836 22816 26852 22880
rect 26916 22816 26924 22880
rect 26604 21792 26924 22816
rect 26604 21728 26612 21792
rect 26676 21728 26692 21792
rect 26756 21728 26772 21792
rect 26836 21728 26852 21792
rect 26916 21728 26924 21792
rect 26604 20704 26924 21728
rect 26604 20640 26612 20704
rect 26676 20640 26692 20704
rect 26756 20640 26772 20704
rect 26836 20640 26852 20704
rect 26916 20640 26924 20704
rect 26604 19616 26924 20640
rect 26604 19552 26612 19616
rect 26676 19552 26692 19616
rect 26756 19552 26772 19616
rect 26836 19552 26852 19616
rect 26916 19552 26924 19616
rect 26604 18528 26924 19552
rect 26604 18464 26612 18528
rect 26676 18464 26692 18528
rect 26756 18464 26772 18528
rect 26836 18464 26852 18528
rect 26916 18464 26924 18528
rect 26604 17440 26924 18464
rect 26604 17376 26612 17440
rect 26676 17376 26692 17440
rect 26756 17376 26772 17440
rect 26836 17376 26852 17440
rect 26916 17376 26924 17440
rect 26604 16352 26924 17376
rect 26604 16288 26612 16352
rect 26676 16288 26692 16352
rect 26756 16288 26772 16352
rect 26836 16288 26852 16352
rect 26916 16288 26924 16352
rect 26604 15264 26924 16288
rect 26604 15200 26612 15264
rect 26676 15200 26692 15264
rect 26756 15200 26772 15264
rect 26836 15200 26852 15264
rect 26916 15200 26924 15264
rect 26604 14176 26924 15200
rect 26604 14112 26612 14176
rect 26676 14112 26692 14176
rect 26756 14112 26772 14176
rect 26836 14112 26852 14176
rect 26916 14112 26924 14176
rect 26604 13088 26924 14112
rect 26604 13024 26612 13088
rect 26676 13024 26692 13088
rect 26756 13024 26772 13088
rect 26836 13024 26852 13088
rect 26916 13024 26924 13088
rect 26604 12000 26924 13024
rect 26604 11936 26612 12000
rect 26676 11936 26692 12000
rect 26756 11936 26772 12000
rect 26836 11936 26852 12000
rect 26916 11936 26924 12000
rect 26604 10912 26924 11936
rect 26604 10848 26612 10912
rect 26676 10848 26692 10912
rect 26756 10848 26772 10912
rect 26836 10848 26852 10912
rect 26916 10848 26924 10912
rect 26604 9824 26924 10848
rect 26604 9760 26612 9824
rect 26676 9760 26692 9824
rect 26756 9760 26772 9824
rect 26836 9760 26852 9824
rect 26916 9760 26924 9824
rect 26604 8736 26924 9760
rect 26604 8672 26612 8736
rect 26676 8672 26692 8736
rect 26756 8672 26772 8736
rect 26836 8672 26852 8736
rect 26916 8672 26924 8736
rect 26604 7648 26924 8672
rect 26604 7584 26612 7648
rect 26676 7584 26692 7648
rect 26756 7584 26772 7648
rect 26836 7584 26852 7648
rect 26916 7584 26924 7648
rect 26604 6560 26924 7584
rect 26604 6496 26612 6560
rect 26676 6496 26692 6560
rect 26756 6496 26772 6560
rect 26836 6496 26852 6560
rect 26916 6496 26924 6560
rect 26604 5472 26924 6496
rect 26604 5408 26612 5472
rect 26676 5408 26692 5472
rect 26756 5408 26772 5472
rect 26836 5408 26852 5472
rect 26916 5408 26924 5472
rect 26604 4384 26924 5408
rect 26604 4320 26612 4384
rect 26676 4320 26692 4384
rect 26756 4320 26772 4384
rect 26836 4320 26852 4384
rect 26916 4320 26924 4384
rect 26604 3296 26924 4320
rect 26604 3232 26612 3296
rect 26676 3232 26692 3296
rect 26756 3232 26772 3296
rect 26836 3232 26852 3296
rect 26916 3232 26924 3296
rect 26604 2208 26924 3232
rect 26604 2144 26612 2208
rect 26676 2144 26692 2208
rect 26756 2144 26772 2208
rect 26836 2144 26852 2208
rect 26916 2144 26924 2208
rect 26604 2128 26924 2144
use sky130_fd_sc_hd__and2_1  _00_
timestamp -25199
transform 1 0 26956 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _01_
timestamp -25199
transform -1 0 26864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _02_
timestamp -25199
transform 1 0 26956 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _03_
timestamp -25199
transform 1 0 26956 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _04_
timestamp -25199
transform 1 0 26956 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _05_
timestamp -25199
transform 1 0 26864 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _06_
timestamp -25199
transform -1 0 27784 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _07_
timestamp -25199
transform -1 0 27784 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _08_
timestamp -25199
transform -1 0 27784 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _09_
timestamp -25199
transform -1 0 27784 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _10_
timestamp -25199
transform -1 0 27784 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _11_
timestamp -25199
transform -1 0 27784 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp -25199
transform -1 0 27784 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _13_
timestamp -25199
transform -1 0 27784 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _14_
timestamp -25199
transform -1 0 27784 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp -25199
transform -1 0 27784 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -25199
transform -1 0 27692 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636943256
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636943256
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -25199
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636943256
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636943256
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -25199
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636943256
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636943256
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -25199
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636943256
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636943256
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -25199
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636943256
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636943256
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -25199
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636943256
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636943256
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -25199
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636943256
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636943256
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -25199
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636943256
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636943256
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -25199
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636943256
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636943256
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -25199
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636943256
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636943256
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -25199
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636943256
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_293
timestamp -25199
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636943256
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636943256
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636943256
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636943256
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp -25199
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -25199
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636943256
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636943256
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636943256
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636943256
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp -25199
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -25199
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636943256
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636943256
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636943256
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636943256
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp -25199
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -25199
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636943256
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636943256
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636943256
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636943256
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp -25199
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp -25199
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636943256
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636943256
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636943256
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636943256
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp -25199
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp -25199
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636943256
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636943256
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636943256
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -25199
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636943256
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636943256
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636943256
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636943256
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp -25199
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -25199
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636943256
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636943256
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636943256
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636943256
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp -25199
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -25199
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636943256
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636943256
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636943256
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636943256
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp -25199
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp -25199
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636943256
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636943256
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636943256
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636943256
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp -25199
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp -25199
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636943256
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636943256
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636943256
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_289
timestamp -25199
transform 1 0 27692 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_297
timestamp -25199
transform 1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636943256
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636943256
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636943256
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636943256
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp -25199
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -25199
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636943256
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636943256
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636943256
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636943256
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp -25199
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -25199
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636943256
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636943256
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636943256
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636943256
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp -25199
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -25199
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636943256
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636943256
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636943256
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636943256
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp -25199
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp -25199
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636943256
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636943256
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636943256
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636943256
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp -25199
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp -25199
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636943256
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp -25199
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636943256
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636943256
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -25199
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636943256
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636943256
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636943256
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636943256
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp -25199
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -25199
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636943256
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636943256
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636943256
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636943256
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp -25199
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp -25199
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636943256
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636943256
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636943256
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636943256
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp -25199
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp -25199
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636943256
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636943256
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636943256
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636943256
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp -25199
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp -25199
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636943256
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636943256
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636943256
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_289
timestamp -25199
transform 1 0 27692 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636943256
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636943256
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636943256
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636943256
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp -25199
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp -25199
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636943256
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636943256
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636943256
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636943256
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp -25199
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -25199
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636943256
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636943256
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636943256
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636943256
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp -25199
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -25199
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636943256
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636943256
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636943256
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636943256
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp -25199
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp -25199
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636943256
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636943256
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636943256
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636943256
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp -25199
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp -25199
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636943256
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp -25199
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636943256
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636943256
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -25199
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636943256
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636943256
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636943256
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636943256
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp -25199
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp -25199
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636943256
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636943256
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636943256
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636943256
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp -25199
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp -25199
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636943256
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636943256
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636943256
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636943256
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp -25199
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp -25199
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636943256
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636943256
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1636943256
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1636943256
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp -25199
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp -25199
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636943256
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636943256
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_277
timestamp -25199
transform 1 0 26588 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_285
timestamp -25199
transform 1 0 27324 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_290
timestamp -25199
transform 1 0 27784 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_298
timestamp -25199
transform 1 0 28520 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636943256
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636943256
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636943256
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636943256
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp -25199
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -25199
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636943256
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636943256
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636943256
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636943256
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp -25199
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp -25199
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636943256
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636943256
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1636943256
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1636943256
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp -25199
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -25199
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636943256
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636943256
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636943256
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1636943256
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp -25199
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp -25199
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636943256
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636943256
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636943256
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1636943256
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp -25199
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp -25199
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636943256
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636943256
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636943256
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -25199
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636943256
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636943256
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636943256
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636943256
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp -25199
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp -25199
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636943256
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1636943256
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1636943256
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1636943256
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp -25199
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp -25199
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636943256
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636943256
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636943256
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1636943256
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp -25199
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp -25199
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636943256
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636943256
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1636943256
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1636943256
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp -25199
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp -25199
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636943256
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1636943256
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1636943256
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_289
timestamp -25199
transform 1 0 27692 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_297
timestamp -25199
transform 1 0 28428 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636943256
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636943256
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636943256
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1636943256
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp -25199
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -25199
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636943256
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636943256
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636943256
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1636943256
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp -25199
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp -25199
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636943256
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636943256
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1636943256
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1636943256
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp -25199
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp -25199
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636943256
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1636943256
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1636943256
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1636943256
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp -25199
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp -25199
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636943256
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1636943256
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1636943256
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1636943256
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp -25199
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp -25199
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636943256
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp -25199
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_9
timestamp 1636943256
transform 1 0 1932 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp -25199
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -25199
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636943256
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636943256
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636943256
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1636943256
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp -25199
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp -25199
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636943256
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1636943256
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1636943256
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1636943256
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp -25199
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp -25199
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636943256
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1636943256
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1636943256
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1636943256
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp -25199
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp -25199
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1636943256
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1636943256
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1636943256
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1636943256
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp -25199
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp -25199
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1636943256
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1636943256
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1636943256
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_289
timestamp -25199
transform 1 0 27692 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636943256
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636943256
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636943256
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1636943256
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp -25199
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp -25199
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636943256
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1636943256
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1636943256
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1636943256
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp -25199
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp -25199
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1636943256
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1636943256
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1636943256
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1636943256
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp -25199
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp -25199
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1636943256
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1636943256
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1636943256
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1636943256
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp -25199
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp -25199
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1636943256
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1636943256
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1636943256
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1636943256
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp -25199
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp -25199
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1636943256
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp -25199
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636943256
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636943256
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp -25199
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636943256
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636943256
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1636943256
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1636943256
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp -25199
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp -25199
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1636943256
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1636943256
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1636943256
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1636943256
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp -25199
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp -25199
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1636943256
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1636943256
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1636943256
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1636943256
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp -25199
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp -25199
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1636943256
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1636943256
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1636943256
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1636943256
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp -25199
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp -25199
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1636943256
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1636943256
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_277
timestamp -25199
transform 1 0 26588 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_285
timestamp -25199
transform 1 0 27324 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_290
timestamp -25199
transform 1 0 27784 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_298
timestamp -25199
transform 1 0 28520 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636943256
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636943256
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636943256
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1636943256
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp -25199
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp -25199
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636943256
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1636943256
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1636943256
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1636943256
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp -25199
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp -25199
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1636943256
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1636943256
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1636943256
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1636943256
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp -25199
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp -25199
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1636943256
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1636943256
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1636943256
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1636943256
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp -25199
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp -25199
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1636943256
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1636943256
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1636943256
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1636943256
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp -25199
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp -25199
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_281
timestamp -25199
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_290
timestamp -25199
transform 1 0 27784 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636943256
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636943256
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp -25199
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636943256
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636943256
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1636943256
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1636943256
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp -25199
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp -25199
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1636943256
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1636943256
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1636943256
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1636943256
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp -25199
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp -25199
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1636943256
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1636943256
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1636943256
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1636943256
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp -25199
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp -25199
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1636943256
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1636943256
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1636943256
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1636943256
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp -25199
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp -25199
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1636943256
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1636943256
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1636943256
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_289
timestamp -25199
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp -25199
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636943256
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636943256
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636943256
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1636943256
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp -25199
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp -25199
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636943256
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1636943256
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1636943256
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1636943256
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp -25199
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp -25199
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1636943256
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1636943256
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1636943256
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1636943256
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp -25199
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp -25199
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1636943256
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1636943256
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1636943256
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1636943256
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp -25199
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp -25199
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1636943256
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1636943256
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1636943256
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1636943256
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_273
timestamp -25199
transform 1 0 26220 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_294
timestamp -25199
transform 1 0 28152 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_298
timestamp -25199
transform 1 0 28520 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636943256
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636943256
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp -25199
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636943256
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1636943256
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1636943256
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1636943256
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp -25199
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp -25199
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1636943256
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1636943256
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1636943256
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1636943256
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp -25199
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp -25199
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1636943256
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1636943256
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1636943256
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1636943256
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp -25199
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp -25199
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1636943256
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1636943256
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1636943256
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1636943256
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp -25199
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp -25199
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1636943256
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1636943256
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1636943256
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_289
timestamp -25199
transform 1 0 27692 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636943256
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1636943256
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1636943256
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1636943256
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp -25199
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp -25199
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636943256
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1636943256
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1636943256
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1636943256
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp -25199
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp -25199
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1636943256
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1636943256
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1636943256
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1636943256
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp -25199
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp -25199
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1636943256
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1636943256
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1636943256
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1636943256
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp -25199
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp -25199
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1636943256
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1636943256
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1636943256
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1636943256
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp -25199
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp -25199
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_281
timestamp -25199
transform 1 0 26956 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_290
timestamp -25199
transform 1 0 27784 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_298
timestamp -25199
transform 1 0 28520 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636943256
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636943256
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp -25199
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636943256
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636943256
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1636943256
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1636943256
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp -25199
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp -25199
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1636943256
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1636943256
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1636943256
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1636943256
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp -25199
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp -25199
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1636943256
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1636943256
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1636943256
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1636943256
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp -25199
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp -25199
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1636943256
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1636943256
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1636943256
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1636943256
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp -25199
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp -25199
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1636943256
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1636943256
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1636943256
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_289
timestamp -25199
transform 1 0 27692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_297
timestamp -25199
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636943256
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636943256
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1636943256
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1636943256
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp -25199
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp -25199
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636943256
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1636943256
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1636943256
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1636943256
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp -25199
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp -25199
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1636943256
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1636943256
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1636943256
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1636943256
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp -25199
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp -25199
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1636943256
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1636943256
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1636943256
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1636943256
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp -25199
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp -25199
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1636943256
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1636943256
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1636943256
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1636943256
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp -25199
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp -25199
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_286
timestamp -25199
transform 1 0 27416 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_292
timestamp -25199
transform 1 0 27968 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636943256
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1636943256
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp -25199
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636943256
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1636943256
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1636943256
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1636943256
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp -25199
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp -25199
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1636943256
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1636943256
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1636943256
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1636943256
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp -25199
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp -25199
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1636943256
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1636943256
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1636943256
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1636943256
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp -25199
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp -25199
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1636943256
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1636943256
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1636943256
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1636943256
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp -25199
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp -25199
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1636943256
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1636943256
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_277
timestamp -25199
transform 1 0 26588 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_285
timestamp -25199
transform 1 0 27324 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_290
timestamp -25199
transform 1 0 27784 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_298
timestamp -25199
transform 1 0 28520 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636943256
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636943256
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1636943256
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1636943256
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp -25199
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp -25199
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1636943256
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1636943256
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1636943256
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1636943256
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp -25199
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp -25199
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1636943256
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1636943256
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1636943256
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1636943256
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp -25199
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp -25199
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1636943256
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1636943256
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1636943256
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1636943256
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp -25199
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp -25199
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1636943256
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1636943256
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1636943256
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1636943256
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp -25199
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp -25199
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1636943256
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_293
timestamp -25199
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636943256
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636943256
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp -25199
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636943256
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1636943256
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1636943256
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1636943256
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp -25199
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp -25199
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1636943256
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1636943256
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1636943256
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1636943256
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp -25199
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp -25199
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1636943256
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1636943256
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1636943256
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1636943256
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp -25199
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp -25199
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1636943256
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1636943256
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1636943256
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1636943256
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp -25199
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp -25199
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1636943256
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1636943256
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1636943256
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_289
timestamp -25199
transform 1 0 27692 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636943256
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636943256
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1636943256
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1636943256
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp -25199
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp -25199
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1636943256
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1636943256
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1636943256
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1636943256
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp -25199
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp -25199
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1636943256
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1636943256
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1636943256
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1636943256
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp -25199
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp -25199
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1636943256
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1636943256
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1636943256
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1636943256
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp -25199
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp -25199
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1636943256
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1636943256
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1636943256
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1636943256
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp -25199
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp -25199
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1636943256
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_293
timestamp -25199
transform 1 0 28060 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636943256
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636943256
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp -25199
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636943256
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1636943256
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1636943256
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1636943256
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp -25199
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp -25199
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1636943256
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1636943256
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1636943256
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1636943256
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp -25199
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp -25199
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1636943256
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1636943256
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1636943256
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1636943256
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp -25199
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp -25199
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1636943256
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1636943256
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1636943256
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1636943256
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp -25199
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp -25199
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1636943256
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1636943256
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1636943256
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_289
timestamp -25199
transform 1 0 27692 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1636943256
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1636943256
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1636943256
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1636943256
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp -25199
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp -25199
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636943256
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1636943256
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1636943256
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1636943256
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp -25199
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp -25199
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1636943256
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1636943256
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1636943256
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1636943256
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp -25199
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp -25199
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1636943256
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1636943256
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1636943256
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1636943256
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp -25199
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp -25199
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1636943256
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1636943256
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1636943256
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1636943256
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp -25199
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp -25199
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_294
timestamp -25199
transform 1 0 28152 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_298
timestamp -25199
transform 1 0 28520 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636943256
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636943256
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp -25199
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636943256
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1636943256
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1636943256
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1636943256
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp -25199
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp -25199
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1636943256
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1636943256
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1636943256
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1636943256
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp -25199
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp -25199
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1636943256
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1636943256
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1636943256
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1636943256
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp -25199
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp -25199
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1636943256
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1636943256
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1636943256
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1636943256
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp -25199
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp -25199
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1636943256
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1636943256
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_277
timestamp -25199
transform 1 0 26588 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_286
timestamp 1636943256
transform 1 0 27416 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_298
timestamp -25199
transform 1 0 28520 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636943256
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1636943256
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1636943256
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1636943256
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp -25199
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp -25199
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1636943256
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1636943256
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1636943256
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1636943256
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp -25199
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp -25199
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1636943256
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1636943256
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1636943256
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1636943256
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp -25199
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp -25199
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1636943256
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1636943256
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1636943256
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1636943256
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp -25199
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp -25199
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1636943256
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1636943256
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1636943256
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1636943256
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp -25199
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp -25199
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_289
timestamp -25199
transform 1 0 27692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_297
timestamp -25199
transform 1 0 28428 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636943256
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636943256
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp -25199
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636943256
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636943256
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1636943256
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1636943256
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp -25199
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp -25199
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1636943256
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1636943256
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1636943256
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1636943256
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp -25199
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp -25199
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1636943256
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1636943256
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1636943256
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1636943256
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp -25199
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp -25199
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1636943256
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1636943256
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1636943256
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1636943256
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp -25199
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp -25199
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1636943256
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1636943256
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1636943256
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_289
timestamp -25199
transform 1 0 27692 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636943256
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1636943256
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1636943256
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1636943256
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp -25199
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp -25199
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636943256
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1636943256
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1636943256
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1636943256
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp -25199
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp -25199
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1636943256
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1636943256
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1636943256
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1636943256
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp -25199
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp -25199
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1636943256
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1636943256
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1636943256
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1636943256
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp -25199
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp -25199
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1636943256
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1636943256
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1636943256
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1636943256
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp -25199
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp -25199
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp -25199
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_290
timestamp -25199
transform 1 0 27784 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_298
timestamp -25199
transform 1 0 28520 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636943256
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636943256
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp -25199
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1636943256
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1636943256
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1636943256
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1636943256
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp -25199
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp -25199
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1636943256
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1636943256
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1636943256
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1636943256
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp -25199
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp -25199
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1636943256
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1636943256
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1636943256
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1636943256
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp -25199
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp -25199
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1636943256
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1636943256
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1636943256
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1636943256
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp -25199
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp -25199
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1636943256
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1636943256
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_277
timestamp -25199
transform 1 0 26588 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_285
timestamp -25199
transform 1 0 27324 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_290
timestamp -25199
transform 1 0 27784 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_298
timestamp -25199
transform 1 0 28520 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636943256
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636943256
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1636943256
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1636943256
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp -25199
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp -25199
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1636943256
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1636943256
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1636943256
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1636943256
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp -25199
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp -25199
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1636943256
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1636943256
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1636943256
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1636943256
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp -25199
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp -25199
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1636943256
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1636943256
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1636943256
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1636943256
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp -25199
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp -25199
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1636943256
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1636943256
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1636943256
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1636943256
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp -25199
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp -25199
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1636943256
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636943256
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1636943256
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp -25199
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636943256
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1636943256
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1636943256
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1636943256
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp -25199
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp -25199
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1636943256
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1636943256
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1636943256
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1636943256
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp -25199
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp -25199
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1636943256
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1636943256
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1636943256
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1636943256
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp -25199
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp -25199
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1636943256
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1636943256
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1636943256
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1636943256
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp -25199
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp -25199
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1636943256
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1636943256
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1636943256
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_289
timestamp -25199
transform 1 0 27692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp -25199
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636943256
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1636943256
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1636943256
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1636943256
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp -25199
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp -25199
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1636943256
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1636943256
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1636943256
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1636943256
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp -25199
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp -25199
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1636943256
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1636943256
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1636943256
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1636943256
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp -25199
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp -25199
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1636943256
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1636943256
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1636943256
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1636943256
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp -25199
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp -25199
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1636943256
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1636943256
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1636943256
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1636943256
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp -25199
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp -25199
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1636943256
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_293
timestamp -25199
transform 1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636943256
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636943256
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp -25199
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1636943256
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1636943256
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1636943256
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1636943256
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp -25199
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp -25199
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1636943256
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1636943256
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1636943256
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1636943256
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp -25199
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp -25199
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1636943256
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1636943256
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1636943256
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1636943256
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp -25199
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp -25199
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1636943256
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1636943256
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1636943256
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1636943256
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp -25199
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp -25199
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1636943256
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1636943256
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1636943256
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_289
timestamp -25199
transform 1 0 27692 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1636943256
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1636943256
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1636943256
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1636943256
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp -25199
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp -25199
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1636943256
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1636943256
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1636943256
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1636943256
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp -25199
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp -25199
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1636943256
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1636943256
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1636943256
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1636943256
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp -25199
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp -25199
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1636943256
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1636943256
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1636943256
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1636943256
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp -25199
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp -25199
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1636943256
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1636943256
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1636943256
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1636943256
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp -25199
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp -25199
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1636943256
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_293
timestamp -25199
transform 1 0 28060 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636943256
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636943256
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp -25199
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1636943256
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1636943256
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1636943256
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1636943256
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp -25199
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp -25199
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1636943256
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1636943256
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1636943256
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1636943256
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp -25199
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp -25199
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1636943256
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1636943256
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1636943256
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1636943256
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp -25199
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp -25199
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1636943256
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1636943256
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1636943256
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1636943256
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp -25199
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp -25199
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1636943256
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1636943256
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_277
timestamp -25199
transform 1 0 26588 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_285
timestamp -25199
transform 1 0 27324 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_290
timestamp -25199
transform 1 0 27784 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_298
timestamp -25199
transform 1 0 28520 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_9
timestamp 1636943256
transform 1 0 1932 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_21
timestamp 1636943256
transform 1 0 3036 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_33
timestamp 1636943256
transform 1 0 4140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_45
timestamp -25199
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp -25199
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1636943256
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1636943256
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1636943256
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1636943256
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp -25199
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp -25199
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1636943256
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1636943256
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1636943256
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1636943256
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp -25199
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp -25199
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1636943256
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1636943256
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1636943256
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1636943256
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp -25199
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp -25199
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1636943256
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1636943256
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1636943256
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1636943256
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp -25199
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp -25199
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_281
timestamp -25199
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_37_290
timestamp -25199
transform 1 0 27784 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636943256
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636943256
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp -25199
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1636943256
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1636943256
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1636943256
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1636943256
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp -25199
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp -25199
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1636943256
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1636943256
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1636943256
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1636943256
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp -25199
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp -25199
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1636943256
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1636943256
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1636943256
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1636943256
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp -25199
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp -25199
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1636943256
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1636943256
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1636943256
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1636943256
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp -25199
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp -25199
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1636943256
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1636943256
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1636943256
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_289
timestamp -25199
transform 1 0 27692 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_297
timestamp -25199
transform 1 0 28428 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1636943256
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1636943256
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1636943256
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1636943256
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp -25199
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp -25199
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1636943256
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1636943256
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1636943256
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1636943256
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp -25199
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp -25199
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1636943256
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1636943256
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1636943256
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1636943256
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp -25199
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp -25199
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1636943256
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1636943256
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1636943256
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1636943256
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp -25199
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp -25199
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1636943256
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1636943256
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1636943256
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1636943256
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp -25199
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp -25199
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1636943256
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_293
timestamp -25199
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1636943256
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1636943256
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp -25199
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636943256
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1636943256
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1636943256
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1636943256
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp -25199
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp -25199
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1636943256
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1636943256
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1636943256
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1636943256
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp -25199
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp -25199
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1636943256
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1636943256
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1636943256
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1636943256
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp -25199
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp -25199
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1636943256
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1636943256
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1636943256
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1636943256
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp -25199
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp -25199
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1636943256
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1636943256
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_277
timestamp -25199
transform 1 0 26588 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_285
timestamp -25199
transform 1 0 27324 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_290
timestamp -25199
transform 1 0 27784 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636943256
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1636943256
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1636943256
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1636943256
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp -25199
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp -25199
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1636943256
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1636943256
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1636943256
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1636943256
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp -25199
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp -25199
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1636943256
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1636943256
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1636943256
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1636943256
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp -25199
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp -25199
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1636943256
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1636943256
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1636943256
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1636943256
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp -25199
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp -25199
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1636943256
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1636943256
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1636943256
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1636943256
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp -25199
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp -25199
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1636943256
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp -25199
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636943256
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1636943256
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp -25199
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636943256
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1636943256
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1636943256
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1636943256
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp -25199
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp -25199
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1636943256
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1636943256
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1636943256
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1636943256
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp -25199
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp -25199
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1636943256
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1636943256
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1636943256
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1636943256
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp -25199
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp -25199
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1636943256
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1636943256
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1636943256
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1636943256
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp -25199
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp -25199
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1636943256
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1636943256
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1636943256
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_289
timestamp -25199
transform 1 0 27692 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_297
timestamp -25199
transform 1 0 28428 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636943256
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636943256
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1636943256
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1636943256
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp -25199
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp -25199
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1636943256
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1636943256
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1636943256
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1636943256
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp -25199
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp -25199
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1636943256
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1636943256
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1636943256
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1636943256
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp -25199
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp -25199
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1636943256
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1636943256
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1636943256
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1636943256
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp -25199
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp -25199
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1636943256
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1636943256
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1636943256
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1636943256
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp -25199
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp -25199
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1636943256
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1636943256
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1636943256
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp -25199
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1636943256
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1636943256
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1636943256
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1636943256
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp -25199
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp -25199
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1636943256
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1636943256
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1636943256
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1636943256
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp -25199
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp -25199
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1636943256
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1636943256
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1636943256
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1636943256
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp -25199
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp -25199
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1636943256
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1636943256
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1636943256
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1636943256
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp -25199
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp -25199
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1636943256
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1636943256
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1636943256
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_289
timestamp -25199
transform 1 0 27692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_297
timestamp -25199
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1636943256
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1636943256
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1636943256
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1636943256
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp -25199
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp -25199
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1636943256
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1636943256
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1636943256
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1636943256
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp -25199
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp -25199
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1636943256
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1636943256
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1636943256
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1636943256
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp -25199
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp -25199
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1636943256
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1636943256
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1636943256
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1636943256
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp -25199
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp -25199
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1636943256
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1636943256
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1636943256
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1636943256
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp -25199
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp -25199
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1636943256
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_293
timestamp -25199
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636943256
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636943256
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp -25199
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1636943256
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1636943256
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_53
timestamp -25199
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_57
timestamp 1636943256
transform 1 0 6348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_69
timestamp 1636943256
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp -25199
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1636943256
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1636943256
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_109
timestamp -25199
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_113
timestamp 1636943256
transform 1 0 11500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_125
timestamp 1636943256
transform 1 0 12604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp -25199
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1636943256
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1636943256
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_165
timestamp -25199
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_169
timestamp 1636943256
transform 1 0 16652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_181
timestamp 1636943256
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_193
timestamp -25199
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1636943256
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1636943256
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_221
timestamp -25199
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_225
timestamp 1636943256
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_237
timestamp 1636943256
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp -25199
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1636943256
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1636943256
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_277
timestamp -25199
transform 1 0 26588 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_281
timestamp 1636943256
transform 1 0 26956 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp -25199
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp -25199
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output3
timestamp -25199
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output4
timestamp -25199
transform 1 0 28060 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output5
timestamp -25199
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output6
timestamp -25199
transform 1 0 28060 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output7
timestamp -25199
transform 1 0 28060 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output8
timestamp -25199
transform 1 0 28060 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output9
timestamp -25199
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output10
timestamp -25199
transform 1 0 28060 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output11
timestamp -25199
transform 1 0 28060 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output12
timestamp -25199
transform 1 0 28060 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output13
timestamp -25199
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output14
timestamp -25199
transform 1 0 28060 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output15
timestamp -25199
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output16
timestamp -25199
transform 1 0 28060 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output17
timestamp -25199
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output18
timestamp -25199
transform 1 0 28060 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_47
timestamp -25199
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -25199
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_48
timestamp -25199
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -25199
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_49
timestamp -25199
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -25199
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_50
timestamp -25199
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -25199
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_51
timestamp -25199
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -25199
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_52
timestamp -25199
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -25199
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_53
timestamp -25199
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -25199
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_54
timestamp -25199
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -25199
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_55
timestamp -25199
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -25199
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_56
timestamp -25199
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -25199
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_57
timestamp -25199
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -25199
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_58
timestamp -25199
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -25199
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_59
timestamp -25199
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -25199
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_60
timestamp -25199
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -25199
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_61
timestamp -25199
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -25199
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_62
timestamp -25199
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -25199
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_63
timestamp -25199
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -25199
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_64
timestamp -25199
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -25199
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_65
timestamp -25199
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -25199
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_66
timestamp -25199
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -25199
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_67
timestamp -25199
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -25199
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_68
timestamp -25199
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -25199
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_69
timestamp -25199
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -25199
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_70
timestamp -25199
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -25199
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_71
timestamp -25199
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -25199
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_72
timestamp -25199
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp -25199
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_73
timestamp -25199
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp -25199
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_74
timestamp -25199
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp -25199
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_75
timestamp -25199
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp -25199
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_76
timestamp -25199
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp -25199
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_77
timestamp -25199
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp -25199
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_78
timestamp -25199
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp -25199
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_79
timestamp -25199
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp -25199
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_80
timestamp -25199
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp -25199
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_81
timestamp -25199
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp -25199
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_82
timestamp -25199
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp -25199
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_83
timestamp -25199
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp -25199
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_84
timestamp -25199
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp -25199
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_85
timestamp -25199
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp -25199
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_86
timestamp -25199
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp -25199
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_87
timestamp -25199
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp -25199
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_88
timestamp -25199
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp -25199
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_89
timestamp -25199
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp -25199
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_90
timestamp -25199
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp -25199
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_91
timestamp -25199
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp -25199
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_92
timestamp -25199
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp -25199
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_93
timestamp -25199
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp -25199
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_94
timestamp -25199
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_95
timestamp -25199
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_96
timestamp -25199
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_97
timestamp -25199
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_98
timestamp -25199
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_99
timestamp -25199
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_100
timestamp -25199
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_101
timestamp -25199
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_102
timestamp -25199
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_103
timestamp -25199
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_104
timestamp -25199
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_105
timestamp -25199
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_106
timestamp -25199
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_107
timestamp -25199
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_108
timestamp -25199
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_109
timestamp -25199
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_110
timestamp -25199
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_111
timestamp -25199
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_112
timestamp -25199
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_113
timestamp -25199
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_114
timestamp -25199
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_115
timestamp -25199
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_116
timestamp -25199
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_117
timestamp -25199
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_118
timestamp -25199
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_119
timestamp -25199
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_120
timestamp -25199
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_121
timestamp -25199
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_122
timestamp -25199
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_123
timestamp -25199
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_124
timestamp -25199
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_125
timestamp -25199
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_126
timestamp -25199
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_127
timestamp -25199
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_128
timestamp -25199
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_129
timestamp -25199
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_130
timestamp -25199
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_131
timestamp -25199
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_132
timestamp -25199
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_133
timestamp -25199
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_134
timestamp -25199
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_135
timestamp -25199
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_136
timestamp -25199
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_137
timestamp -25199
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_138
timestamp -25199
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_139
timestamp -25199
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_140
timestamp -25199
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_141
timestamp -25199
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_142
timestamp -25199
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_143
timestamp -25199
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_144
timestamp -25199
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_145
timestamp -25199
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_146
timestamp -25199
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_147
timestamp -25199
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_148
timestamp -25199
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_149
timestamp -25199
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_150
timestamp -25199
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_151
timestamp -25199
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_152
timestamp -25199
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_153
timestamp -25199
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_154
timestamp -25199
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_155
timestamp -25199
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_156
timestamp -25199
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_157
timestamp -25199
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_158
timestamp -25199
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_159
timestamp -25199
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_160
timestamp -25199
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_161
timestamp -25199
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_162
timestamp -25199
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_163
timestamp -25199
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_164
timestamp -25199
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_165
timestamp -25199
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_166
timestamp -25199
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_167
timestamp -25199
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_168
timestamp -25199
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_169
timestamp -25199
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_170
timestamp -25199
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_171
timestamp -25199
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_172
timestamp -25199
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_173
timestamp -25199
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_174
timestamp -25199
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_175
timestamp -25199
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_176
timestamp -25199
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_177
timestamp -25199
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_178
timestamp -25199
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_179
timestamp -25199
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_180
timestamp -25199
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_181
timestamp -25199
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_182
timestamp -25199
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_183
timestamp -25199
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_184
timestamp -25199
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_185
timestamp -25199
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_186
timestamp -25199
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_187
timestamp -25199
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_188
timestamp -25199
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_189
timestamp -25199
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_190
timestamp -25199
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_191
timestamp -25199
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_192
timestamp -25199
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_193
timestamp -25199
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_194
timestamp -25199
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_195
timestamp -25199
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_196
timestamp -25199
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_197
timestamp -25199
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_198
timestamp -25199
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_199
timestamp -25199
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_200
timestamp -25199
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_201
timestamp -25199
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_202
timestamp -25199
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_203
timestamp -25199
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_204
timestamp -25199
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_205
timestamp -25199
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_206
timestamp -25199
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_207
timestamp -25199
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_208
timestamp -25199
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_209
timestamp -25199
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_210
timestamp -25199
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_211
timestamp -25199
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_212
timestamp -25199
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_213
timestamp -25199
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_214
timestamp -25199
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_215
timestamp -25199
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_216
timestamp -25199
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_217
timestamp -25199
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_218
timestamp -25199
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_219
timestamp -25199
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_220
timestamp -25199
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_221
timestamp -25199
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_222
timestamp -25199
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_223
timestamp -25199
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_224
timestamp -25199
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_225
timestamp -25199
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_226
timestamp -25199
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_227
timestamp -25199
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_228
timestamp -25199
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_229
timestamp -25199
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_230
timestamp -25199
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_231
timestamp -25199
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_232
timestamp -25199
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_233
timestamp -25199
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_234
timestamp -25199
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_235
timestamp -25199
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_236
timestamp -25199
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_237
timestamp -25199
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_238
timestamp -25199
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_239
timestamp -25199
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_240
timestamp -25199
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_241
timestamp -25199
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_242
timestamp -25199
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_243
timestamp -25199
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_244
timestamp -25199
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_245
timestamp -25199
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_246
timestamp -25199
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_247
timestamp -25199
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_248
timestamp -25199
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_249
timestamp -25199
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_250
timestamp -25199
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_251
timestamp -25199
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_252
timestamp -25199
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp -25199
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_254
timestamp -25199
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_255
timestamp -25199
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_256
timestamp -25199
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_257
timestamp -25199
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp -25199
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_259
timestamp -25199
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_260
timestamp -25199
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_261
timestamp -25199
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_262
timestamp -25199
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp -25199
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_264
timestamp -25199
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp -25199
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_266
timestamp -25199
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_267
timestamp -25199
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp -25199
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_269
timestamp -25199
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_270
timestamp -25199
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_271
timestamp -25199
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_272
timestamp -25199
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp -25199
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_274
timestamp -25199
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_275
timestamp -25199
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_276
timestamp -25199
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_277
timestamp -25199
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp -25199
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_279
timestamp -25199
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_280
timestamp -25199
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_281
timestamp -25199
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_282
timestamp -25199
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp -25199
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_284
timestamp -25199
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_285
timestamp -25199
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_286
timestamp -25199
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_287
timestamp -25199
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp -25199
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_289
timestamp -25199
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_290
timestamp -25199
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_291
timestamp -25199
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_292
timestamp -25199
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp -25199
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_294
timestamp -25199
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_295
timestamp -25199
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_296
timestamp -25199
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_297
timestamp -25199
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_298
timestamp -25199
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_299
timestamp -25199
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_300
timestamp -25199
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_301
timestamp -25199
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_302
timestamp -25199
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_303
timestamp -25199
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_304
timestamp -25199
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_305
timestamp -25199
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_306
timestamp -25199
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_307
timestamp -25199
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_308
timestamp -25199
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_309
timestamp -25199
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_310
timestamp -25199
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_311
timestamp -25199
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_312
timestamp -25199
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_313
timestamp -25199
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_314
timestamp -25199
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_315
timestamp -25199
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_316
timestamp -25199
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_317
timestamp -25199
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_318
timestamp -25199
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_319
timestamp -25199
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_320
timestamp -25199
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_321
timestamp -25199
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_322
timestamp -25199
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_323
timestamp -25199
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_324
timestamp -25199
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_325
timestamp -25199
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_326
timestamp -25199
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_327
timestamp -25199
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_328
timestamp -25199
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_329
timestamp -25199
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_330
timestamp -25199
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_331
timestamp -25199
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_332
timestamp -25199
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_333
timestamp -25199
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_334
timestamp -25199
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_335
timestamp -25199
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_336
timestamp -25199
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_337
timestamp -25199
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_338
timestamp -25199
transform 1 0 26864 0 1 27200
box -38 -48 130 592
<< labels >>
flabel metal3 s 29200 2456 30000 2576 0 FreeSans 480 0 0 0 bm_s0_s0_o[0]
port 0 nsew signal output
flabel metal3 s 29200 4088 30000 4208 0 FreeSans 480 0 0 0 bm_s0_s0_o[1]
port 1 nsew signal output
flabel metal3 s 29200 5720 30000 5840 0 FreeSans 480 0 0 0 bm_s0_s2_o[0]
port 2 nsew signal output
flabel metal3 s 29200 7352 30000 7472 0 FreeSans 480 0 0 0 bm_s0_s2_o[1]
port 3 nsew signal output
flabel metal3 s 29200 8984 30000 9104 0 FreeSans 480 0 0 0 bm_s1_s0_o[0]
port 4 nsew signal output
flabel metal3 s 29200 10616 30000 10736 0 FreeSans 480 0 0 0 bm_s1_s0_o[1]
port 5 nsew signal output
flabel metal3 s 29200 12248 30000 12368 0 FreeSans 480 0 0 0 bm_s1_s2_o[0]
port 6 nsew signal output
flabel metal3 s 29200 13880 30000 14000 0 FreeSans 480 0 0 0 bm_s1_s2_o[1]
port 7 nsew signal output
flabel metal3 s 29200 15512 30000 15632 0 FreeSans 480 0 0 0 bm_s2_s1_o[0]
port 8 nsew signal output
flabel metal3 s 29200 17144 30000 17264 0 FreeSans 480 0 0 0 bm_s2_s1_o[1]
port 9 nsew signal output
flabel metal3 s 29200 18776 30000 18896 0 FreeSans 480 0 0 0 bm_s2_s3_o[0]
port 10 nsew signal output
flabel metal3 s 29200 20408 30000 20528 0 FreeSans 480 0 0 0 bm_s2_s3_o[1]
port 11 nsew signal output
flabel metal3 s 29200 22040 30000 22160 0 FreeSans 480 0 0 0 bm_s3_s1_o[0]
port 12 nsew signal output
flabel metal3 s 29200 23672 30000 23792 0 FreeSans 480 0 0 0 bm_s3_s1_o[1]
port 13 nsew signal output
flabel metal3 s 29200 25304 30000 25424 0 FreeSans 480 0 0 0 bm_s3_s3_o[0]
port 14 nsew signal output
flabel metal3 s 29200 26936 30000 27056 0 FreeSans 480 0 0 0 bm_s3_s3_o[1]
port 15 nsew signal output
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 piso_data_i[0]
port 16 nsew signal input
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 piso_data_i[1]
port 17 nsew signal input
flabel metal4 s 1944 2128 2264 27792 0 FreeSans 1920 90 0 0 vccd1
port 18 nsew power bidirectional
flabel metal4 s 9944 2128 10264 27792 0 FreeSans 1920 90 0 0 vccd1
port 18 nsew power bidirectional
flabel metal4 s 17944 2128 18264 27792 0 FreeSans 1920 90 0 0 vccd1
port 18 nsew power bidirectional
flabel metal4 s 25944 2128 26264 27792 0 FreeSans 1920 90 0 0 vccd1
port 18 nsew power bidirectional
flabel metal4 s 2604 2128 2924 27792 0 FreeSans 1920 90 0 0 vssd1
port 19 nsew ground bidirectional
flabel metal4 s 10604 2128 10924 27792 0 FreeSans 1920 90 0 0 vssd1
port 19 nsew ground bidirectional
flabel metal4 s 18604 2128 18924 27792 0 FreeSans 1920 90 0 0 vssd1
port 19 nsew ground bidirectional
flabel metal4 s 26604 2128 26924 27792 0 FreeSans 1920 90 0 0 vssd1
port 19 nsew ground bidirectional
rlabel metal1 14996 27744 14996 27744 0 vccd1
rlabel metal1 14996 27200 14996 27200 0 vssd1
rlabel metal2 28382 2737 28382 2737 0 bm_s0_s0_o[0]
rlabel metal2 28382 4335 28382 4335 0 bm_s0_s0_o[1]
rlabel metal2 28382 6001 28382 6001 0 bm_s0_s2_o[0]
rlabel metal2 28382 7599 28382 7599 0 bm_s0_s2_o[1]
rlabel metal2 28382 9265 28382 9265 0 bm_s1_s0_o[0]
rlabel metal2 28382 10863 28382 10863 0 bm_s1_s0_o[1]
rlabel metal2 28382 12529 28382 12529 0 bm_s1_s2_o[0]
rlabel metal2 28382 14127 28382 14127 0 bm_s1_s2_o[1]
rlabel via2 28382 15555 28382 15555 0 bm_s2_s1_o[0]
rlabel metal2 28382 17391 28382 17391 0 bm_s2_s1_o[1]
rlabel metal2 28382 19091 28382 19091 0 bm_s2_s3_o[0]
rlabel metal2 28382 20655 28382 20655 0 bm_s2_s3_o[1]
rlabel metal2 28382 22321 28382 22321 0 bm_s3_s1_o[0]
rlabel metal2 28382 23919 28382 23919 0 bm_s3_s1_o[1]
rlabel metal2 28382 25585 28382 25585 0 bm_s3_s3_o[0]
rlabel metal2 28382 27183 28382 27183 0 bm_s3_s3_o[1]
rlabel metal1 27094 16694 27094 16694 0 net1
rlabel metal1 27922 13498 27922 13498 0 net10
rlabel metal2 27554 20366 27554 20366 0 net11
rlabel metal1 27738 17646 27738 17646 0 net12
rlabel metal1 27922 18938 27922 18938 0 net13
rlabel metal1 27784 20910 27784 20910 0 net14
rlabel metal1 27922 22202 27922 22202 0 net15
rlabel metal1 27922 22746 27922 22746 0 net16
rlabel metal1 27922 24378 27922 24378 0 net17
rlabel metal1 27692 18394 27692 18394 0 net18
rlabel metal2 1794 19686 1794 19686 0 net2
rlabel metal2 27554 4352 27554 4352 0 net3
rlabel metal1 28152 4590 28152 4590 0 net4
rlabel metal2 27738 6086 27738 6086 0 net5
rlabel metal2 27554 10030 27554 10030 0 net6
rlabel metal2 27738 9350 27738 9350 0 net7
rlabel metal1 27922 9418 27922 9418 0 net8
rlabel metal1 27922 11866 27922 11866 0 net9
rlabel metal3 751 7412 751 7412 0 piso_data_i[0]
rlabel metal3 751 22372 751 22372 0 piso_data_i[1]
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
