* NGSPICE file created from acsu.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

.subckt acsu bm_s0_s0_i[0] bm_s0_s0_i[1] bm_s0_s2_i[0] bm_s0_s2_i[1] bm_s1_s0_i[0]
+ bm_s1_s0_i[1] bm_s1_s2_i[0] bm_s1_s2_i[1] bm_s2_s1_i[0] bm_s2_s1_i[1] bm_s2_s3_i[0]
+ bm_s2_s3_i[1] bm_s3_s1_i[0] bm_s3_s1_i[1] bm_s3_s3_i[0] bm_s3_s3_i[1] dec_bits_o[0]
+ dec_bits_o[1] dec_bits_o[2] dec_bits_o[3] pm_s0_i[0] pm_s0_i[1] pm_s0_i[2] pm_s0_i[3]
+ pm_s0_i[4] pm_s0_i[5] pm_s0_i[6] pm_s0_i[7] pm_s0_o[0] pm_s0_o[1] pm_s0_o[2] pm_s0_o[3]
+ pm_s0_o[4] pm_s0_o[5] pm_s0_o[6] pm_s0_o[7] pm_s1_i[0] pm_s1_i[1] pm_s1_i[2] pm_s1_i[3]
+ pm_s1_i[4] pm_s1_i[5] pm_s1_i[6] pm_s1_i[7] pm_s1_o[0] pm_s1_o[1] pm_s1_o[2] pm_s1_o[3]
+ pm_s1_o[4] pm_s1_o[5] pm_s1_o[6] pm_s1_o[7] pm_s2_i[0] pm_s2_i[1] pm_s2_i[2] pm_s2_i[3]
+ pm_s2_i[4] pm_s2_i[5] pm_s2_i[6] pm_s2_i[7] pm_s2_o[0] pm_s2_o[1] pm_s2_o[2] pm_s2_o[3]
+ pm_s2_o[4] pm_s2_o[5] pm_s2_o[6] pm_s2_o[7] pm_s3_i[0] pm_s3_i[1] pm_s3_i[2] pm_s3_i[3]
+ pm_s3_i[4] pm_s3_i[5] pm_s3_i[6] pm_s3_i[7] pm_s3_o[0] pm_s3_o[1] pm_s3_o[2] pm_s3_o[3]
+ pm_s3_o[4] pm_s3_o[5] pm_s3_o[6] pm_s3_o[7] vccd1 vssd1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_363_ net42 net14 vssd1 vssd1 vccd1 vccd1 _103_ sky130_fd_sc_hd__xnor2_2
X_294_ _020_ _023_ _045_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_432_ net26 net6 vssd1 vssd1 vccd1 vccd1 _163_ sky130_fd_sc_hd__nand2_1
XFILLER_9_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout105 net30 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_2
X_415_ _146_ _150_ _153_ _154_ vssd1 vssd1 vccd1 vccd1 _155_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_20_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_346_ net30 _080_ net31 vssd1 vssd1 vccd1 vccd1 _095_ sky130_fd_sc_hd__a21oi_1
XFILLER_12_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_277_ net39 net100 net94 vssd1 vssd1 vccd1 vccd1 _035_ sky130_fd_sc_hd__and3_1
XFILLER_23_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_329_ net20 net19 _053_ net21 vssd1 vssd1 vccd1 vccd1 _078_ sky130_fd_sc_hd__a31o_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input18_A pm_s0_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 pm_s2_o[6] sky130_fd_sc_hd__buf_4
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 pm_s1_o[3] sky130_fd_sc_hd__buf_4
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 pm_s0_o[0] sky130_fd_sc_hd__buf_4
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_362_ net42 net14 vssd1 vssd1 vccd1 vccd1 _102_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_21_Left_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_293_ _223_ _003_ net91 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__mux2_1
X_431_ _214_ _161_ vssd1 vssd1 vccd1 vccd1 _162_ sky130_fd_sc_hd__xnor2_1
XANTENNA_output49_A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout106 net28 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_20_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_276_ _032_ _033_ vssd1 vssd1 vccd1 vccd1 _034_ sky130_fd_sc_hd__nor2_1
X_414_ net40 _148_ vssd1 vssd1 vccd1 vccd1 _154_ sky130_fd_sc_hd__xor2_1
X_345_ net31 net105 net93 vssd1 vssd1 vccd1 vccd1 _094_ sky130_fd_sc_hd__and3_1
XFILLER_23_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_259_ net45 net97 net99 _220_ vssd1 vssd1 vccd1 vccd1 _017_ sky130_fd_sc_hd__and4_1
XANTENNA_input48_A pm_s3_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_328_ _213_ _214_ _216_ _053_ vssd1 vssd1 vccd1 vccd1 _077_ sky130_fd_sc_hd__or4b_2
XFILLER_9_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_24_Left_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input30_A pm_s1_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 pm_s2_o[7] sky130_fd_sc_hd__buf_4
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 pm_s1_o[4] sky130_fd_sc_hd__buf_4
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 pm_s0_o[1] sky130_fd_sc_hd__buf_4
XFILLER_22_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_292_ _006_ _007_ net91 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__mux2_1
XFILLER_13_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_430_ net111 net1 _160_ _159_ vssd1 vssd1 vccd1 vccd1 _161_ sky130_fd_sc_hd__a31o_1
X_361_ _099_ _100_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__and2b_1
Xfanout107 net27 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_2
XFILLER_12_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_275_ net95 _017_ net47 vssd1 vssd1 vccd1 vccd1 _033_ sky130_fd_sc_hd__a21oi_1
X_413_ net48 _144_ vssd1 vssd1 vccd1 vccd1 _153_ sky130_fd_sc_hd__xnor2_1
X_344_ _091_ _092_ vssd1 vssd1 vccd1 vccd1 _093_ sky130_fd_sc_hd__nor2_1
XFILLER_23_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_258_ _005_ _007_ vssd1 vssd1 vccd1 vccd1 _016_ sky130_fd_sc_hd__nor2_1
X_327_ net20 net19 net21 _053_ vssd1 vssd1 vccd1 vccd1 _076_ sky130_fd_sc_hd__and4_1
XFILLER_15_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input23_A pm_s0_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 pm_s3_o[0] sky130_fd_sc_hd__buf_4
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 pm_s1_o[5] sky130_fd_sc_hd__buf_4
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 pm_s0_o[2] sky130_fd_sc_hd__buf_4
XFILLER_22_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_291_ _008_ net91 _046_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__o21bai_1
XFILLER_13_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_360_ _093_ _097_ net89 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__mux2_1
X_489_ _209_ _210_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__and2b_1
XFILLER_12_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout108 net27 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__buf_1
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_274_ net47 net95 _017_ vssd1 vssd1 vccd1 vccd1 _032_ sky130_fd_sc_hd__and3_1
X_412_ _139_ _143_ _146_ _150_ _151_ vssd1 vssd1 vccd1 vccd1 _152_ sky130_fd_sc_hd__a221o_1
X_343_ net22 _076_ net23 vssd1 vssd1 vccd1 vccd1 _092_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_257_ _005_ _007_ _014_ vssd1 vssd1 vccd1 vccd1 _015_ sky130_fd_sc_hd__a21oi_1
X_326_ _067_ _068_ _070_ _071_ vssd1 vssd1 vccd1 vccd1 _075_ sky130_fd_sc_hd__o211ai_1
Xfanout90 net51 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_1
XFILLER_18_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__488__S net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_309_ net7 net25 _057_ _055_ vssd1 vssd1 vccd1 vccd1 _058_ sky130_fd_sc_hd__a31o_2
XFILLER_6_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_90 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 pm_s3_o[1] sky130_fd_sc_hd__buf_4
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 pm_s1_o[6] sky130_fd_sc_hd__buf_4
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 pm_s0_o[3] sky130_fd_sc_hd__buf_4
XANTENNA_input16_A bm_s3_s3_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input8_A bm_s1_s2_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_290_ _041_ _043_ _044_ _040_ _013_ vssd1 vssd1 vccd1 vccd1 _046_ sky130_fd_sc_hd__o221a_1
XFILLER_13_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_488_ _203_ _207_ net86 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__mux2_1
XFILLER_3_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout109 net20 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_3_70 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_411_ _140_ _142_ vssd1 vssd1 vccd1 vccd1 _151_ sky130_fd_sc_hd__and2_1
X_273_ _028_ _029_ _030_ vssd1 vssd1 vccd1 vccd1 _031_ sky130_fd_sc_hd__a21o_1
X_342_ net23 net22 _076_ vssd1 vssd1 vccd1 vccd1 _091_ sky130_fd_sc_hd__and3_1
XFILLER_12_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout91 _045_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_2
X_256_ _008_ _012_ _013_ _011_ vssd1 vssd1 vccd1 vccd1 _014_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_0_60 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_325_ _059_ _065_ vssd1 vssd1 vccd1 vccd1 _074_ sky130_fd_sc_hd__nor2_1
XFILLER_9_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input46_A pm_s3_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_239_ net12 net34 vssd1 vssd1 vccd1 vccd1 _224_ sky130_fd_sc_hd__and2_1
X_308_ net8 net26 vssd1 vssd1 vccd1 vccd1 _057_ sky130_fd_sc_hd__xor2_1
XFILLER_20_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_91 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 pm_s0_o[4] sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 pm_s3_o[2] sky130_fd_sc_hd__buf_4
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 pm_s1_o[7] sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_15_Left_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_487_ _197_ _196_ net85 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__mux2_1
XFILLER_8_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_410_ _148_ _149_ vssd1 vssd1 vccd1 vccd1 _150_ sky130_fd_sc_hd__nor2_1
X_272_ net94 _022_ _018_ _019_ vssd1 vssd1 vccd1 vccd1 _030_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_0_Left_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_341_ _086_ _087_ vssd1 vssd1 vccd1 vccd1 _090_ sky130_fd_sc_hd__or2_1
XFILLER_5_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout92 _130_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_2
X_255_ _225_ _226_ vssd1 vssd1 vccd1 vccd1 _013_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_324_ _070_ _071_ _067_ _068_ vssd1 vssd1 vccd1 vccd1 _073_ sky130_fd_sc_hd__a211oi_1
XFILLER_9_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_61 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__304__A1 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input39_A pm_s2_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Left_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_238_ _221_ _222_ vssd1 vssd1 vccd1 vccd1 _223_ sky130_fd_sc_hd__and2_1
X_307_ net7 net25 vssd1 vssd1 vccd1 vccd1 _056_ sky130_fd_sc_hd__nand2_1
XFILLER_1_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 pm_s2_o[0] sky130_fd_sc_hd__buf_4
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 pm_s0_o[5] sky130_fd_sc_hd__buf_4
XFILLER_7_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input21_A pm_s0_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_486_ _189_ _192_ net85 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__mux2_1
XFILLER_8_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_271_ net95 _018_ vssd1 vssd1 vccd1 vccd1 _029_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_340_ _086_ _087_ _088_ vssd1 vssd1 vccd1 vccd1 _089_ sky130_fd_sc_hd__a21o_1
X_469_ _195_ _197_ vssd1 vssd1 vccd1 vccd1 _200_ sky130_fd_sc_hd__or2_1
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_254_ _009_ _010_ _226_ vssd1 vssd1 vccd1 vccd1 _012_ sky130_fd_sc_hd__and3b_1
Xfanout93 _080_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_2
X_323_ _070_ _071_ vssd1 vssd1 vccd1 vccd1 _072_ sky130_fd_sc_hd__and2_1
XFILLER_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_237_ net99 _220_ net96 vssd1 vssd1 vccd1 vccd1 _222_ sky130_fd_sc_hd__a21o_1
X_306_ net8 net26 vssd1 vssd1 vccd1 vccd1 _055_ sky130_fd_sc_hd__and2_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 pm_s0_o[6] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_17_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input14_A bm_s3_s1_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_485_ _179_ _182_ net85 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__mux2_1
XFILLER_8_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input6_A bm_s1_s0_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input17_X net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_270_ net38 _021_ vssd1 vssd1 vccd1 vccd1 _028_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_399_ _121_ _128_ _129_ _137_ _138_ vssd1 vssd1 vccd1 vccd1 _139_ sky130_fd_sc_hd__a311o_1
X_468_ _195_ _197_ _198_ vssd1 vssd1 vccd1 vccd1 _199_ sky130_fd_sc_hd__a21o_1
XFILLER_4_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_322_ net107 _058_ net106 vssd1 vssd1 vccd1 vccd1 _071_ sky130_fd_sc_hd__a21o_1
Xfanout94 _021_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_2
X_253_ _009_ _010_ vssd1 vssd1 vccd1 vccd1 _011_ sky130_fd_sc_hd__and2b_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_236_ net96 net99 _220_ vssd1 vssd1 vccd1 vccd1 _221_ sky130_fd_sc_hd__nand3_1
X_305_ _214_ _053_ vssd1 vssd1 vccd1 vccd1 _054_ sky130_fd_sc_hd__xnor2_1
XFILLER_1_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input44_A pm_s3_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput49 net86 vssd1 vssd1 vccd1 vccd1 dec_bits_o[0] sky130_fd_sc_hd__buf_4
XFILLER_22_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_484_ _162_ _167_ net85 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__mux2_1
XFILLER_8_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_398_ _125_ _126_ _122_ _123_ vssd1 vssd1 vccd1 vccd1 _138_ sky130_fd_sc_hd__o211a_1
XFILLER_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_467_ _190_ _191_ _187_ _188_ vssd1 vssd1 vccd1 vccd1 _198_ sky130_fd_sc_hd__o211a_1
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout95 net46 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_2
X_252_ net11 net33 vssd1 vssd1 vccd1 vccd1 _010_ sky130_fd_sc_hd__xor2_1
XFILLER_13_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_321_ net107 net106 _058_ vssd1 vssd1 vccd1 vccd1 _070_ sky130_fd_sc_hd__nand3_1
X_235_ _218_ _219_ _217_ vssd1 vssd1 vccd1 vccd1 _220_ sky130_fd_sc_hd__o21ai_4
X_304_ net17 net3 _052_ _051_ vssd1 vssd1 vccd1 vccd1 _053_ sky130_fd_sc_hd__a31o_1
XFILLER_1_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_7_Left_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input37_A pm_s2_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_483_ _171_ _169_ net85 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__mux2_1
X_397_ net92 _131_ _134_ _135_ vssd1 vssd1 vccd1 vccd1 _137_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_20_Left_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_466_ net22 _187_ vssd1 vssd1 vccd1 vccd1 _197_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_251_ net15 net41 vssd1 vssd1 vccd1 vccd1 _009_ sky130_fd_sc_hd__xor2_1
Xfanout96 net44 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_2
Xfanout85 net86 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_320_ _067_ _068_ vssd1 vssd1 vccd1 vccd1 _069_ sky130_fd_sc_hd__nor2_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_449_ net107 net106 _166_ vssd1 vssd1 vccd1 vccd1 _180_ sky130_fd_sc_hd__and3_1
X_234_ net16 net42 vssd1 vssd1 vccd1 vccd1 _219_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_23_Left_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_303_ net18 net4 vssd1 vssd1 vccd1 vccd1 _052_ sky130_fd_sc_hd__xor2_2
XFILLER_19_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_482_ _158_ _173_ net85 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__mux2_1
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_396_ _134_ _135_ vssd1 vssd1 vccd1 vccd1 _136_ sky130_fd_sc_hd__and2_1
XANTENNA_input12_A bm_s2_s3_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_465_ _195_ vssd1 vssd1 vccd1 vccd1 _196_ sky130_fd_sc_hd__inv_2
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout97 net44 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__buf_1
X_250_ _218_ _219_ vssd1 vssd1 vccd1 vccd1 _008_ sky130_fd_sc_hd__xnor2_1
Xfanout86 net49 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input4_A bm_s0_s2_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_379_ _117_ _118_ vssd1 vssd1 vccd1 vccd1 _119_ sky130_fd_sc_hd__and2b_1
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_448_ _177_ _178_ vssd1 vssd1 vccd1 vccd1 _179_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_9_86 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_233_ net15 net41 vssd1 vssd1 vccd1 vccd1 _218_ sky130_fd_sc_hd__nand2_1
X_302_ net18 net4 vssd1 vssd1 vccd1 vccd1 _051_ sky130_fd_sc_hd__and2_1
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input42_A pm_s3_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_481_ _209_ _210_ _211_ _208_ vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__o22a_1
XFILLER_12_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_464_ net105 _190_ vssd1 vssd1 vccd1 vccd1 _195_ sky130_fd_sc_hd__xnor2_1
X_395_ net102 net104 _111_ net37 vssd1 vssd1 vccd1 vccd1 _135_ sky130_fd_sc_hd__a31o_1
XFILLER_4_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout87 net88 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_2
Xfanout98 net43 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_378_ net33 net9 vssd1 vssd1 vccd1 vccd1 _118_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_0_56 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_447_ net110 _161_ net109 vssd1 vssd1 vccd1 vccd1 _178_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_9_87 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_232_ net16 net42 vssd1 vssd1 vccd1 vccd1 _217_ sky130_fd_sc_hd__nand2_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_301_ net111 net3 vssd1 vssd1 vccd1 vccd1 _050_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_77 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input35_A pm_s2_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_480_ _203_ _206_ _209_ _210_ vssd1 vssd1 vccd1 vccd1 _211_ sky130_fd_sc_hd__a22o_1
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout85_A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_394_ net37 net102 net104 _111_ vssd1 vssd1 vccd1 vccd1 _134_ sky130_fd_sc_hd__nand4_2
X_463_ _176_ _183_ _184_ _185_ _193_ vssd1 vssd1 vccd1 vccd1 _194_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_13_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout99 net43 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_2
Xfanout88 net50 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dlymetal6s2s_1
X_377_ net41 net13 vssd1 vssd1 vccd1 vccd1 _117_ sky130_fd_sc_hd__xor2_1
XFILLER_1_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_57 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_446_ _213_ _214_ _161_ vssd1 vssd1 vccd1 vccd1 _177_ sky130_fd_sc_hd__or3b_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_88 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_300_ _047_ _048_ vssd1 vssd1 vccd1 vccd1 _049_ sky130_fd_sc_hd__and2_1
X_231_ net21 vssd1 vssd1 vccd1 vccd1 _216_ sky130_fd_sc_hd__inv_2
X_429_ net18 net2 vssd1 vssd1 vccd1 vccd1 _160_ sky130_fd_sc_hd__xor2_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput1 bm_s0_s0_i[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_27_Left_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Left_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_78 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input28_A pm_s1_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_68 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_393_ net37 net102 net104 _111_ vssd1 vssd1 vccd1 vccd1 _133_ sky130_fd_sc_hd__and4_1
XFILLER_4_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_462_ _187_ _188_ _190_ _191_ vssd1 vssd1 vccd1 vccd1 _193_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_13_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input10_A bm_s2_s1_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_58 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout89 net90 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_2
X_376_ _113_ _114_ vssd1 vssd1 vccd1 vccd1 _116_ sky130_fd_sc_hd__or2_1
X_445_ _162_ _168_ _170_ _171_ _175_ vssd1 vssd1 vccd1 vccd1 _176_ sky130_fd_sc_hd__o221a_1
XFILLER_24_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input2_A bm_s0_s0_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_230_ net107 vssd1 vssd1 vccd1 vccd1 _215_ sky130_fd_sc_hd__inv_2
X_428_ net18 net2 vssd1 vssd1 vccd1 vccd1 _159_ sky130_fd_sc_hd__and2_1
X_359_ _087_ _085_ net90 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__mux2_1
Xinput2 bm_s0_s0_i[1] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_10_89 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_79 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input40_A pm_s2_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_69 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_392_ net92 _131_ vssd1 vssd1 vccd1 vccd1 _132_ sky130_fd_sc_hd__nor2_1
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_461_ _190_ _191_ vssd1 vssd1 vccd1 vccd1 _192_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_59 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_375_ _114_ vssd1 vssd1 vccd1 vccd1 _115_ sky130_fd_sc_hd__inv_2
X_444_ _170_ _171_ _174_ _158_ vssd1 vssd1 vccd1 vccd1 _175_ sky130_fd_sc_hd__a22o_1
X_358_ _079_ _082_ net89 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__mux2_1
X_427_ _156_ _157_ vssd1 vssd1 vccd1 vccd1 _158_ sky130_fd_sc_hd__and2_1
XFILLER_1_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_289_ _009_ _010_ net91 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__mux2_1
Xinput3 bm_s0_s2_i[0] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_1
XFILLER_19_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input33_A pm_s2_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_391_ net96 net98 _105_ net45 vssd1 vssd1 vccd1 vccd1 _131_ sky130_fd_sc_hd__a31oi_2
X_460_ net108 net106 _166_ net29 vssd1 vssd1 vccd1 vccd1 _191_ sky130_fd_sc_hd__a31oi_2
XFILLER_4_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_374_ _103_ _104_ vssd1 vssd1 vccd1 vccd1 _114_ sky130_fd_sc_hd__xnor2_1
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_443_ _164_ _172_ vssd1 vssd1 vccd1 vccd1 _174_ sky130_fd_sc_hd__nand2_1
XFILLER_24_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout86_X net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_288_ _045_ vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__inv_2
X_426_ net111 net1 vssd1 vssd1 vccd1 vccd1 _157_ sky130_fd_sc_hd__or2_1
X_357_ _069_ _072_ net89 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__mux2_1
Xinput4 bm_s0_s2_i[1] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_1
XFILLER_19_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_409_ net100 _133_ net39 vssd1 vssd1 vccd1 vccd1 _149_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput40 pm_s2_i[7] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_7_80 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input26_A pm_s1_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_390_ net45 net96 net98 _105_ vssd1 vssd1 vccd1 vccd1 _130_ sky130_fd_sc_hd__and4_1
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_373_ _109_ _110_ vssd1 vssd1 vccd1 vccd1 _113_ sky130_fd_sc_hd__xnor2_1
X_442_ _164_ _172_ vssd1 vssd1 vccd1 vccd1 _173_ sky130_fd_sc_hd__and2_1
XFILLER_24_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_287_ _041_ _043_ _044_ _040_ vssd1 vssd1 vccd1 vccd1 _045_ sky130_fd_sc_hd__o22a_1
XFILLER_14_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_356_ _054_ _059_ net89 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__mux2_1
X_425_ net111 net1 vssd1 vssd1 vccd1 vccd1 _156_ sky130_fd_sc_hd__nand2_1
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput5 bm_s1_s0_i[0] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_408_ net39 net100 _133_ vssd1 vssd1 vccd1 vccd1 _148_ sky130_fd_sc_hd__and3_1
X_339_ net93 _081_ _077_ _078_ vssd1 vssd1 vccd1 vccd1 _088_ sky130_fd_sc_hd__o211a_1
XFILLER_21_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput41 pm_s3_i[0] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_2
Xinput30 pm_s1_i[5] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_81 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input19_A pm_s0_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_71 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_372_ _212_ _111_ vssd1 vssd1 vccd1 vccd1 _112_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_441_ net25 net5 vssd1 vssd1 vccd1 vccd1 _172_ sky130_fd_sc_hd__or2_1
XFILLER_5_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_424_ _153_ _154_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__and2b_1
X_286_ _034_ _037_ _041_ _043_ vssd1 vssd1 vccd1 vccd1 _044_ sky130_fd_sc_hd__a22o_1
X_355_ _064_ _060_ net89 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__mux2_1
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 bm_s1_s0_i[1] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_407_ _146_ vssd1 vssd1 vccd1 vccd1 _147_ sky130_fd_sc_hd__inv_2
XFILLER_24_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Left_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_269_ net100 net94 vssd1 vssd1 vccd1 vccd1 _027_ sky130_fd_sc_hd__xor2_1
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_338_ net22 _077_ vssd1 vssd1 vccd1 vccd1 _087_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_92 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput31 pm_s1_i[6] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_1
Xinput20 pm_s0_i[3] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_1
XFILLER_23_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_82 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput42 pm_s3_i[1] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_2
XFILLER_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input31_A pm_s1_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_72 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_371_ net33 net9 _109_ _108_ vssd1 vssd1 vccd1 vccd1 _111_ sky130_fd_sc_hd__a31o_2
X_440_ _156_ _160_ vssd1 vssd1 vccd1 vccd1 _171_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_423_ _150_ _147_ net88 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__mux2_1
X_285_ net40 _035_ vssd1 vssd1 vccd1 vccd1 _043_ sky130_fd_sc_hd__xnor2_2
X_354_ _049_ _061_ net89 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_62 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 bm_s1_s2_i[0] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_406_ _144_ _145_ vssd1 vssd1 vccd1 vccd1 _146_ sky130_fd_sc_hd__or2_1
X_268_ _004_ _015_ _016_ _024_ _025_ vssd1 vssd1 vccd1 vccd1 _026_ sky130_fd_sc_hd__o311a_1
X_337_ net105 net93 vssd1 vssd1 vccd1 vccd1 _086_ sky130_fd_sc_hd__xnor2_1
XFILLER_2_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_93 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput43 pm_s3_i[2] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_1
Xinput32 pm_s1_i[7] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_1
Xinput21 pm_s0_i[4] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_22_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput10 bm_s2_s1_i[1] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input24_A pm_s0_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_73 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_370_ net33 net9 vssd1 vssd1 vccd1 vccd1 _110_ sky130_fd_sc_hd__nand2_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_422_ _140_ _141_ net87 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__mux2_1
X_284_ _041_ vssd1 vssd1 vccd1 vccd1 _042_ sky130_fd_sc_hd__inv_2
X_353_ _099_ _100_ _101_ _098_ vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__o22a_1
Xinput8 bm_s1_s2_i[1] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_1_63 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_405_ net95 _130_ net47 vssd1 vssd1 vccd1 vccd1 _145_ sky130_fd_sc_hd__a21oi_1
XFILLER_25_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_267_ _221_ _222_ _001_ _002_ vssd1 vssd1 vccd1 vccd1 _025_ sky130_fd_sc_hd__a211o_1
X_336_ net105 net93 vssd1 vssd1 vccd1 vccd1 _085_ sky130_fd_sc_hd__xor2_1
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput44 pm_s3_i[3] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
Xinput33 pm_s2_i[0] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_2
Xinput22 pm_s0_i[5] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_2
Xinput11 bm_s2_s3_i[0] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_1
X_319_ net110 _053_ net109 vssd1 vssd1 vccd1 vccd1 _068_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_22_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input17_A pm_s0_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input9_A bm_s2_s1_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_421_ _136_ _132_ net87 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__mux2_1
X_283_ net48 _032_ vssd1 vssd1 vccd1 vccd1 _041_ sky130_fd_sc_hd__xor2_2
Xinput9 bm_s2_s1_i[0] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_64 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_352_ _093_ _096_ _099_ _100_ vssd1 vssd1 vccd1 vccd1 _101_ sky130_fd_sc_hd__a22o_1
XFILLER_27_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_404_ net47 net46 net92 vssd1 vssd1 vccd1 vccd1 _144_ sky130_fd_sc_hd__and3_1
X_266_ _018_ _019_ net94 _022_ vssd1 vssd1 vccd1 vccd1 _024_ sky130_fd_sc_hd__a211o_1
X_335_ _066_ _073_ _074_ _075_ _083_ vssd1 vssd1 vccd1 vccd1 _084_ sky130_fd_sc_hd__o311a_1
XFILLER_24_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input47_A pm_s3_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_73 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput45 pm_s3_i[4] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_2
Xinput34 pm_s2_i[1] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput23 pm_s0_i[6] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_26_Left_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput12 bm_s2_s3_i[1] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_1
X_249_ _212_ _000_ vssd1 vssd1 vccd1 vccd1 _007_ sky130_fd_sc_hd__xnor2_1
X_318_ net109 net110 _053_ vssd1 vssd1 vccd1 vccd1 _067_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_10_Left_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_282_ _026_ _031_ _034_ _037_ _039_ vssd1 vssd1 vccd1 vccd1 _040_ sky130_fd_sc_hd__o221a_1
X_420_ _124_ _127_ net87 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__mux2_1
X_351_ net24 _091_ vssd1 vssd1 vccd1 vccd1 _100_ sky130_fd_sc_hd__xor2_1
X_403_ net92 _131_ _136_ _140_ _142_ vssd1 vssd1 vccd1 vccd1 _143_ sky130_fd_sc_hd__o32a_1
XFILLER_18_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_334_ _077_ _078_ net93 _081_ vssd1 vssd1 vccd1 vccd1 _083_ sky130_fd_sc_hd__a211o_1
X_265_ net94 _022_ vssd1 vssd1 vccd1 vccd1 _023_ sky130_fd_sc_hd__nor2_1
XFILLER_2_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput46 pm_s3_i[5] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
Xinput35 pm_s2_i[2] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
Xinput24 pm_s0_i[7] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_1
Xinput13 bm_s3_s1_i[0] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_1
X_248_ _005_ vssd1 vssd1 vccd1 vccd1 _006_ sky130_fd_sc_hd__inv_2
XFILLER_14_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_317_ _059_ _065_ _054_ vssd1 vssd1 vccd1 vccd1 _066_ sky130_fd_sc_hd__a21boi_1
XFILLER_14_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input22_A pm_s0_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_281_ _028_ _029_ vssd1 vssd1 vccd1 vccd1 _039_ sky130_fd_sc_hd__or2_1
XFILLER_14_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_350_ net32 _094_ vssd1 vssd1 vccd1 vccd1 _099_ sky130_fd_sc_hd__xnor2_1
X_479_ net24 _201_ vssd1 vssd1 vccd1 vccd1 _210_ sky130_fd_sc_hd__xor2_1
X_402_ net95 net92 vssd1 vssd1 vccd1 vccd1 _142_ sky130_fd_sc_hd__xnor2_1
X_264_ net101 net104 _000_ net37 vssd1 vssd1 vccd1 vccd1 _022_ sky130_fd_sc_hd__a31oi_2
XFILLER_2_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_333_ net93 _081_ vssd1 vssd1 vccd1 vccd1 _082_ sky130_fd_sc_hd__nor2_1
XFILLER_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput36 pm_s2_i[3] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
Xinput25 pm_s1_i[0] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_2
Xinput14 bm_s3_s1_i[1] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_1
X_247_ net99 _220_ vssd1 vssd1 vccd1 vccd1 _005_ sky130_fd_sc_hd__xnor2_1
X_316_ _062_ _064_ _063_ _060_ vssd1 vssd1 vccd1 vccd1 _065_ sky130_fd_sc_hd__a2bb2o_1
Xinput47 pm_s3_i[6] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__buf_1
XFILLER_11_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input15_A bm_s3_s3_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_280_ _037_ vssd1 vssd1 vccd1 vccd1 _038_ sky130_fd_sc_hd__inv_2
XFILLER_14_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input7_A bm_s1_s2_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_478_ net32 _204_ vssd1 vssd1 vccd1 vccd1 _209_ sky130_fd_sc_hd__xnor2_1
X_401_ net95 net92 vssd1 vssd1 vccd1 vccd1 _141_ sky130_fd_sc_hd__xor2_1
XFILLER_25_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_263_ net37 net101 net103 _000_ vssd1 vssd1 vccd1 vccd1 _021_ sky130_fd_sc_hd__and4_1
XFILLER_18_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_332_ net108 net28 _058_ net29 vssd1 vssd1 vccd1 vccd1 _081_ sky130_fd_sc_hd__a31oi_2
XFILLER_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput48 pm_s3_i[7] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput37 pm_s2_i[4] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput26 pm_s1_i[1] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_2
Xinput15 bm_s3_s3_i[0] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_1
X_246_ _001_ _002_ _221_ _222_ vssd1 vssd1 vccd1 vccd1 _004_ sky130_fd_sc_hd__o211a_1
X_315_ _047_ _052_ vssd1 vssd1 vccd1 vccd1 _064_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input45_A pm_s3_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_229_ net110 vssd1 vssd1 vccd1 vccd1 _214_ sky130_fd_sc_hd__inv_2
XFILLER_8_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_477_ _194_ _199_ _203_ _206_ _200_ vssd1 vssd1 vccd1 vccd1 _208_ sky130_fd_sc_hd__o221a_1
X_400_ net100 _134_ vssd1 vssd1 vccd1 vccd1 _140_ sky130_fd_sc_hd__xnor2_1
X_262_ _018_ _019_ vssd1 vssd1 vccd1 vccd1 _020_ sky130_fd_sc_hd__and2_1
X_331_ net108 net28 net29 _058_ vssd1 vssd1 vccd1 vccd1 _080_ sky130_fd_sc_hd__and4_1
XFILLER_23_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput38 pm_s2_i[5] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_1
Xinput27 pm_s1_i[2] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_1
Xinput16 bm_s3_s3_i[1] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_1
X_245_ _001_ _002_ vssd1 vssd1 vccd1 vccd1 _003_ sky130_fd_sc_hd__nor2_1
XFILLER_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_314_ _050_ _061_ _052_ vssd1 vssd1 vccd1 vccd1 _063_ sky130_fd_sc_hd__or3b_1
XFILLER_20_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input38_A pm_s2_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_228_ net109 vssd1 vssd1 vccd1 vccd1 _213_ sky130_fd_sc_hd__inv_2
XFILLER_3_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input20_A pm_s0_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_476_ _206_ vssd1 vssd1 vccd1 vccd1 _207_ sky130_fd_sc_hd__inv_2
XFILLER_14_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_261_ net97 net99 _220_ net45 vssd1 vssd1 vccd1 vccd1 _019_ sky130_fd_sc_hd__a31o_1
X_330_ _077_ _078_ vssd1 vssd1 vccd1 vccd1 _079_ sky130_fd_sc_hd__and2_1
X_459_ net108 net106 net29 _166_ vssd1 vssd1 vccd1 vccd1 _190_ sky130_fd_sc_hd__and4_2
XFILLER_23_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput39 pm_s2_i[6] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_1
Xinput28 pm_s1_i[3] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_1
Xinput17 pm_s0_i[0] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
X_244_ net103 _000_ net101 vssd1 vssd1 vccd1 vccd1 _002_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_16_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_313_ _050_ _061_ vssd1 vssd1 vccd1 vccd1 _062_ sky130_fd_sc_hd__nor2_1
X_227_ net103 vssd1 vssd1 vccd1 vccd1 _212_ sky130_fd_sc_hd__inv_2
XFILLER_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input13_A bm_s3_s1_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_475_ _204_ _205_ vssd1 vssd1 vccd1 vccd1 _206_ sky130_fd_sc_hd__or2_1
XFILLER_25_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_260_ net45 net97 net99 _220_ vssd1 vssd1 vccd1 vccd1 _018_ sky130_fd_sc_hd__nand4_2
XANTENNA_input5_A bm_s1_s0_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_389_ _107_ _112_ vssd1 vssd1 vccd1 vccd1 _129_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_19_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_458_ _187_ _188_ vssd1 vssd1 vccd1 vccd1 _189_ sky130_fd_sc_hd__and2_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput29 pm_s1_i[4] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_2
Xinput18 pm_s0_i[1] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_2
X_243_ net101 net103 _000_ vssd1 vssd1 vccd1 vccd1 _001_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_16_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_312_ net7 net25 vssd1 vssd1 vccd1 vccd1 _061_ sky130_fd_sc_hd__xor2_2
XFILLER_22_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input43_A pm_s3_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_474_ net105 _190_ net31 vssd1 vssd1 vccd1 vccd1 _205_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_19_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_388_ _122_ _123_ _125_ _126_ vssd1 vssd1 vccd1 vccd1 _128_ sky130_fd_sc_hd__a211o_1
X_457_ net109 net110 _161_ net21 vssd1 vssd1 vccd1 vccd1 _188_ sky130_fd_sc_hd__a31o_1
Xinput19 pm_s0_i[2] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_24_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_242_ net11 net33 _226_ _224_ vssd1 vssd1 vccd1 vccd1 _000_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_16_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_311_ _056_ _057_ vssd1 vssd1 vccd1 vccd1 _060_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input36_A pm_s2_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_9_Left_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_473_ net31 net105 _190_ vssd1 vssd1 vccd1 vccd1 _204_ sky130_fd_sc_hd__and3_1
XFILLER_25_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_387_ _125_ _126_ vssd1 vssd1 vccd1 vccd1 _127_ sky130_fd_sc_hd__nor2_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_456_ _213_ _214_ _216_ _161_ vssd1 vssd1 vccd1 vccd1 _187_ sky130_fd_sc_hd__or4b_2
XTAP_TAPCELL_ROW_24_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_310_ _215_ _058_ vssd1 vssd1 vccd1 vccd1 _059_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_241_ net12 net34 vssd1 vssd1 vccd1 vccd1 _226_ sky130_fd_sc_hd__xor2_1
X_439_ _164_ _165_ vssd1 vssd1 vccd1 vccd1 _170_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_21_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input29_A pm_s1_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_12_Left_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_472_ _201_ _202_ vssd1 vssd1 vccd1 vccd1 _203_ sky130_fd_sc_hd__nor2_1
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_386_ net98 _105_ net96 vssd1 vssd1 vccd1 vccd1 _126_ sky130_fd_sc_hd__a21oi_1
XANTENNA_input11_A bm_s2_s3_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_455_ net109 net110 net21 _161_ vssd1 vssd1 vccd1 vccd1 _186_ sky130_fd_sc_hd__and4_1
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input3_A bm_s0_s2_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_240_ net11 net33 vssd1 vssd1 vccd1 vccd1 _225_ sky130_fd_sc_hd__nand2_1
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_369_ net34 net10 vssd1 vssd1 vccd1 vccd1 _109_ sky130_fd_sc_hd__xor2_1
XFILLER_13_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_438_ _164_ _165_ vssd1 vssd1 vccd1 vccd1 _169_ sky130_fd_sc_hd__xor2_1
XFILLER_9_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout110 net19 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout111_A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input41_A pm_s3_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_471_ net22 _186_ net23 vssd1 vssd1 vccd1 vccd1 _202_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_27_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_385_ net96 net98 _105_ vssd1 vssd1 vccd1 vccd1 _125_ sky130_fd_sc_hd__and3_1
XFILLER_17_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_454_ _177_ _178_ _180_ _181_ vssd1 vssd1 vccd1 vccd1 _185_ sky130_fd_sc_hd__a211o_1
XFILLER_11_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 pm_s3_o[3] sky130_fd_sc_hd__buf_4
XFILLER_20_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_368_ net34 net10 vssd1 vssd1 vccd1 vccd1 _108_ sky130_fd_sc_hd__and2_1
X_299_ net111 net3 vssd1 vssd1 vccd1 vccd1 _048_ sky130_fd_sc_hd__or2_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_437_ net107 _166_ vssd1 vssd1 vccd1 vccd1 _168_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout100 net38 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout111 net17 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_83 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input34_A pm_s2_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_470_ net23 net22 _186_ vssd1 vssd1 vccd1 vccd1 _201_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_27_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_384_ _122_ _123_ vssd1 vssd1 vccd1 vccd1 _124_ sky130_fd_sc_hd__and2_1
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_453_ _162_ _168_ vssd1 vssd1 vccd1 vccd1 _184_ sky130_fd_sc_hd__and2_1
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 pm_s3_o[4] sky130_fd_sc_hd__buf_4
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 pm_s2_o[1] sky130_fd_sc_hd__buf_4
X_367_ net98 _105_ vssd1 vssd1 vccd1 vccd1 _107_ sky130_fd_sc_hd__xnor2_1
X_298_ net111 net3 vssd1 vssd1 vccd1 vccd1 _047_ sky130_fd_sc_hd__nand2_1
X_436_ _215_ _166_ vssd1 vssd1 vccd1 vccd1 _167_ sky130_fd_sc_hd__xnor2_1
Xfanout101 net36 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_419_ _112_ _106_ net87 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_84 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input27_A pm_s1_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_74 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Left_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_383_ net103 _111_ net101 vssd1 vssd1 vccd1 vccd1 _123_ sky130_fd_sc_hd__a21o_1
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_452_ _180_ _181_ _177_ _178_ vssd1 vssd1 vccd1 vccd1 _183_ sky130_fd_sc_hd__o211a_1
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 pm_s3_o[5] sky130_fd_sc_hd__buf_4
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 pm_s2_o[2] sky130_fd_sc_hd__buf_4
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 pm_s0_o[7] sky130_fd_sc_hd__buf_4
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_366_ net98 _105_ vssd1 vssd1 vccd1 vccd1 _106_ sky130_fd_sc_hd__xor2_1
X_297_ _042_ _043_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__nor2_1
X_435_ _164_ _165_ _163_ vssd1 vssd1 vccd1 vccd1 _166_ sky130_fd_sc_hd__o21ai_4
XFILLER_9_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout102 net36 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__buf_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input1_A bm_s0_s0_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_418_ _113_ _115_ net87 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__mux2_1
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_349_ _084_ _089_ _093_ _096_ _090_ vssd1 vssd1 vccd1 vccd1 _098_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_8_85 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_75 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_382_ net101 net103 _111_ vssd1 vssd1 vccd1 vccd1 _122_ sky130_fd_sc_hd__nand3_1
XFILLER_15_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput50 net88 vssd1 vssd1 vccd1 vccd1 dec_bits_o[1] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_2_65 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 pm_s3_o[6] sky130_fd_sc_hd__buf_4
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 pm_s2_o[3] sky130_fd_sc_hd__buf_4
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 pm_s1_o[0] sky130_fd_sc_hd__buf_4
X_451_ _180_ _181_ vssd1 vssd1 vccd1 vccd1 _182_ sky130_fd_sc_hd__nor2_1
X_365_ _103_ _104_ _102_ vssd1 vssd1 vccd1 vccd1 _105_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_15_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_296_ _034_ _038_ net91 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__mux2_1
X_434_ net26 net6 vssd1 vssd1 vccd1 vccd1 _165_ sky130_fd_sc_hd__xnor2_2
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_76 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout103 net35 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_12_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_279_ _035_ _036_ vssd1 vssd1 vccd1 vccd1 _037_ sky130_fd_sc_hd__or2_1
X_417_ _118_ _117_ net87 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_348_ _096_ vssd1 vssd1 vccd1 vccd1 _097_ sky130_fd_sc_hd__inv_2
XFILLER_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_76 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input32_A pm_s1_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_381_ _107_ _112_ _116_ _120_ vssd1 vssd1 vccd1 vccd1 _121_ sky130_fd_sc_hd__a22o_1
Xoutput51 net90 vssd1 vssd1 vccd1 vccd1 dec_bits_o[2] sky130_fd_sc_hd__buf_4
XFILLER_15_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_66 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 pm_s2_o[4] sky130_fd_sc_hd__buf_4
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 pm_s1_o[1] sky130_fd_sc_hd__buf_4
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 pm_s3_o[7] sky130_fd_sc_hd__buf_4
X_450_ net107 _166_ net106 vssd1 vssd1 vccd1 vccd1 _181_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_18_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_433_ net25 net5 vssd1 vssd1 vccd1 vccd1 _164_ sky130_fd_sc_hd__nand2_2
X_364_ net41 net13 vssd1 vssd1 vccd1 vccd1 _104_ sky130_fd_sc_hd__nand2_1
X_295_ _029_ _027_ net91 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__mux2_1
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout104 net35 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_12_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_416_ _153_ _154_ _155_ _152_ vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__a22o_1
X_278_ net100 net94 net39 vssd1 vssd1 vccd1 vccd1 _036_ sky130_fd_sc_hd__a21oi_1
X_347_ _094_ _095_ vssd1 vssd1 vccd1 vccd1 _096_ sky130_fd_sc_hd__or2_1
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input25_A pm_s1_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 dec_bits_o[3] sky130_fd_sc_hd__buf_4
X_380_ _113_ _114_ _119_ vssd1 vssd1 vccd1 vccd1 _120_ sky130_fd_sc_hd__a21o_1
XFILLER_15_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_67 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 pm_s2_o[5] sky130_fd_sc_hd__buf_4
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 pm_s1_o[2] sky130_fd_sc_hd__buf_4
.ends

