magic
tech sky130A
magscale 1 2
timestamp 1769196442
<< viali >>
rect 1501 25177 1535 25211
rect 1777 25177 1811 25211
rect 1593 25109 1627 25143
rect 1501 24769 1535 24803
rect 1777 24769 1811 24803
rect 1593 24565 1627 24599
rect 1409 24157 1443 24191
rect 1685 24157 1719 24191
rect 6837 24157 6871 24191
rect 7205 24157 7239 24191
rect 7021 24089 7055 24123
rect 7113 24089 7147 24123
rect 1593 24021 1627 24055
rect 7389 24021 7423 24055
rect 7297 23817 7331 23851
rect 7481 23817 7515 23851
rect 8033 23817 8067 23851
rect 1501 23681 1535 23715
rect 1961 23681 1995 23715
rect 2881 23681 2915 23715
rect 2973 23681 3007 23715
rect 3249 23681 3283 23715
rect 3525 23681 3559 23715
rect 4445 23681 4479 23715
rect 6561 23681 6595 23715
rect 7300 23681 7334 23715
rect 7849 23681 7883 23715
rect 7941 23681 7975 23715
rect 8401 23681 8435 23715
rect 8585 23681 8619 23715
rect 6837 23613 6871 23647
rect 7665 23613 7699 23647
rect 8309 23613 8343 23647
rect 1777 23545 1811 23579
rect 3157 23545 3191 23579
rect 4353 23545 4387 23579
rect 6929 23545 6963 23579
rect 8217 23545 8251 23579
rect 1593 23477 1627 23511
rect 2697 23477 2731 23511
rect 3433 23477 3467 23511
rect 6653 23477 6687 23511
rect 8769 23477 8803 23511
rect 7389 23273 7423 23307
rect 8033 23273 8067 23307
rect 2973 23205 3007 23239
rect 7573 23205 7607 23239
rect 8125 23205 8159 23239
rect 8217 23205 8251 23239
rect 4629 23137 4663 23171
rect 6929 23137 6963 23171
rect 1409 23069 1443 23103
rect 1685 23069 1719 23103
rect 2421 23069 2455 23103
rect 2605 23069 2639 23103
rect 2789 23069 2823 23103
rect 3065 23069 3099 23103
rect 3341 23069 3375 23103
rect 3433 23069 3467 23103
rect 3801 23069 3835 23103
rect 3985 23069 4019 23103
rect 4077 23069 4111 23103
rect 4261 23069 4295 23103
rect 4721 23069 4755 23103
rect 6837 23069 6871 23103
rect 7113 23069 7147 23103
rect 7205 23069 7239 23103
rect 7481 23069 7515 23103
rect 7757 23069 7791 23103
rect 7849 23069 7883 23103
rect 2697 23001 2731 23035
rect 3249 23001 3283 23035
rect 3893 23001 3927 23035
rect 8585 23001 8619 23035
rect 3617 22933 3651 22967
rect 4169 22933 4203 22967
rect 3617 22729 3651 22763
rect 7757 22729 7791 22763
rect 1501 22593 1535 22627
rect 1777 22593 1811 22627
rect 2145 22593 2179 22627
rect 2237 22593 2271 22627
rect 2513 22593 2547 22627
rect 3709 22593 3743 22627
rect 7665 22593 7699 22627
rect 7941 22593 7975 22627
rect 28089 22593 28123 22627
rect 2605 22525 2639 22559
rect 2881 22525 2915 22559
rect 28365 22525 28399 22559
rect 1961 22457 1995 22491
rect 7941 22457 7975 22491
rect 1593 22389 1627 22423
rect 2421 22389 2455 22423
rect 2513 22185 2547 22219
rect 9045 22185 9079 22219
rect 7113 22117 7147 22151
rect 8953 22049 8987 22083
rect 2651 21981 2685 22015
rect 2881 21981 2915 22015
rect 3009 21981 3043 22015
rect 3157 21981 3191 22015
rect 3985 21981 4019 22015
rect 4353 21981 4387 22015
rect 5273 21981 5307 22015
rect 5457 21981 5491 22015
rect 5549 21981 5583 22015
rect 5641 21981 5675 22015
rect 6009 21981 6043 22015
rect 6193 21981 6227 22015
rect 6401 21981 6435 22015
rect 6837 21981 6871 22015
rect 6929 21981 6963 22015
rect 7205 21981 7239 22015
rect 9416 21981 9450 22015
rect 1501 21913 1535 21947
rect 1777 21913 1811 21947
rect 2789 21913 2823 21947
rect 4077 21913 4111 21947
rect 4169 21913 4203 21947
rect 6285 21913 6319 21947
rect 1593 21845 1627 21879
rect 3801 21845 3835 21879
rect 5825 21845 5859 21879
rect 6561 21845 6595 21879
rect 6653 21845 6687 21879
rect 9413 21845 9447 21879
rect 9597 21845 9631 21879
rect 4905 21641 4939 21675
rect 5917 21573 5951 21607
rect 8493 21573 8527 21607
rect 1409 21505 1443 21539
rect 1869 21505 1903 21539
rect 2421 21505 2455 21539
rect 2697 21505 2731 21539
rect 2789 21505 2823 21539
rect 4997 21505 5031 21539
rect 6101 21505 6135 21539
rect 6193 21505 6227 21539
rect 6561 21505 6595 21539
rect 6653 21505 6687 21539
rect 7021 21505 7055 21539
rect 7481 21505 7515 21539
rect 7757 21505 7791 21539
rect 7941 21505 7975 21539
rect 7297 21437 7331 21471
rect 8033 21437 8067 21471
rect 1685 21369 1719 21403
rect 8217 21369 8251 21403
rect 1593 21301 1627 21335
rect 2513 21301 2547 21335
rect 2973 21301 3007 21335
rect 5917 21301 5951 21335
rect 6929 21301 6963 21335
rect 7205 21301 7239 21335
rect 3893 21097 3927 21131
rect 5365 21097 5399 21131
rect 7113 21097 7147 21131
rect 1685 20961 1719 20995
rect 1409 20893 1443 20927
rect 2881 20893 2915 20927
rect 2973 20893 3007 20927
rect 3157 20893 3191 20927
rect 3341 20893 3375 20927
rect 3801 20893 3835 20927
rect 4261 20893 4295 20927
rect 5457 20893 5491 20927
rect 7021 20893 7055 20927
rect 7297 20893 7331 20927
rect 7389 20893 7423 20927
rect 9413 20893 9447 20927
rect 9506 20893 9540 20927
rect 7573 20825 7607 20859
rect 4077 20757 4111 20791
rect 4169 20757 4203 20791
rect 4537 20757 4571 20791
rect 9781 20757 9815 20791
rect 3157 20553 3191 20587
rect 2789 20485 2823 20519
rect 1409 20417 1443 20451
rect 1685 20417 1719 20451
rect 2605 20417 2639 20451
rect 2881 20417 2915 20451
rect 2973 20417 3007 20451
rect 9045 20417 9079 20451
rect 9138 20417 9172 20451
rect 9505 20417 9539 20451
rect 9643 20417 9677 20451
rect 9965 20417 9999 20451
rect 10058 20417 10092 20451
rect 9413 20281 9447 20315
rect 9873 20281 9907 20315
rect 1593 20213 1627 20247
rect 10149 20213 10183 20247
rect 6469 20009 6503 20043
rect 7481 20009 7515 20043
rect 9137 20009 9171 20043
rect 20808 20009 20842 20043
rect 22385 20009 22419 20043
rect 26157 20009 26191 20043
rect 3157 19941 3191 19975
rect 23305 19941 23339 19975
rect 10425 19873 10459 19907
rect 12357 19873 12391 19907
rect 13093 19873 13127 19907
rect 18797 19873 18831 19907
rect 20545 19873 20579 19907
rect 22845 19873 22879 19907
rect 24409 19873 24443 19907
rect 1409 19805 1443 19839
rect 1685 19805 1719 19839
rect 6377 19805 6411 19839
rect 7389 19805 7423 19839
rect 9321 19805 9355 19839
rect 9505 19805 9539 19839
rect 9781 19805 9815 19839
rect 10057 19805 10091 19839
rect 10241 19805 10275 19839
rect 13277 19805 13311 19839
rect 22753 19805 22787 19839
rect 23581 19805 23615 19839
rect 2789 19737 2823 19771
rect 9413 19737 9447 19771
rect 9623 19737 9657 19771
rect 10149 19737 10183 19771
rect 12449 19737 12483 19771
rect 13369 19737 13403 19771
rect 18613 19737 18647 19771
rect 23305 19737 23339 19771
rect 24685 19737 24719 19771
rect 1593 19669 1627 19703
rect 3249 19669 3283 19703
rect 9873 19669 9907 19703
rect 12541 19669 12575 19703
rect 12909 19669 12943 19703
rect 13737 19669 13771 19703
rect 18153 19669 18187 19703
rect 18521 19669 18555 19703
rect 19073 19669 19107 19703
rect 22293 19669 22327 19703
rect 23489 19669 23523 19703
rect 1593 19465 1627 19499
rect 2329 19465 2363 19499
rect 6193 19465 6227 19499
rect 8217 19465 8251 19499
rect 8309 19465 8343 19499
rect 9689 19465 9723 19499
rect 12357 19465 12391 19499
rect 24777 19465 24811 19499
rect 18153 19397 18187 19431
rect 1409 19329 1443 19363
rect 1685 19329 1719 19363
rect 2237 19329 2271 19363
rect 2973 19329 3007 19363
rect 3893 19329 3927 19363
rect 5365 19329 5399 19363
rect 5641 19329 5675 19363
rect 5825 19329 5859 19363
rect 5917 19329 5951 19363
rect 6009 19329 6043 19363
rect 6645 19319 6679 19353
rect 6745 19329 6779 19363
rect 7021 19329 7055 19363
rect 7113 19329 7147 19363
rect 7389 19329 7423 19363
rect 7573 19329 7607 19363
rect 8033 19329 8067 19363
rect 8401 19329 8435 19363
rect 9597 19329 9631 19363
rect 9781 19329 9815 19363
rect 12725 19329 12759 19363
rect 15301 19329 15335 19363
rect 17877 19329 17911 19363
rect 22753 19329 22787 19363
rect 22937 19329 22971 19363
rect 23029 19329 23063 19363
rect 3801 19261 3835 19295
rect 6837 19261 6871 19295
rect 7941 19261 7975 19295
rect 12817 19261 12851 19295
rect 12909 19261 12943 19295
rect 22845 19261 22879 19295
rect 23305 19261 23339 19295
rect 3249 19193 3283 19227
rect 6561 19193 6595 19227
rect 3433 19125 3467 19159
rect 3525 19125 3559 19159
rect 3709 19125 3743 19159
rect 5457 19125 5491 19159
rect 7297 19125 7331 19159
rect 7481 19125 7515 19159
rect 8677 19125 8711 19159
rect 15485 19125 15519 19159
rect 19625 19125 19659 19159
rect 19809 19125 19843 19159
rect 2973 18921 3007 18955
rect 3433 18921 3467 18955
rect 4169 18921 4203 18955
rect 13185 18921 13219 18955
rect 14473 18921 14507 18955
rect 22201 18921 22235 18955
rect 23213 18921 23247 18955
rect 23397 18921 23431 18955
rect 24409 18921 24443 18955
rect 3341 18785 3375 18819
rect 4261 18785 4295 18819
rect 11253 18785 11287 18819
rect 1409 18717 1443 18751
rect 1685 18717 1719 18751
rect 2421 18717 2455 18751
rect 2789 18717 2823 18751
rect 3065 18717 3099 18751
rect 4077 18717 4111 18751
rect 4537 18717 4571 18751
rect 11437 18717 11471 18751
rect 16221 18717 16255 18751
rect 21833 18717 21867 18751
rect 24593 18717 24627 18751
rect 24685 18717 24719 18751
rect 2605 18649 2639 18683
rect 2697 18649 2731 18683
rect 11713 18649 11747 18683
rect 15945 18649 15979 18683
rect 23365 18649 23399 18683
rect 23581 18649 23615 18683
rect 1593 18581 1627 18615
rect 3617 18581 3651 18615
rect 3801 18581 3835 18615
rect 4445 18581 4479 18615
rect 22201 18581 22235 18615
rect 22385 18581 22419 18615
rect 3157 18377 3191 18411
rect 9137 18377 9171 18411
rect 12173 18377 12207 18411
rect 12541 18377 12575 18411
rect 15945 18377 15979 18411
rect 3801 18309 3835 18343
rect 4077 18309 4111 18343
rect 9781 18309 9815 18343
rect 1501 18241 1535 18275
rect 1777 18241 1811 18275
rect 3617 18241 3651 18275
rect 3893 18241 3927 18275
rect 3985 18241 4019 18275
rect 9321 18241 9355 18275
rect 9413 18241 9447 18275
rect 9689 18241 9723 18275
rect 9965 18241 9999 18275
rect 10057 18241 10091 18275
rect 14197 18241 14231 18275
rect 16221 18241 16255 18275
rect 20913 18241 20947 18275
rect 21097 18241 21131 18275
rect 23213 18241 23247 18275
rect 23305 18241 23339 18275
rect 2697 18173 2731 18207
rect 12633 18173 12667 18207
rect 12725 18173 12759 18207
rect 14473 18173 14507 18207
rect 23397 18173 23431 18207
rect 23489 18173 23523 18207
rect 3065 18105 3099 18139
rect 9781 18105 9815 18139
rect 12081 18105 12115 18139
rect 1593 18037 1627 18071
rect 3433 18037 3467 18071
rect 9597 18037 9631 18071
rect 16037 18037 16071 18071
rect 20913 18037 20947 18071
rect 23029 18037 23063 18071
rect 2329 17833 2363 17867
rect 3341 17833 3375 17867
rect 7297 17833 7331 17867
rect 14749 17833 14783 17867
rect 16313 17833 16347 17867
rect 21557 17833 21591 17867
rect 1685 17765 1719 17799
rect 2697 17697 2731 17731
rect 6837 17697 6871 17731
rect 15301 17697 15335 17731
rect 15669 17697 15703 17731
rect 18245 17697 18279 17731
rect 19809 17697 19843 17731
rect 21649 17697 21683 17731
rect 2237 17629 2271 17663
rect 3065 17629 3099 17663
rect 3157 17629 3191 17663
rect 5825 17629 5859 17663
rect 5918 17629 5952 17663
rect 6745 17629 6779 17663
rect 7021 17629 7055 17663
rect 7113 17629 7147 17663
rect 15945 17629 15979 17663
rect 21925 17629 21959 17663
rect 1501 17561 1535 17595
rect 1777 17561 1811 17595
rect 2789 17561 2823 17595
rect 15117 17561 15151 17595
rect 15209 17561 15243 17595
rect 18061 17561 18095 17595
rect 20085 17561 20119 17595
rect 6193 17493 6227 17527
rect 15853 17493 15887 17527
rect 17693 17493 17727 17527
rect 18153 17493 18187 17527
rect 7113 17289 7147 17323
rect 7757 17289 7791 17323
rect 9321 17289 9355 17323
rect 18613 17289 18647 17323
rect 21005 17289 21039 17323
rect 24593 17289 24627 17323
rect 8953 17221 8987 17255
rect 9169 17221 9203 17255
rect 18705 17221 18739 17255
rect 18889 17221 18923 17255
rect 22017 17221 22051 17255
rect 23121 17221 23155 17255
rect 1501 17153 1535 17187
rect 1777 17153 1811 17187
rect 5457 17153 5491 17187
rect 6377 17153 6411 17187
rect 6561 17153 6595 17187
rect 6929 17153 6963 17187
rect 7205 17153 7239 17187
rect 7389 17153 7423 17187
rect 7481 17153 7515 17187
rect 7573 17153 7607 17187
rect 21189 17153 21223 17187
rect 21465 17153 21499 17187
rect 21649 17153 21683 17187
rect 22385 17153 22419 17187
rect 22845 17153 22879 17187
rect 5733 17085 5767 17119
rect 6193 17085 6227 17119
rect 6653 17085 6687 17119
rect 6745 17085 6779 17119
rect 16865 17085 16899 17119
rect 17141 17085 17175 17119
rect 19073 17085 19107 17119
rect 6009 17017 6043 17051
rect 21833 17017 21867 17051
rect 1593 16949 1627 16983
rect 5549 16949 5583 16983
rect 9137 16949 9171 16983
rect 22017 16949 22051 16983
rect 2697 16745 2731 16779
rect 6377 16745 6411 16779
rect 6837 16745 6871 16779
rect 8585 16745 8619 16779
rect 11253 16745 11287 16779
rect 17220 16745 17254 16779
rect 18705 16745 18739 16779
rect 23857 16745 23891 16779
rect 1685 16677 1719 16711
rect 6193 16677 6227 16711
rect 6561 16677 6595 16711
rect 11345 16609 11379 16643
rect 11621 16609 11655 16643
rect 16957 16609 16991 16643
rect 23581 16609 23615 16643
rect 24409 16609 24443 16643
rect 24685 16609 24719 16643
rect 2835 16541 2869 16575
rect 3248 16541 3282 16575
rect 3341 16541 3375 16575
rect 3433 16541 3467 16575
rect 3617 16541 3651 16575
rect 5917 16541 5951 16575
rect 6469 16541 6503 16575
rect 6929 16541 6963 16575
rect 7941 16541 7975 16575
rect 8089 16541 8123 16575
rect 8406 16541 8440 16575
rect 19901 16541 19935 16575
rect 19993 16541 20027 16575
rect 23489 16541 23523 16575
rect 1501 16473 1535 16507
rect 1777 16473 1811 16507
rect 2973 16473 3007 16507
rect 3065 16473 3099 16507
rect 3525 16473 3559 16507
rect 8217 16473 8251 16507
rect 8309 16473 8343 16507
rect 13093 16405 13127 16439
rect 26157 16405 26191 16439
rect 1593 16201 1627 16235
rect 2789 16201 2823 16235
rect 6193 16201 6227 16235
rect 6945 16201 6979 16235
rect 7113 16201 7147 16235
rect 9321 16201 9355 16235
rect 9873 16201 9907 16235
rect 12081 16201 12115 16235
rect 12449 16201 12483 16235
rect 6745 16133 6779 16167
rect 7205 16133 7239 16167
rect 7405 16133 7439 16167
rect 9229 16133 9263 16167
rect 9689 16133 9723 16167
rect 10041 16133 10075 16167
rect 10241 16133 10275 16167
rect 1501 16065 1535 16099
rect 1777 16065 1811 16099
rect 2237 16065 2271 16099
rect 2513 16065 2547 16099
rect 2605 16065 2639 16099
rect 2881 16065 2915 16099
rect 3065 16065 3099 16099
rect 3341 16065 3375 16099
rect 3433 16065 3467 16099
rect 3617 16065 3651 16099
rect 5825 16065 5859 16099
rect 5918 16065 5952 16099
rect 8861 16065 8895 16099
rect 8954 16065 8988 16099
rect 9505 16065 9539 16099
rect 9781 16065 9815 16099
rect 11989 16065 12023 16099
rect 18429 16065 18463 16099
rect 18613 16065 18647 16099
rect 3249 15997 3283 16031
rect 12541 15997 12575 16031
rect 12725 15997 12759 16031
rect 15025 15997 15059 16031
rect 15301 15997 15335 16031
rect 2329 15929 2363 15963
rect 7573 15929 7607 15963
rect 6929 15861 6963 15895
rect 7389 15861 7423 15895
rect 10057 15861 10091 15895
rect 13553 15861 13587 15895
rect 18797 15861 18831 15895
rect 2973 15657 3007 15691
rect 3893 15657 3927 15691
rect 6101 15657 6135 15691
rect 9597 15657 9631 15691
rect 10333 15657 10367 15691
rect 10609 15657 10643 15691
rect 12725 15657 12759 15691
rect 14841 15657 14875 15691
rect 6929 15589 6963 15623
rect 9413 15589 9447 15623
rect 1685 15521 1719 15555
rect 3065 15521 3099 15555
rect 5917 15521 5951 15555
rect 9137 15521 9171 15555
rect 13369 15521 13403 15555
rect 14289 15521 14323 15555
rect 17049 15521 17083 15555
rect 1409 15453 1443 15487
rect 2329 15453 2363 15487
rect 2422 15453 2456 15487
rect 2605 15453 2639 15487
rect 2835 15453 2869 15487
rect 3340 15453 3374 15487
rect 3433 15453 3467 15487
rect 3801 15453 3835 15487
rect 5825 15453 5859 15487
rect 6561 15453 6595 15487
rect 6654 15453 6688 15487
rect 9689 15453 9723 15487
rect 9873 15453 9907 15487
rect 10149 15453 10183 15487
rect 10425 15453 10459 15487
rect 10518 15453 10552 15487
rect 13093 15453 13127 15487
rect 14473 15453 14507 15487
rect 16957 15453 16991 15487
rect 18797 15453 18831 15487
rect 19993 15453 20027 15487
rect 20177 15453 20211 15487
rect 2697 15385 2731 15419
rect 13185 15317 13219 15351
rect 14381 15317 14415 15351
rect 21465 15317 21499 15351
rect 1777 15113 1811 15147
rect 2513 15113 2547 15147
rect 9321 15113 9355 15147
rect 9781 15113 9815 15147
rect 12725 15113 12759 15147
rect 13093 15113 13127 15147
rect 21557 15113 21591 15147
rect 2605 15045 2639 15079
rect 9413 15045 9447 15079
rect 18981 15045 19015 15079
rect 20269 15045 20303 15079
rect 22109 15045 22143 15079
rect 1501 14977 1535 15011
rect 1685 14977 1719 15011
rect 2880 14977 2914 15011
rect 2973 14977 3007 15011
rect 3433 14977 3467 15011
rect 9505 14977 9539 15011
rect 9873 14977 9907 15011
rect 18797 14977 18831 15011
rect 18889 14977 18923 15011
rect 19165 14977 19199 15011
rect 21005 14977 21039 15011
rect 21189 14977 21223 15011
rect 21281 14977 21315 15011
rect 21373 14977 21407 15011
rect 21833 14977 21867 15011
rect 2053 14909 2087 14943
rect 3709 14909 3743 14943
rect 9045 14909 9079 14943
rect 9137 14909 9171 14943
rect 9965 14909 9999 14943
rect 13185 14909 13219 14943
rect 13369 14909 13403 14943
rect 2329 14841 2363 14875
rect 18613 14773 18647 14807
rect 23581 14773 23615 14807
rect 1685 14569 1719 14603
rect 4261 14569 4295 14603
rect 16129 14569 16163 14603
rect 16221 14569 16255 14603
rect 1593 14501 1627 14535
rect 19257 14501 19291 14535
rect 15485 14433 15519 14467
rect 16773 14433 16807 14467
rect 17325 14433 17359 14467
rect 17601 14433 17635 14467
rect 21373 14433 21407 14467
rect 1409 14365 1443 14399
rect 1869 14365 1903 14399
rect 2973 14365 3007 14399
rect 3341 14365 3375 14399
rect 3801 14365 3835 14399
rect 4077 14365 4111 14399
rect 19441 14365 19475 14399
rect 19625 14365 19659 14399
rect 19809 14365 19843 14399
rect 20729 14365 20763 14399
rect 20913 14365 20947 14399
rect 21097 14365 21131 14399
rect 3157 14297 3191 14331
rect 3249 14297 3283 14331
rect 15669 14297 15703 14331
rect 16681 14297 16715 14331
rect 19533 14297 19567 14331
rect 21005 14297 21039 14331
rect 21649 14297 21683 14331
rect 3525 14229 3559 14263
rect 3893 14229 3927 14263
rect 15209 14229 15243 14263
rect 15761 14229 15795 14263
rect 16589 14229 16623 14263
rect 19073 14229 19107 14263
rect 21281 14229 21315 14263
rect 23121 14229 23155 14263
rect 3525 14025 3559 14059
rect 3617 14025 3651 14059
rect 8401 14025 8435 14059
rect 9597 14025 9631 14059
rect 11989 14025 12023 14059
rect 19441 14025 19475 14059
rect 21925 14025 21959 14059
rect 23397 14025 23431 14059
rect 1685 13957 1719 13991
rect 8033 13957 8067 13991
rect 9229 13957 9263 13991
rect 9445 13957 9479 13991
rect 17969 13957 18003 13991
rect 1501 13889 1535 13923
rect 1777 13889 1811 13923
rect 2973 13889 3007 13923
rect 3249 13889 3283 13923
rect 3341 13889 3375 13923
rect 3801 13889 3835 13923
rect 3893 13889 3927 13923
rect 4077 13889 4111 13923
rect 4169 13889 4203 13923
rect 6469 13889 6503 13923
rect 6623 13889 6657 13923
rect 7757 13889 7791 13923
rect 7905 13889 7939 13923
rect 8125 13889 8159 13923
rect 8222 13889 8256 13923
rect 12449 13889 12483 13923
rect 14197 13889 14231 13923
rect 17693 13889 17727 13923
rect 22293 13889 22327 13923
rect 23489 13889 23523 13923
rect 23949 13889 23983 13923
rect 12541 13821 12575 13855
rect 12633 13821 12667 13855
rect 14473 13821 14507 13855
rect 15945 13821 15979 13855
rect 16129 13821 16163 13855
rect 22385 13821 22419 13855
rect 22477 13821 22511 13855
rect 23213 13821 23247 13855
rect 24225 13821 24259 13855
rect 25697 13821 25731 13855
rect 6837 13753 6871 13787
rect 3065 13685 3099 13719
rect 9413 13685 9447 13719
rect 12081 13685 12115 13719
rect 23857 13685 23891 13719
rect 3525 13481 3559 13515
rect 4537 13481 4571 13515
rect 6837 13481 6871 13515
rect 7021 13481 7055 13515
rect 7297 13481 7331 13515
rect 7665 13481 7699 13515
rect 8953 13481 8987 13515
rect 14473 13481 14507 13515
rect 24409 13481 24443 13515
rect 7481 13413 7515 13447
rect 1685 13345 1719 13379
rect 4077 13345 4111 13379
rect 4261 13345 4295 13379
rect 6469 13345 6503 13379
rect 8769 13345 8803 13379
rect 9229 13345 9263 13379
rect 15025 13345 15059 13379
rect 24869 13345 24903 13379
rect 24961 13345 24995 13379
rect 1409 13277 1443 13311
rect 3617 13277 3651 13311
rect 3985 13277 4019 13311
rect 4169 13277 4203 13311
rect 4445 13277 4479 13311
rect 6009 13277 6043 13311
rect 6163 13277 6197 13311
rect 7573 13277 7607 13311
rect 8401 13277 8435 13311
rect 8494 13277 8528 13311
rect 9137 13277 9171 13311
rect 9689 13277 9723 13311
rect 9903 13277 9937 13311
rect 10057 13277 10091 13311
rect 11345 13277 11379 13311
rect 13001 13277 13035 13311
rect 14841 13277 14875 13311
rect 24777 13277 24811 13311
rect 6377 13209 6411 13243
rect 6837 13209 6871 13243
rect 7113 13209 7147 13243
rect 11437 13209 11471 13243
rect 13277 13209 13311 13243
rect 14933 13209 14967 13243
rect 3801 13141 3835 13175
rect 7313 13141 7347 13175
rect 9597 13141 9631 13175
rect 13461 13141 13495 13175
rect 1685 12937 1719 12971
rect 3433 12937 3467 12971
rect 6929 12937 6963 12971
rect 9229 12937 9263 12971
rect 13277 12937 13311 12971
rect 15853 12937 15887 12971
rect 19165 12937 19199 12971
rect 19809 12937 19843 12971
rect 2421 12869 2455 12903
rect 11805 12869 11839 12903
rect 15761 12869 15795 12903
rect 19073 12869 19107 12903
rect 19901 12869 19935 12903
rect 1409 12801 1443 12835
rect 1869 12801 1903 12835
rect 2635 12801 2669 12835
rect 2789 12801 2823 12835
rect 3065 12801 3099 12835
rect 6561 12801 6595 12835
rect 8861 12801 8895 12835
rect 8954 12801 8988 12835
rect 11529 12801 11563 12835
rect 13369 12801 13403 12835
rect 13645 12801 13679 12835
rect 3157 12733 3191 12767
rect 6469 12733 6503 12767
rect 19257 12733 19291 12767
rect 19717 12733 19751 12767
rect 1593 12665 1627 12699
rect 3249 12597 3283 12631
rect 11345 12597 11379 12631
rect 16773 12597 16807 12631
rect 18705 12597 18739 12631
rect 20269 12597 20303 12631
rect 3065 12393 3099 12427
rect 12817 12393 12851 12427
rect 2973 12325 3007 12359
rect 11897 12325 11931 12359
rect 12725 12325 12759 12359
rect 21925 12325 21959 12359
rect 24685 12325 24719 12359
rect 1961 12257 1995 12291
rect 12173 12257 12207 12291
rect 13461 12257 13495 12291
rect 14933 12257 14967 12291
rect 23673 12257 23707 12291
rect 23857 12257 23891 12291
rect 2237 12189 2271 12223
rect 2329 12189 2363 12223
rect 4261 12189 4295 12223
rect 11713 12189 11747 12223
rect 13277 12189 13311 12223
rect 16773 12189 16807 12223
rect 17049 12189 17083 12223
rect 24501 12189 24535 12223
rect 2605 12121 2639 12155
rect 15209 12121 15243 12155
rect 21741 12121 21775 12155
rect 4169 12053 4203 12087
rect 12265 12053 12299 12087
rect 12357 12053 12391 12087
rect 13185 12053 13219 12087
rect 16681 12053 16715 12087
rect 23213 12053 23247 12087
rect 23581 12053 23615 12087
rect 2421 11849 2455 11883
rect 9321 11849 9355 11883
rect 15301 11849 15335 11883
rect 16221 11849 16255 11883
rect 18797 11849 18831 11883
rect 22293 11849 22327 11883
rect 24777 11849 24811 11883
rect 15669 11781 15703 11815
rect 23305 11781 23339 11815
rect 1961 11713 1995 11747
rect 2329 11713 2363 11747
rect 2881 11713 2915 11747
rect 13277 11713 13311 11747
rect 16313 11713 16347 11747
rect 16957 11713 16991 11747
rect 18705 11713 18739 11747
rect 22201 11713 22235 11747
rect 2237 11645 2271 11679
rect 2605 11645 2639 11679
rect 3157 11645 3191 11679
rect 9413 11645 9447 11679
rect 9689 11645 9723 11679
rect 15761 11645 15795 11679
rect 15945 11645 15979 11679
rect 16681 11645 16715 11679
rect 18889 11645 18923 11679
rect 22385 11645 22419 11679
rect 23029 11645 23063 11679
rect 13093 11577 13127 11611
rect 3249 11509 3283 11543
rect 3433 11509 3467 11543
rect 11161 11509 11195 11543
rect 14565 11509 14599 11543
rect 15117 11509 15151 11543
rect 18337 11509 18371 11543
rect 21833 11509 21867 11543
rect 1593 11305 1627 11339
rect 2329 11305 2363 11339
rect 3157 11305 3191 11339
rect 3801 11305 3835 11339
rect 14473 11305 14507 11339
rect 16037 11305 16071 11339
rect 19073 11305 19107 11339
rect 4629 11237 4663 11271
rect 2053 11169 2087 11203
rect 4537 11169 4571 11203
rect 4721 11169 4755 11203
rect 15025 11169 15059 11203
rect 15393 11169 15427 11203
rect 17601 11169 17635 11203
rect 19993 11169 20027 11203
rect 20085 11169 20119 11203
rect 22385 11169 22419 11203
rect 24869 11169 24903 11203
rect 24961 11169 24995 11203
rect 1409 11101 1443 11135
rect 1961 11101 1995 11135
rect 3341 11101 3375 11135
rect 3617 11101 3651 11135
rect 3985 11101 4019 11135
rect 4077 11101 4111 11135
rect 4261 11101 4295 11135
rect 4353 11101 4387 11135
rect 4445 11101 4479 11135
rect 4813 11101 4847 11135
rect 8677 11101 8711 11135
rect 16589 11101 16623 11135
rect 17325 11101 17359 11135
rect 10701 11033 10735 11067
rect 10885 11033 10919 11067
rect 14105 11033 14139 11067
rect 14289 11033 14323 11067
rect 14841 11033 14875 11067
rect 15669 11033 15703 11067
rect 19901 11033 19935 11067
rect 22109 11033 22143 11067
rect 24777 11033 24811 11067
rect 3525 10965 3559 10999
rect 9413 10965 9447 10999
rect 14933 10965 14967 10999
rect 15577 10965 15611 10999
rect 19533 10965 19567 10999
rect 20637 10965 20671 10999
rect 24409 10965 24443 10999
rect 1685 10761 1719 10795
rect 3617 10761 3651 10795
rect 4077 10761 4111 10795
rect 9689 10761 9723 10795
rect 10057 10761 10091 10795
rect 20821 10761 20855 10795
rect 21281 10761 21315 10795
rect 24685 10761 24719 10795
rect 20913 10693 20947 10727
rect 23857 10693 23891 10727
rect 1409 10625 1443 10659
rect 1869 10625 1903 10659
rect 3249 10625 3283 10659
rect 3342 10625 3376 10659
rect 3709 10625 3743 10659
rect 3863 10625 3897 10659
rect 9045 10625 9079 10659
rect 11529 10625 11563 10659
rect 13829 10625 13863 10659
rect 19257 10625 19291 10659
rect 23765 10625 23799 10659
rect 24593 10625 24627 10659
rect 6377 10557 6411 10591
rect 6653 10557 6687 10591
rect 8861 10557 8895 10591
rect 8953 10557 8987 10591
rect 10149 10557 10183 10591
rect 10333 10557 10367 10591
rect 11805 10557 11839 10591
rect 14105 10557 14139 10591
rect 15577 10557 15611 10591
rect 20729 10557 20763 10591
rect 23949 10557 23983 10591
rect 24777 10557 24811 10591
rect 1593 10489 1627 10523
rect 9413 10489 9447 10523
rect 8125 10421 8159 10455
rect 9597 10421 9631 10455
rect 13277 10421 13311 10455
rect 19441 10421 19475 10455
rect 23397 10421 23431 10455
rect 24225 10421 24259 10455
rect 1593 10217 1627 10251
rect 6763 10217 6797 10251
rect 7113 10217 7147 10251
rect 11621 10217 11655 10251
rect 14105 10217 14139 10251
rect 7573 10081 7607 10115
rect 7665 10081 7699 10115
rect 8769 10081 8803 10115
rect 9137 10081 9171 10115
rect 12173 10081 12207 10115
rect 14749 10081 14783 10115
rect 19717 10081 19751 10115
rect 19901 10081 19935 10115
rect 1409 10013 1443 10047
rect 1685 10013 1719 10047
rect 7021 10013 7055 10047
rect 11989 10013 12023 10047
rect 14473 10013 14507 10047
rect 7481 9945 7515 9979
rect 9321 9945 9355 9979
rect 14565 9945 14599 9979
rect 5273 9877 5307 9911
rect 9229 9877 9263 9911
rect 9689 9877 9723 9911
rect 12081 9877 12115 9911
rect 19257 9877 19291 9911
rect 19625 9877 19659 9911
rect 1593 9673 1627 9707
rect 7113 9673 7147 9707
rect 12265 9673 12299 9707
rect 19625 9673 19659 9707
rect 22477 9673 22511 9707
rect 6745 9605 6779 9639
rect 18153 9605 18187 9639
rect 23673 9605 23707 9639
rect 1409 9537 1443 9571
rect 1685 9537 1719 9571
rect 11897 9537 11931 9571
rect 14381 9537 14415 9571
rect 17877 9537 17911 9571
rect 22385 9537 22419 9571
rect 6561 9469 6595 9503
rect 6653 9469 6687 9503
rect 11621 9469 11655 9503
rect 11805 9469 11839 9503
rect 14105 9469 14139 9503
rect 14289 9469 14323 9503
rect 22661 9469 22695 9503
rect 23397 9469 23431 9503
rect 25145 9469 25179 9503
rect 11253 9333 11287 9367
rect 14749 9333 14783 9367
rect 22017 9333 22051 9367
rect 3985 9129 4019 9163
rect 7297 9129 7331 9163
rect 12449 9129 12483 9163
rect 15853 9129 15887 9163
rect 20453 9129 20487 9163
rect 3525 9061 3559 9095
rect 7205 8993 7239 9027
rect 7849 8993 7883 9027
rect 9873 8993 9907 9027
rect 11805 8993 11839 9027
rect 11989 8993 12023 9027
rect 14381 8993 14415 9027
rect 1777 8925 1811 8959
rect 4169 8925 4203 8959
rect 14105 8925 14139 8959
rect 20637 8925 20671 8959
rect 22937 8925 22971 8959
rect 2053 8857 2087 8891
rect 3893 8857 3927 8891
rect 10149 8857 10183 8891
rect 12081 8857 12115 8891
rect 1409 8789 1443 8823
rect 4353 8789 4387 8823
rect 4537 8789 4571 8823
rect 7665 8789 7699 8823
rect 7757 8789 7791 8823
rect 11621 8789 11655 8823
rect 21925 8789 21959 8823
rect 23121 8789 23155 8823
rect 2605 8585 2639 8619
rect 2973 8585 3007 8619
rect 4261 8585 4295 8619
rect 7941 8585 7975 8619
rect 10241 8585 10275 8619
rect 10609 8585 10643 8619
rect 20821 8585 20855 8619
rect 24317 8585 24351 8619
rect 8033 8517 8067 8551
rect 19533 8517 19567 8551
rect 22109 8517 22143 8551
rect 1409 8449 1443 8483
rect 3065 8449 3099 8483
rect 3801 8449 3835 8483
rect 3893 8449 3927 8483
rect 4353 8449 4387 8483
rect 11529 8449 11563 8483
rect 24409 8449 24443 8483
rect 1685 8381 1719 8415
rect 3249 8381 3283 8415
rect 3617 8381 3651 8415
rect 7849 8381 7883 8415
rect 10701 8381 10735 8415
rect 10885 8381 10919 8415
rect 17693 8381 17727 8415
rect 19165 8381 19199 8415
rect 19441 8381 19475 8415
rect 21833 8381 21867 8415
rect 24225 8381 24259 8415
rect 4537 8313 4571 8347
rect 7481 8313 7515 8347
rect 8401 8313 8435 8347
rect 23581 8313 23615 8347
rect 24777 8245 24811 8279
rect 3801 8041 3835 8075
rect 8217 8041 8251 8075
rect 17601 8041 17635 8075
rect 19349 8041 19383 8075
rect 19533 8041 19567 8075
rect 27905 8041 27939 8075
rect 2513 7973 2547 8007
rect 17969 7973 18003 8007
rect 1409 7905 1443 7939
rect 1685 7905 1719 7939
rect 4353 7905 4387 7939
rect 4721 7905 4755 7939
rect 17325 7905 17359 7939
rect 20085 7905 20119 7939
rect 20913 7905 20947 7939
rect 21281 7905 21315 7939
rect 24685 7905 24719 7939
rect 2329 7837 2363 7871
rect 2605 7837 2639 7871
rect 6469 7837 6503 7871
rect 17785 7837 17819 7871
rect 18153 7837 18187 7871
rect 20821 7837 20855 7871
rect 21465 7837 21499 7871
rect 24409 7837 24443 7871
rect 28089 7837 28123 7871
rect 4261 7769 4295 7803
rect 6745 7769 6779 7803
rect 17049 7769 17083 7803
rect 17509 7769 17543 7803
rect 20729 7769 20763 7803
rect 21557 7769 21591 7803
rect 28365 7769 28399 7803
rect 4169 7701 4203 7735
rect 15577 7701 15611 7735
rect 19901 7701 19935 7735
rect 19993 7701 20027 7735
rect 20361 7701 20395 7735
rect 21925 7701 21959 7735
rect 26157 7701 26191 7735
rect 1409 7497 1443 7531
rect 7205 7497 7239 7531
rect 7573 7497 7607 7531
rect 8861 7497 8895 7531
rect 14749 7497 14783 7531
rect 15393 7497 15427 7531
rect 16681 7497 16715 7531
rect 17141 7497 17175 7531
rect 18429 7497 18463 7531
rect 18889 7497 18923 7531
rect 24869 7497 24903 7531
rect 24961 7497 24995 7531
rect 14841 7429 14875 7463
rect 15301 7429 15335 7463
rect 24041 7429 24075 7463
rect 1593 7361 1627 7395
rect 3801 7361 3835 7395
rect 4353 7361 4387 7395
rect 14565 7361 14599 7395
rect 15025 7361 15059 7395
rect 15577 7361 15611 7395
rect 15853 7361 15887 7395
rect 17049 7361 17083 7395
rect 18797 7361 18831 7395
rect 24133 7361 24167 7395
rect 1869 7293 1903 7327
rect 3893 7293 3927 7327
rect 3985 7293 4019 7327
rect 4629 7293 4663 7327
rect 7665 7293 7699 7327
rect 7849 7293 7883 7327
rect 17325 7293 17359 7327
rect 18981 7293 19015 7327
rect 21833 7293 21867 7327
rect 22109 7293 22143 7327
rect 24225 7293 24259 7327
rect 25053 7293 25087 7327
rect 3433 7225 3467 7259
rect 15761 7225 15795 7259
rect 3341 7157 3375 7191
rect 6101 7157 6135 7191
rect 14381 7157 14415 7191
rect 23581 7157 23615 7191
rect 23673 7157 23707 7191
rect 24501 7157 24535 7191
rect 4813 6953 4847 6987
rect 22201 6953 22235 6987
rect 1961 6885 1995 6919
rect 5457 6817 5491 6851
rect 7021 6817 7055 6851
rect 13093 6817 13127 6851
rect 14105 6817 14139 6851
rect 19717 6817 19751 6851
rect 19901 6817 19935 6851
rect 22753 6817 22787 6851
rect 1777 6749 1811 6783
rect 2237 6749 2271 6783
rect 5181 6749 5215 6783
rect 10701 6749 10735 6783
rect 10977 6749 11011 6783
rect 22569 6749 22603 6783
rect 22661 6749 22695 6783
rect 1501 6681 1535 6715
rect 1685 6681 1719 6715
rect 2053 6681 2087 6715
rect 8769 6681 8803 6715
rect 10425 6681 10459 6715
rect 12817 6681 12851 6715
rect 13737 6681 13771 6715
rect 14381 6681 14415 6715
rect 19625 6681 19659 6715
rect 2421 6613 2455 6647
rect 5273 6613 5307 6647
rect 8953 6613 8987 6647
rect 11345 6613 11379 6647
rect 13829 6613 13863 6647
rect 15853 6613 15887 6647
rect 19257 6613 19291 6647
rect 7849 6409 7883 6443
rect 8861 6409 8895 6443
rect 14381 6409 14415 6443
rect 14749 6409 14783 6443
rect 14841 6409 14875 6443
rect 16681 6409 16715 6443
rect 17141 6409 17175 6443
rect 21189 6409 21223 6443
rect 7113 6341 7147 6375
rect 11529 6341 11563 6375
rect 13369 6341 13403 6375
rect 14013 6341 14047 6375
rect 21281 6341 21315 6375
rect 1501 6273 1535 6307
rect 1961 6273 1995 6307
rect 8217 6273 8251 6307
rect 9965 6273 9999 6307
rect 10977 6273 11011 6307
rect 13277 6273 13311 6307
rect 13921 6273 13955 6307
rect 15209 6273 15243 6307
rect 17049 6273 17083 6307
rect 3249 6205 3283 6239
rect 8309 6205 8343 6239
rect 8493 6205 8527 6239
rect 9505 6205 9539 6239
rect 9781 6205 9815 6239
rect 9873 6205 9907 6239
rect 11069 6205 11103 6239
rect 11253 6205 11287 6239
rect 14197 6205 14231 6239
rect 14933 6205 14967 6239
rect 17325 6205 17359 6239
rect 1685 6137 1719 6171
rect 1869 6137 1903 6171
rect 7757 6137 7791 6171
rect 10333 6137 10367 6171
rect 10609 6137 10643 6171
rect 15577 6137 15611 6171
rect 3709 6069 3743 6103
rect 13553 6069 13587 6103
rect 15393 6069 15427 6103
rect 2973 5865 3007 5899
rect 5549 5865 5583 5899
rect 7573 5865 7607 5899
rect 12173 5865 12207 5899
rect 12265 5865 12299 5899
rect 2237 5797 2271 5831
rect 2421 5797 2455 5831
rect 2697 5797 2731 5831
rect 14105 5797 14139 5831
rect 4997 5729 5031 5763
rect 8033 5729 8067 5763
rect 8125 5729 8159 5763
rect 10793 5729 10827 5763
rect 11437 5729 11471 5763
rect 12817 5729 12851 5763
rect 14565 5729 14599 5763
rect 14657 5729 14691 5763
rect 16681 5729 16715 5763
rect 18521 5729 18555 5763
rect 18613 5729 18647 5763
rect 21649 5729 21683 5763
rect 1409 5661 1443 5695
rect 1685 5661 1719 5695
rect 2513 5661 2547 5695
rect 2789 5661 2823 5695
rect 3525 5661 3559 5695
rect 4077 5661 4111 5695
rect 4445 5661 4479 5695
rect 7941 5661 7975 5695
rect 11345 5661 11379 5695
rect 12633 5661 12667 5695
rect 12725 5661 12759 5695
rect 14473 5661 14507 5695
rect 16497 5661 16531 5695
rect 21833 5661 21867 5695
rect 3341 5593 3375 5627
rect 4261 5593 4295 5627
rect 16405 5593 16439 5627
rect 21373 5593 21407 5627
rect 22017 5593 22051 5627
rect 1593 5525 1627 5559
rect 3893 5525 3927 5559
rect 5089 5525 5123 5559
rect 5181 5525 5215 5559
rect 5733 5525 5767 5559
rect 10885 5525 10919 5559
rect 11253 5525 11287 5559
rect 16037 5525 16071 5559
rect 18061 5525 18095 5559
rect 18429 5525 18463 5559
rect 19901 5525 19935 5559
rect 1593 5321 1627 5355
rect 3249 5321 3283 5355
rect 3709 5321 3743 5355
rect 5181 5321 5215 5355
rect 19165 5321 19199 5355
rect 21189 5321 21223 5355
rect 21557 5321 21591 5355
rect 2145 5253 2179 5287
rect 3617 5253 3651 5287
rect 6193 5253 6227 5287
rect 17693 5253 17727 5287
rect 1409 5185 1443 5219
rect 1685 5185 1719 5219
rect 2697 5185 2731 5219
rect 3065 5185 3099 5219
rect 3433 5185 3467 5219
rect 4353 5185 4387 5219
rect 5089 5185 5123 5219
rect 5549 5185 5583 5219
rect 17417 5185 17451 5219
rect 25053 5185 25087 5219
rect 4077 5117 4111 5151
rect 5365 5117 5399 5151
rect 20913 5117 20947 5151
rect 21097 5117 21131 5151
rect 24777 5117 24811 5151
rect 2329 5049 2363 5083
rect 2881 5049 2915 5083
rect 2513 4981 2547 5015
rect 4261 4981 4295 5015
rect 4537 4981 4571 5015
rect 4721 4981 4755 5015
rect 5733 4981 5767 5015
rect 6009 4981 6043 5015
rect 23305 4981 23339 5015
rect 3157 4777 3191 4811
rect 8677 4777 8711 4811
rect 18153 4777 18187 4811
rect 18521 4777 18555 4811
rect 21925 4777 21959 4811
rect 25145 4777 25179 4811
rect 3525 4709 3559 4743
rect 1409 4641 1443 4675
rect 3801 4641 3835 4675
rect 4077 4641 4111 4675
rect 6929 4641 6963 4675
rect 14841 4641 14875 4675
rect 15209 4641 15243 4675
rect 22569 4641 22603 4675
rect 24501 4641 24535 4675
rect 24685 4641 24719 4675
rect 3249 4573 3283 4607
rect 14749 4573 14783 4607
rect 18337 4573 18371 4607
rect 22293 4573 22327 4607
rect 24777 4573 24811 4607
rect 1685 4505 1719 4539
rect 7205 4505 7239 4539
rect 15393 4505 15427 4539
rect 5549 4437 5583 4471
rect 14289 4437 14323 4471
rect 14657 4437 14691 4471
rect 15485 4437 15519 4471
rect 15853 4437 15887 4471
rect 22385 4437 22419 4471
rect 2605 4233 2639 4267
rect 2973 4233 3007 4267
rect 4629 4233 4663 4267
rect 7481 4233 7515 4267
rect 7849 4233 7883 4267
rect 17877 4233 17911 4267
rect 18337 4233 18371 4267
rect 19165 4233 19199 4267
rect 22201 4233 22235 4267
rect 23029 4233 23063 4267
rect 4537 4165 4571 4199
rect 8677 4165 8711 4199
rect 10885 4165 10919 4199
rect 11897 4165 11931 4199
rect 11989 4165 12023 4199
rect 15669 4165 15703 4199
rect 18245 4165 18279 4199
rect 19073 4165 19107 4199
rect 23121 4165 23155 4199
rect 5089 4097 5123 4131
rect 12449 4097 12483 4131
rect 15945 4097 15979 4131
rect 22293 4097 22327 4131
rect 3065 4029 3099 4063
rect 3249 4029 3283 4063
rect 4813 4029 4847 4063
rect 7941 4029 7975 4063
rect 8125 4029 8159 4063
rect 8769 4029 8803 4063
rect 8953 4029 8987 4063
rect 10701 4029 10735 4063
rect 10793 4029 10827 4063
rect 12081 4029 12115 4063
rect 14197 4029 14231 4063
rect 18521 4029 18555 4063
rect 19257 4029 19291 4063
rect 22385 4029 22419 4063
rect 23305 4029 23339 4063
rect 4169 3961 4203 3995
rect 8309 3961 8343 3995
rect 11253 3893 11287 3927
rect 11529 3893 11563 3927
rect 18705 3893 18739 3927
rect 21833 3893 21867 3927
rect 22661 3893 22695 3927
rect 5549 3689 5583 3723
rect 8493 3689 8527 3723
rect 10425 3689 10459 3723
rect 12265 3689 12299 3723
rect 15853 3689 15887 3723
rect 18613 3689 18647 3723
rect 22845 3689 22879 3723
rect 3801 3553 3835 3587
rect 6561 3553 6595 3587
rect 8769 3553 8803 3587
rect 9597 3553 9631 3587
rect 11897 3553 11931 3587
rect 12725 3553 12759 3587
rect 12817 3553 12851 3587
rect 14105 3553 14139 3587
rect 14381 3553 14415 3587
rect 18061 3553 18095 3587
rect 19257 3553 19291 3587
rect 21097 3553 21131 3587
rect 9321 3485 9355 3519
rect 12173 3485 12207 3519
rect 18429 3485 18463 3519
rect 4077 3417 4111 3451
rect 6837 3417 6871 3451
rect 9413 3417 9447 3451
rect 17785 3417 17819 3451
rect 19533 3417 19567 3451
rect 21373 3417 21407 3451
rect 8309 3349 8343 3383
rect 8953 3349 8987 3383
rect 12633 3349 12667 3383
rect 16313 3349 16347 3383
rect 18245 3349 18279 3383
rect 21005 3349 21039 3383
rect 4445 3145 4479 3179
rect 4813 3145 4847 3179
rect 7573 3145 7607 3179
rect 7941 3145 7975 3179
rect 9505 3145 9539 3179
rect 12173 3145 12207 3179
rect 12541 3145 12575 3179
rect 17509 3145 17543 3179
rect 17877 3145 17911 3179
rect 20085 3145 20119 3179
rect 20453 3145 20487 3179
rect 20545 3145 20579 3179
rect 4905 3077 4939 3111
rect 10977 3077 11011 3111
rect 17417 3077 17451 3111
rect 8033 3009 8067 3043
rect 11253 3009 11287 3043
rect 12633 3009 12667 3043
rect 5089 2941 5123 2975
rect 8125 2941 8159 2975
rect 12081 2941 12115 2975
rect 12725 2941 12759 2975
rect 17233 2941 17267 2975
rect 20729 2941 20763 2975
<< metal1 >>
rect 1104 27770 28888 27792
rect 1104 27718 2918 27770
rect 2970 27718 2982 27770
rect 3034 27718 3046 27770
rect 3098 27718 3110 27770
rect 3162 27718 3174 27770
rect 3226 27718 3238 27770
rect 3290 27718 10918 27770
rect 10970 27718 10982 27770
rect 11034 27718 11046 27770
rect 11098 27718 11110 27770
rect 11162 27718 11174 27770
rect 11226 27718 11238 27770
rect 11290 27718 18918 27770
rect 18970 27718 18982 27770
rect 19034 27718 19046 27770
rect 19098 27718 19110 27770
rect 19162 27718 19174 27770
rect 19226 27718 19238 27770
rect 19290 27718 26918 27770
rect 26970 27718 26982 27770
rect 27034 27718 27046 27770
rect 27098 27718 27110 27770
rect 27162 27718 27174 27770
rect 27226 27718 27238 27770
rect 27290 27718 28888 27770
rect 1104 27696 28888 27718
rect 1104 27226 28888 27248
rect 1104 27174 3658 27226
rect 3710 27174 3722 27226
rect 3774 27174 3786 27226
rect 3838 27174 3850 27226
rect 3902 27174 3914 27226
rect 3966 27174 3978 27226
rect 4030 27174 11658 27226
rect 11710 27174 11722 27226
rect 11774 27174 11786 27226
rect 11838 27174 11850 27226
rect 11902 27174 11914 27226
rect 11966 27174 11978 27226
rect 12030 27174 19658 27226
rect 19710 27174 19722 27226
rect 19774 27174 19786 27226
rect 19838 27174 19850 27226
rect 19902 27174 19914 27226
rect 19966 27174 19978 27226
rect 20030 27174 27658 27226
rect 27710 27174 27722 27226
rect 27774 27174 27786 27226
rect 27838 27174 27850 27226
rect 27902 27174 27914 27226
rect 27966 27174 27978 27226
rect 28030 27174 28888 27226
rect 1104 27152 28888 27174
rect 1104 26682 28888 26704
rect 1104 26630 2918 26682
rect 2970 26630 2982 26682
rect 3034 26630 3046 26682
rect 3098 26630 3110 26682
rect 3162 26630 3174 26682
rect 3226 26630 3238 26682
rect 3290 26630 10918 26682
rect 10970 26630 10982 26682
rect 11034 26630 11046 26682
rect 11098 26630 11110 26682
rect 11162 26630 11174 26682
rect 11226 26630 11238 26682
rect 11290 26630 18918 26682
rect 18970 26630 18982 26682
rect 19034 26630 19046 26682
rect 19098 26630 19110 26682
rect 19162 26630 19174 26682
rect 19226 26630 19238 26682
rect 19290 26630 26918 26682
rect 26970 26630 26982 26682
rect 27034 26630 27046 26682
rect 27098 26630 27110 26682
rect 27162 26630 27174 26682
rect 27226 26630 27238 26682
rect 27290 26630 28888 26682
rect 1104 26608 28888 26630
rect 1104 26138 28888 26160
rect 1104 26086 3658 26138
rect 3710 26086 3722 26138
rect 3774 26086 3786 26138
rect 3838 26086 3850 26138
rect 3902 26086 3914 26138
rect 3966 26086 3978 26138
rect 4030 26086 11658 26138
rect 11710 26086 11722 26138
rect 11774 26086 11786 26138
rect 11838 26086 11850 26138
rect 11902 26086 11914 26138
rect 11966 26086 11978 26138
rect 12030 26086 19658 26138
rect 19710 26086 19722 26138
rect 19774 26086 19786 26138
rect 19838 26086 19850 26138
rect 19902 26086 19914 26138
rect 19966 26086 19978 26138
rect 20030 26086 27658 26138
rect 27710 26086 27722 26138
rect 27774 26086 27786 26138
rect 27838 26086 27850 26138
rect 27902 26086 27914 26138
rect 27966 26086 27978 26138
rect 28030 26086 28888 26138
rect 1104 26064 28888 26086
rect 1104 25594 28888 25616
rect 1104 25542 2918 25594
rect 2970 25542 2982 25594
rect 3034 25542 3046 25594
rect 3098 25542 3110 25594
rect 3162 25542 3174 25594
rect 3226 25542 3238 25594
rect 3290 25542 10918 25594
rect 10970 25542 10982 25594
rect 11034 25542 11046 25594
rect 11098 25542 11110 25594
rect 11162 25542 11174 25594
rect 11226 25542 11238 25594
rect 11290 25542 18918 25594
rect 18970 25542 18982 25594
rect 19034 25542 19046 25594
rect 19098 25542 19110 25594
rect 19162 25542 19174 25594
rect 19226 25542 19238 25594
rect 19290 25542 26918 25594
rect 26970 25542 26982 25594
rect 27034 25542 27046 25594
rect 27098 25542 27110 25594
rect 27162 25542 27174 25594
rect 27226 25542 27238 25594
rect 27290 25542 28888 25594
rect 1104 25520 28888 25542
rect 1210 25168 1216 25220
rect 1268 25208 1274 25220
rect 1489 25211 1547 25217
rect 1489 25208 1501 25211
rect 1268 25180 1501 25208
rect 1268 25168 1274 25180
rect 1489 25177 1501 25180
rect 1535 25208 1547 25211
rect 1765 25211 1823 25217
rect 1765 25208 1777 25211
rect 1535 25180 1777 25208
rect 1535 25177 1547 25180
rect 1489 25171 1547 25177
rect 1765 25177 1777 25180
rect 1811 25177 1823 25211
rect 1765 25171 1823 25177
rect 1581 25143 1639 25149
rect 1581 25109 1593 25143
rect 1627 25140 1639 25143
rect 2498 25140 2504 25152
rect 1627 25112 2504 25140
rect 1627 25109 1639 25112
rect 1581 25103 1639 25109
rect 2498 25100 2504 25112
rect 2556 25100 2562 25152
rect 1104 25050 28888 25072
rect 1104 24998 3658 25050
rect 3710 24998 3722 25050
rect 3774 24998 3786 25050
rect 3838 24998 3850 25050
rect 3902 24998 3914 25050
rect 3966 24998 3978 25050
rect 4030 24998 11658 25050
rect 11710 24998 11722 25050
rect 11774 24998 11786 25050
rect 11838 24998 11850 25050
rect 11902 24998 11914 25050
rect 11966 24998 11978 25050
rect 12030 24998 19658 25050
rect 19710 24998 19722 25050
rect 19774 24998 19786 25050
rect 19838 24998 19850 25050
rect 19902 24998 19914 25050
rect 19966 24998 19978 25050
rect 20030 24998 27658 25050
rect 27710 24998 27722 25050
rect 27774 24998 27786 25050
rect 27838 24998 27850 25050
rect 27902 24998 27914 25050
rect 27966 24998 27978 25050
rect 28030 24998 28888 25050
rect 1104 24976 28888 24998
rect 1302 24760 1308 24812
rect 1360 24800 1366 24812
rect 1489 24803 1547 24809
rect 1489 24800 1501 24803
rect 1360 24772 1501 24800
rect 1360 24760 1366 24772
rect 1489 24769 1501 24772
rect 1535 24800 1547 24803
rect 1765 24803 1823 24809
rect 1765 24800 1777 24803
rect 1535 24772 1777 24800
rect 1535 24769 1547 24772
rect 1489 24763 1547 24769
rect 1765 24769 1777 24772
rect 1811 24769 1823 24803
rect 1765 24763 1823 24769
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24596 1639 24599
rect 2682 24596 2688 24608
rect 1627 24568 2688 24596
rect 1627 24565 1639 24568
rect 1581 24559 1639 24565
rect 2682 24556 2688 24568
rect 2740 24556 2746 24608
rect 1104 24506 28888 24528
rect 1104 24454 2918 24506
rect 2970 24454 2982 24506
rect 3034 24454 3046 24506
rect 3098 24454 3110 24506
rect 3162 24454 3174 24506
rect 3226 24454 3238 24506
rect 3290 24454 10918 24506
rect 10970 24454 10982 24506
rect 11034 24454 11046 24506
rect 11098 24454 11110 24506
rect 11162 24454 11174 24506
rect 11226 24454 11238 24506
rect 11290 24454 18918 24506
rect 18970 24454 18982 24506
rect 19034 24454 19046 24506
rect 19098 24454 19110 24506
rect 19162 24454 19174 24506
rect 19226 24454 19238 24506
rect 19290 24454 26918 24506
rect 26970 24454 26982 24506
rect 27034 24454 27046 24506
rect 27098 24454 27110 24506
rect 27162 24454 27174 24506
rect 27226 24454 27238 24506
rect 27290 24454 28888 24506
rect 1104 24432 28888 24454
rect 5442 24216 5448 24268
rect 5500 24256 5506 24268
rect 5500 24228 7236 24256
rect 5500 24216 5506 24228
rect 1302 24148 1308 24200
rect 1360 24188 1366 24200
rect 1397 24191 1455 24197
rect 1397 24188 1409 24191
rect 1360 24160 1409 24188
rect 1360 24148 1366 24160
rect 1397 24157 1409 24160
rect 1443 24188 1455 24191
rect 1673 24191 1731 24197
rect 1673 24188 1685 24191
rect 1443 24160 1685 24188
rect 1443 24157 1455 24160
rect 1397 24151 1455 24157
rect 1673 24157 1685 24160
rect 1719 24157 1731 24191
rect 1673 24151 1731 24157
rect 6822 24148 6828 24200
rect 6880 24148 6886 24200
rect 7208 24197 7236 24228
rect 7193 24191 7251 24197
rect 7193 24157 7205 24191
rect 7239 24157 7251 24191
rect 7193 24151 7251 24157
rect 6914 24080 6920 24132
rect 6972 24120 6978 24132
rect 7009 24123 7067 24129
rect 7009 24120 7021 24123
rect 6972 24092 7021 24120
rect 6972 24080 6978 24092
rect 7009 24089 7021 24092
rect 7055 24089 7067 24123
rect 7009 24083 7067 24089
rect 7098 24080 7104 24132
rect 7156 24080 7162 24132
rect 1581 24055 1639 24061
rect 1581 24021 1593 24055
rect 1627 24052 1639 24055
rect 2038 24052 2044 24064
rect 1627 24024 2044 24052
rect 1627 24021 1639 24024
rect 1581 24015 1639 24021
rect 2038 24012 2044 24024
rect 2096 24012 2102 24064
rect 7377 24055 7435 24061
rect 7377 24021 7389 24055
rect 7423 24052 7435 24055
rect 8386 24052 8392 24064
rect 7423 24024 8392 24052
rect 7423 24021 7435 24024
rect 7377 24015 7435 24021
rect 8386 24012 8392 24024
rect 8444 24012 8450 24064
rect 1104 23962 28888 23984
rect 1104 23910 3658 23962
rect 3710 23910 3722 23962
rect 3774 23910 3786 23962
rect 3838 23910 3850 23962
rect 3902 23910 3914 23962
rect 3966 23910 3978 23962
rect 4030 23910 11658 23962
rect 11710 23910 11722 23962
rect 11774 23910 11786 23962
rect 11838 23910 11850 23962
rect 11902 23910 11914 23962
rect 11966 23910 11978 23962
rect 12030 23910 19658 23962
rect 19710 23910 19722 23962
rect 19774 23910 19786 23962
rect 19838 23910 19850 23962
rect 19902 23910 19914 23962
rect 19966 23910 19978 23962
rect 20030 23910 27658 23962
rect 27710 23910 27722 23962
rect 27774 23910 27786 23962
rect 27838 23910 27850 23962
rect 27902 23910 27914 23962
rect 27966 23910 27978 23962
rect 28030 23910 28888 23962
rect 1104 23888 28888 23910
rect 6822 23808 6828 23860
rect 6880 23848 6886 23860
rect 7285 23851 7343 23857
rect 7285 23848 7297 23851
rect 6880 23820 7297 23848
rect 6880 23808 6886 23820
rect 7285 23817 7297 23820
rect 7331 23817 7343 23851
rect 7285 23811 7343 23817
rect 7469 23851 7527 23857
rect 7469 23817 7481 23851
rect 7515 23848 7527 23851
rect 8021 23851 8079 23857
rect 8021 23848 8033 23851
rect 7515 23820 8033 23848
rect 7515 23817 7527 23820
rect 7469 23811 7527 23817
rect 8021 23817 8033 23820
rect 8067 23817 8079 23851
rect 8021 23811 8079 23817
rect 2884 23752 4476 23780
rect 1302 23672 1308 23724
rect 1360 23712 1366 23724
rect 1489 23715 1547 23721
rect 1489 23712 1501 23715
rect 1360 23684 1501 23712
rect 1360 23672 1366 23684
rect 1489 23681 1501 23684
rect 1535 23712 1547 23715
rect 1949 23715 2007 23721
rect 1949 23712 1961 23715
rect 1535 23684 1961 23712
rect 1535 23681 1547 23684
rect 1489 23675 1547 23681
rect 1949 23681 1961 23684
rect 1995 23681 2007 23715
rect 1949 23675 2007 23681
rect 2682 23672 2688 23724
rect 2740 23712 2746 23724
rect 2884 23721 2912 23752
rect 2869 23715 2927 23721
rect 2869 23712 2881 23715
rect 2740 23684 2881 23712
rect 2740 23672 2746 23684
rect 2869 23681 2881 23684
rect 2915 23681 2927 23715
rect 2869 23675 2927 23681
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23681 3019 23715
rect 2961 23675 3019 23681
rect 3237 23715 3295 23721
rect 3237 23681 3249 23715
rect 3283 23712 3295 23715
rect 3418 23712 3424 23724
rect 3283 23684 3424 23712
rect 3283 23681 3295 23684
rect 3237 23675 3295 23681
rect 2774 23604 2780 23656
rect 2832 23644 2838 23656
rect 2976 23644 3004 23675
rect 3418 23672 3424 23684
rect 3476 23672 3482 23724
rect 3513 23715 3571 23721
rect 3513 23681 3525 23715
rect 3559 23712 3571 23715
rect 3786 23712 3792 23724
rect 3559 23684 3792 23712
rect 3559 23681 3571 23684
rect 3513 23675 3571 23681
rect 3786 23672 3792 23684
rect 3844 23672 3850 23724
rect 4448 23721 4476 23752
rect 7944 23752 8616 23780
rect 7944 23724 7972 23752
rect 4433 23715 4491 23721
rect 4433 23681 4445 23715
rect 4479 23712 4491 23715
rect 5442 23712 5448 23724
rect 4479 23684 5448 23712
rect 4479 23681 4491 23684
rect 4433 23675 4491 23681
rect 5442 23672 5448 23684
rect 5500 23672 5506 23724
rect 6549 23715 6607 23721
rect 6549 23681 6561 23715
rect 6595 23681 6607 23715
rect 6549 23675 6607 23681
rect 2832 23616 3004 23644
rect 2832 23604 2838 23616
rect 3694 23604 3700 23656
rect 3752 23644 3758 23656
rect 6564 23644 6592 23675
rect 6914 23672 6920 23724
rect 6972 23712 6978 23724
rect 7288 23715 7346 23721
rect 7288 23712 7300 23715
rect 6972 23684 7300 23712
rect 6972 23672 6978 23684
rect 7288 23681 7300 23684
rect 7334 23681 7346 23715
rect 7288 23675 7346 23681
rect 7834 23672 7840 23724
rect 7892 23672 7898 23724
rect 7926 23672 7932 23724
rect 7984 23672 7990 23724
rect 8386 23672 8392 23724
rect 8444 23672 8450 23724
rect 8588 23721 8616 23752
rect 8573 23715 8631 23721
rect 8573 23681 8585 23715
rect 8619 23681 8631 23715
rect 8573 23675 8631 23681
rect 6730 23644 6736 23656
rect 3752 23616 6736 23644
rect 3752 23604 3758 23616
rect 6730 23604 6736 23616
rect 6788 23644 6794 23656
rect 6825 23647 6883 23653
rect 6825 23644 6837 23647
rect 6788 23616 6837 23644
rect 6788 23604 6794 23616
rect 6825 23613 6837 23616
rect 6871 23613 6883 23647
rect 6825 23607 6883 23613
rect 7650 23604 7656 23656
rect 7708 23644 7714 23656
rect 8297 23647 8355 23653
rect 8297 23644 8309 23647
rect 7708 23616 8309 23644
rect 7708 23604 7714 23616
rect 8297 23613 8309 23616
rect 8343 23613 8355 23647
rect 8297 23607 8355 23613
rect 1394 23536 1400 23588
rect 1452 23576 1458 23588
rect 1765 23579 1823 23585
rect 1765 23576 1777 23579
rect 1452 23548 1777 23576
rect 1452 23536 1458 23548
rect 1765 23545 1777 23548
rect 1811 23545 1823 23579
rect 1765 23539 1823 23545
rect 2498 23536 2504 23588
rect 2556 23576 2562 23588
rect 3145 23579 3203 23585
rect 3145 23576 3157 23579
rect 2556 23548 3157 23576
rect 2556 23536 2562 23548
rect 3145 23545 3157 23548
rect 3191 23576 3203 23579
rect 3191 23548 4200 23576
rect 3191 23545 3203 23548
rect 3145 23539 3203 23545
rect 1581 23511 1639 23517
rect 1581 23477 1593 23511
rect 1627 23508 1639 23511
rect 1946 23508 1952 23520
rect 1627 23480 1952 23508
rect 1627 23477 1639 23480
rect 1581 23471 1639 23477
rect 1946 23468 1952 23480
rect 2004 23468 2010 23520
rect 2590 23468 2596 23520
rect 2648 23508 2654 23520
rect 2685 23511 2743 23517
rect 2685 23508 2697 23511
rect 2648 23480 2697 23508
rect 2648 23468 2654 23480
rect 2685 23477 2697 23480
rect 2731 23477 2743 23511
rect 2685 23471 2743 23477
rect 3418 23468 3424 23520
rect 3476 23468 3482 23520
rect 4172 23508 4200 23548
rect 4246 23536 4252 23588
rect 4304 23576 4310 23588
rect 4341 23579 4399 23585
rect 4341 23576 4353 23579
rect 4304 23548 4353 23576
rect 4304 23536 4310 23548
rect 4341 23545 4353 23548
rect 4387 23576 4399 23579
rect 6917 23579 6975 23585
rect 6917 23576 6929 23579
rect 4387 23548 6929 23576
rect 4387 23545 4399 23548
rect 4341 23539 4399 23545
rect 6917 23545 6929 23548
rect 6963 23545 6975 23579
rect 6917 23539 6975 23545
rect 8205 23579 8263 23585
rect 8205 23545 8217 23579
rect 8251 23576 8263 23579
rect 9030 23576 9036 23588
rect 8251 23548 9036 23576
rect 8251 23545 8263 23548
rect 8205 23539 8263 23545
rect 9030 23536 9036 23548
rect 9088 23536 9094 23588
rect 5626 23508 5632 23520
rect 4172 23480 5632 23508
rect 5626 23468 5632 23480
rect 5684 23468 5690 23520
rect 6641 23511 6699 23517
rect 6641 23477 6653 23511
rect 6687 23508 6699 23511
rect 7098 23508 7104 23520
rect 6687 23480 7104 23508
rect 6687 23477 6699 23480
rect 6641 23471 6699 23477
rect 7098 23468 7104 23480
rect 7156 23508 7162 23520
rect 7742 23508 7748 23520
rect 7156 23480 7748 23508
rect 7156 23468 7162 23480
rect 7742 23468 7748 23480
rect 7800 23468 7806 23520
rect 8754 23468 8760 23520
rect 8812 23468 8818 23520
rect 1104 23418 28888 23440
rect 1104 23366 2918 23418
rect 2970 23366 2982 23418
rect 3034 23366 3046 23418
rect 3098 23366 3110 23418
rect 3162 23366 3174 23418
rect 3226 23366 3238 23418
rect 3290 23366 10918 23418
rect 10970 23366 10982 23418
rect 11034 23366 11046 23418
rect 11098 23366 11110 23418
rect 11162 23366 11174 23418
rect 11226 23366 11238 23418
rect 11290 23366 18918 23418
rect 18970 23366 18982 23418
rect 19034 23366 19046 23418
rect 19098 23366 19110 23418
rect 19162 23366 19174 23418
rect 19226 23366 19238 23418
rect 19290 23366 26918 23418
rect 26970 23366 26982 23418
rect 27034 23366 27046 23418
rect 27098 23366 27110 23418
rect 27162 23366 27174 23418
rect 27226 23366 27238 23418
rect 27290 23366 28888 23418
rect 1104 23344 28888 23366
rect 1762 23264 1768 23316
rect 1820 23304 1826 23316
rect 4706 23304 4712 23316
rect 1820 23276 4712 23304
rect 1820 23264 1826 23276
rect 2961 23239 3019 23245
rect 2961 23205 2973 23239
rect 3007 23236 3019 23239
rect 3326 23236 3332 23248
rect 3007 23208 3332 23236
rect 3007 23205 3019 23208
rect 2961 23199 3019 23205
rect 3326 23196 3332 23208
rect 3384 23196 3390 23248
rect 3418 23196 3424 23248
rect 3476 23196 3482 23248
rect 2498 23128 2504 23180
rect 2556 23168 2562 23180
rect 3436 23168 3464 23196
rect 2556 23140 2820 23168
rect 2556 23128 2562 23140
rect 1394 23060 1400 23112
rect 1452 23060 1458 23112
rect 1673 23103 1731 23109
rect 1673 23069 1685 23103
rect 1719 23100 1731 23103
rect 2314 23100 2320 23112
rect 1719 23072 2320 23100
rect 1719 23069 1731 23072
rect 1673 23063 1731 23069
rect 2314 23060 2320 23072
rect 2372 23060 2378 23112
rect 2406 23060 2412 23112
rect 2464 23060 2470 23112
rect 2590 23060 2596 23112
rect 2648 23060 2654 23112
rect 2792 23109 2820 23140
rect 3344 23140 3464 23168
rect 2777 23103 2835 23109
rect 2777 23069 2789 23103
rect 2823 23069 2835 23103
rect 2777 23063 2835 23069
rect 2866 23060 2872 23112
rect 2924 23100 2930 23112
rect 3344 23109 3372 23140
rect 3053 23103 3111 23109
rect 3053 23100 3065 23103
rect 2924 23072 3065 23100
rect 2924 23060 2930 23072
rect 3053 23069 3065 23072
rect 3099 23069 3111 23103
rect 3329 23103 3387 23109
rect 3329 23100 3341 23103
rect 3053 23063 3111 23069
rect 3160 23072 3341 23100
rect 2685 23035 2743 23041
rect 2685 23001 2697 23035
rect 2731 23032 2743 23035
rect 3160 23032 3188 23072
rect 3329 23069 3341 23072
rect 3375 23069 3387 23103
rect 3329 23063 3387 23069
rect 3421 23103 3479 23109
rect 3421 23069 3433 23103
rect 3467 23100 3479 23103
rect 3528 23100 3556 23276
rect 4706 23264 4712 23276
rect 4764 23264 4770 23316
rect 7377 23307 7435 23313
rect 7377 23273 7389 23307
rect 7423 23304 7435 23307
rect 7650 23304 7656 23316
rect 7423 23276 7656 23304
rect 7423 23273 7435 23276
rect 7377 23267 7435 23273
rect 7650 23264 7656 23276
rect 7708 23264 7714 23316
rect 7926 23264 7932 23316
rect 7984 23304 7990 23316
rect 8021 23307 8079 23313
rect 8021 23304 8033 23307
rect 7984 23276 8033 23304
rect 7984 23264 7990 23276
rect 8021 23273 8033 23276
rect 8067 23273 8079 23307
rect 8021 23267 8079 23273
rect 5626 23196 5632 23248
rect 5684 23236 5690 23248
rect 7561 23239 7619 23245
rect 7561 23236 7573 23239
rect 5684 23208 7573 23236
rect 5684 23196 5690 23208
rect 7561 23205 7573 23208
rect 7607 23205 7619 23239
rect 7561 23199 7619 23205
rect 4617 23171 4675 23177
rect 4617 23168 4629 23171
rect 3988 23140 4629 23168
rect 3467 23072 3556 23100
rect 3467 23069 3479 23072
rect 3421 23063 3479 23069
rect 3786 23060 3792 23112
rect 3844 23060 3850 23112
rect 3988 23109 4016 23140
rect 4617 23137 4629 23140
rect 4663 23168 4675 23171
rect 4663 23140 5396 23168
rect 4663 23137 4675 23140
rect 4617 23131 4675 23137
rect 3973 23103 4031 23109
rect 3973 23069 3985 23103
rect 4019 23069 4031 23103
rect 3973 23063 4031 23069
rect 4062 23060 4068 23112
rect 4120 23060 4126 23112
rect 4246 23060 4252 23112
rect 4304 23060 4310 23112
rect 4706 23060 4712 23112
rect 4764 23060 4770 23112
rect 2731 23004 3188 23032
rect 3237 23035 3295 23041
rect 2731 23001 2743 23004
rect 2685 22995 2743 23001
rect 3237 23001 3249 23035
rect 3283 23032 3295 23035
rect 3694 23032 3700 23044
rect 3283 23004 3700 23032
rect 3283 23001 3295 23004
rect 3237 22995 3295 23001
rect 2498 22924 2504 22976
rect 2556 22964 2562 22976
rect 3252 22964 3280 22995
rect 3694 22992 3700 23004
rect 3752 22992 3758 23044
rect 3881 23035 3939 23041
rect 3881 23001 3893 23035
rect 3927 23032 3939 23035
rect 3927 23004 4292 23032
rect 3927 23001 3939 23004
rect 3881 22995 3939 23001
rect 4264 22976 4292 23004
rect 2556 22936 3280 22964
rect 2556 22924 2562 22936
rect 3510 22924 3516 22976
rect 3568 22964 3574 22976
rect 3605 22967 3663 22973
rect 3605 22964 3617 22967
rect 3568 22936 3617 22964
rect 3568 22924 3574 22936
rect 3605 22933 3617 22936
rect 3651 22933 3663 22967
rect 3605 22927 3663 22933
rect 4154 22924 4160 22976
rect 4212 22924 4218 22976
rect 4246 22924 4252 22976
rect 4304 22924 4310 22976
rect 4724 22964 4752 23060
rect 5368 23032 5396 23140
rect 6362 23128 6368 23180
rect 6420 23168 6426 23180
rect 6914 23168 6920 23180
rect 6420 23140 6920 23168
rect 6420 23128 6426 23140
rect 6914 23128 6920 23140
rect 6972 23128 6978 23180
rect 7576 23168 7604 23199
rect 8110 23196 8116 23248
rect 8168 23196 8174 23248
rect 8205 23239 8263 23245
rect 8205 23205 8217 23239
rect 8251 23205 8263 23239
rect 8205 23199 8263 23205
rect 8220 23168 8248 23199
rect 8478 23168 8484 23180
rect 7576 23140 8484 23168
rect 8478 23128 8484 23140
rect 8536 23128 8542 23180
rect 6822 23060 6828 23112
rect 6880 23060 6886 23112
rect 7098 23060 7104 23112
rect 7156 23060 7162 23112
rect 7190 23060 7196 23112
rect 7248 23060 7254 23112
rect 7469 23103 7527 23109
rect 7469 23069 7481 23103
rect 7515 23069 7527 23103
rect 7469 23063 7527 23069
rect 7484 23032 7512 23063
rect 7742 23060 7748 23112
rect 7800 23060 7806 23112
rect 7837 23103 7895 23109
rect 7837 23069 7849 23103
rect 7883 23069 7895 23103
rect 7837 23063 7895 23069
rect 5368 23004 7512 23032
rect 7558 22992 7564 23044
rect 7616 23032 7622 23044
rect 7852 23032 7880 23063
rect 7616 23004 7880 23032
rect 8573 23035 8631 23041
rect 7616 22992 7622 23004
rect 8573 23001 8585 23035
rect 8619 23001 8631 23035
rect 8573 22995 8631 23001
rect 8588 22964 8616 22995
rect 8938 22964 8944 22976
rect 4724 22936 8944 22964
rect 8938 22924 8944 22936
rect 8996 22924 9002 22976
rect 1104 22874 28888 22896
rect 1104 22822 3658 22874
rect 3710 22822 3722 22874
rect 3774 22822 3786 22874
rect 3838 22822 3850 22874
rect 3902 22822 3914 22874
rect 3966 22822 3978 22874
rect 4030 22822 11658 22874
rect 11710 22822 11722 22874
rect 11774 22822 11786 22874
rect 11838 22822 11850 22874
rect 11902 22822 11914 22874
rect 11966 22822 11978 22874
rect 12030 22822 19658 22874
rect 19710 22822 19722 22874
rect 19774 22822 19786 22874
rect 19838 22822 19850 22874
rect 19902 22822 19914 22874
rect 19966 22822 19978 22874
rect 20030 22822 27658 22874
rect 27710 22822 27722 22874
rect 27774 22822 27786 22874
rect 27838 22822 27850 22874
rect 27902 22822 27914 22874
rect 27966 22822 27978 22874
rect 28030 22822 28888 22874
rect 1104 22800 28888 22822
rect 2866 22720 2872 22772
rect 2924 22760 2930 22772
rect 3418 22760 3424 22772
rect 2924 22732 3424 22760
rect 2924 22720 2930 22732
rect 3418 22720 3424 22732
rect 3476 22760 3482 22772
rect 3605 22763 3663 22769
rect 3605 22760 3617 22763
rect 3476 22732 3617 22760
rect 3476 22720 3482 22732
rect 3605 22729 3617 22732
rect 3651 22729 3663 22763
rect 3605 22723 3663 22729
rect 7098 22720 7104 22772
rect 7156 22760 7162 22772
rect 7466 22760 7472 22772
rect 7156 22732 7472 22760
rect 7156 22720 7162 22732
rect 7466 22720 7472 22732
rect 7524 22760 7530 22772
rect 7745 22763 7803 22769
rect 7745 22760 7757 22763
rect 7524 22732 7757 22760
rect 7524 22720 7530 22732
rect 7745 22729 7757 22732
rect 7791 22729 7803 22763
rect 7745 22723 7803 22729
rect 6178 22692 6184 22704
rect 2148 22664 6184 22692
rect 1210 22584 1216 22636
rect 1268 22624 1274 22636
rect 1489 22627 1547 22633
rect 1489 22624 1501 22627
rect 1268 22596 1501 22624
rect 1268 22584 1274 22596
rect 1489 22593 1501 22596
rect 1535 22624 1547 22627
rect 1765 22627 1823 22633
rect 1765 22624 1777 22627
rect 1535 22596 1777 22624
rect 1535 22593 1547 22596
rect 1489 22587 1547 22593
rect 1765 22593 1777 22596
rect 1811 22593 1823 22627
rect 1765 22587 1823 22593
rect 1946 22584 1952 22636
rect 2004 22624 2010 22636
rect 2148 22633 2176 22664
rect 6178 22652 6184 22664
rect 6236 22692 6242 22704
rect 7190 22692 7196 22704
rect 6236 22664 7196 22692
rect 6236 22652 6242 22664
rect 7190 22652 7196 22664
rect 7248 22652 7254 22704
rect 2133 22627 2191 22633
rect 2133 22624 2145 22627
rect 2004 22596 2145 22624
rect 2004 22584 2010 22596
rect 2133 22593 2145 22596
rect 2179 22593 2191 22627
rect 2133 22587 2191 22593
rect 2222 22584 2228 22636
rect 2280 22584 2286 22636
rect 2501 22627 2559 22633
rect 2501 22593 2513 22627
rect 2547 22624 2559 22627
rect 2682 22624 2688 22636
rect 2547 22596 2688 22624
rect 2547 22593 2559 22596
rect 2501 22587 2559 22593
rect 2682 22584 2688 22596
rect 2740 22584 2746 22636
rect 3697 22627 3755 22633
rect 3697 22593 3709 22627
rect 3743 22624 3755 22627
rect 3970 22624 3976 22636
rect 3743 22596 3976 22624
rect 3743 22593 3755 22596
rect 3697 22587 3755 22593
rect 3970 22584 3976 22596
rect 4028 22584 4034 22636
rect 7208 22624 7236 22652
rect 7653 22627 7711 22633
rect 7653 22624 7665 22627
rect 7208 22596 7665 22624
rect 7653 22593 7665 22596
rect 7699 22624 7711 22627
rect 7742 22624 7748 22636
rect 7699 22596 7748 22624
rect 7699 22593 7711 22596
rect 7653 22587 7711 22593
rect 7742 22584 7748 22596
rect 7800 22584 7806 22636
rect 7926 22584 7932 22636
rect 7984 22584 7990 22636
rect 28074 22584 28080 22636
rect 28132 22584 28138 22636
rect 2038 22516 2044 22568
rect 2096 22556 2102 22568
rect 2593 22559 2651 22565
rect 2593 22556 2605 22559
rect 2096 22528 2605 22556
rect 2096 22516 2102 22528
rect 2593 22525 2605 22528
rect 2639 22525 2651 22559
rect 2593 22519 2651 22525
rect 2869 22559 2927 22565
rect 2869 22525 2881 22559
rect 2915 22525 2927 22559
rect 2869 22519 2927 22525
rect 1949 22491 2007 22497
rect 1949 22457 1961 22491
rect 1995 22488 2007 22491
rect 2774 22488 2780 22500
rect 1995 22460 2780 22488
rect 1995 22457 2007 22460
rect 1949 22451 2007 22457
rect 2774 22448 2780 22460
rect 2832 22448 2838 22500
rect 1581 22423 1639 22429
rect 1581 22389 1593 22423
rect 1627 22420 1639 22423
rect 2038 22420 2044 22432
rect 1627 22392 2044 22420
rect 1627 22389 1639 22392
rect 1581 22383 1639 22389
rect 2038 22380 2044 22392
rect 2096 22380 2102 22432
rect 2409 22423 2467 22429
rect 2409 22389 2421 22423
rect 2455 22420 2467 22423
rect 2590 22420 2596 22432
rect 2455 22392 2596 22420
rect 2455 22389 2467 22392
rect 2409 22383 2467 22389
rect 2590 22380 2596 22392
rect 2648 22420 2654 22432
rect 2884 22420 2912 22519
rect 28350 22516 28356 22568
rect 28408 22516 28414 22568
rect 7834 22448 7840 22500
rect 7892 22488 7898 22500
rect 7929 22491 7987 22497
rect 7929 22488 7941 22491
rect 7892 22460 7941 22488
rect 7892 22448 7898 22460
rect 7929 22457 7941 22460
rect 7975 22457 7987 22491
rect 7929 22451 7987 22457
rect 6362 22420 6368 22432
rect 2648 22392 6368 22420
rect 2648 22380 2654 22392
rect 6362 22380 6368 22392
rect 6420 22380 6426 22432
rect 1104 22330 28888 22352
rect 1104 22278 2918 22330
rect 2970 22278 2982 22330
rect 3034 22278 3046 22330
rect 3098 22278 3110 22330
rect 3162 22278 3174 22330
rect 3226 22278 3238 22330
rect 3290 22278 10918 22330
rect 10970 22278 10982 22330
rect 11034 22278 11046 22330
rect 11098 22278 11110 22330
rect 11162 22278 11174 22330
rect 11226 22278 11238 22330
rect 11290 22278 18918 22330
rect 18970 22278 18982 22330
rect 19034 22278 19046 22330
rect 19098 22278 19110 22330
rect 19162 22278 19174 22330
rect 19226 22278 19238 22330
rect 19290 22278 26918 22330
rect 26970 22278 26982 22330
rect 27034 22278 27046 22330
rect 27098 22278 27110 22330
rect 27162 22278 27174 22330
rect 27226 22278 27238 22330
rect 27290 22278 28888 22330
rect 1104 22256 28888 22278
rect 2406 22176 2412 22228
rect 2464 22216 2470 22228
rect 2501 22219 2559 22225
rect 2501 22216 2513 22219
rect 2464 22188 2513 22216
rect 2464 22176 2470 22188
rect 2501 22185 2513 22188
rect 2547 22185 2559 22219
rect 2501 22179 2559 22185
rect 3234 22176 3240 22228
rect 3292 22216 3298 22228
rect 3418 22216 3424 22228
rect 3292 22188 3424 22216
rect 3292 22176 3298 22188
rect 3418 22176 3424 22188
rect 3476 22176 3482 22228
rect 5442 22176 5448 22228
rect 5500 22216 5506 22228
rect 5500 22188 6132 22216
rect 5500 22176 5506 22188
rect 6104 22148 6132 22188
rect 7926 22176 7932 22228
rect 7984 22216 7990 22228
rect 9033 22219 9091 22225
rect 9033 22216 9045 22219
rect 7984 22188 9045 22216
rect 7984 22176 7990 22188
rect 9033 22185 9045 22188
rect 9079 22185 9091 22219
rect 9033 22179 9091 22185
rect 7101 22151 7159 22157
rect 7101 22148 7113 22151
rect 6104 22120 7113 22148
rect 7101 22117 7113 22120
rect 7147 22148 7159 22151
rect 7558 22148 7564 22160
rect 7147 22120 7564 22148
rect 7147 22117 7159 22120
rect 7101 22111 7159 22117
rect 7558 22108 7564 22120
rect 7616 22108 7622 22160
rect 2774 22040 2780 22092
rect 2832 22080 2838 22092
rect 4154 22080 4160 22092
rect 2832 22052 2912 22080
rect 2832 22040 2838 22052
rect 2590 21972 2596 22024
rect 2648 22021 2654 22024
rect 2884 22021 2912 22052
rect 3160 22052 4160 22080
rect 3160 22021 3188 22052
rect 4154 22040 4160 22052
rect 4212 22040 4218 22092
rect 4890 22040 4896 22092
rect 4948 22080 4954 22092
rect 4948 22052 5580 22080
rect 4948 22040 4954 22052
rect 2648 22015 2697 22021
rect 2648 21981 2651 22015
rect 2685 21981 2697 22015
rect 2648 21975 2697 21981
rect 2869 22015 2927 22021
rect 2869 21981 2881 22015
rect 2915 21981 2927 22015
rect 2869 21975 2927 21981
rect 2997 22015 3055 22021
rect 2997 21981 3009 22015
rect 3043 21981 3055 22015
rect 2997 21975 3055 21981
rect 3145 22015 3203 22021
rect 3145 21981 3157 22015
rect 3191 21981 3203 22015
rect 3145 21975 3203 21981
rect 3973 22015 4031 22021
rect 3973 21981 3985 22015
rect 4019 22012 4031 22015
rect 4341 22015 4399 22021
rect 4019 21984 4292 22012
rect 4019 21981 4031 21984
rect 3973 21975 4031 21981
rect 2648 21972 2654 21975
rect 1210 21904 1216 21956
rect 1268 21944 1274 21956
rect 1489 21947 1547 21953
rect 1489 21944 1501 21947
rect 1268 21916 1501 21944
rect 1268 21904 1274 21916
rect 1489 21913 1501 21916
rect 1535 21944 1547 21947
rect 1765 21947 1823 21953
rect 1765 21944 1777 21947
rect 1535 21916 1777 21944
rect 1535 21913 1547 21916
rect 1489 21907 1547 21913
rect 1765 21913 1777 21916
rect 1811 21913 1823 21947
rect 1765 21907 1823 21913
rect 2774 21904 2780 21956
rect 2832 21904 2838 21956
rect 1581 21879 1639 21885
rect 1581 21845 1593 21879
rect 1627 21876 1639 21879
rect 1854 21876 1860 21888
rect 1627 21848 1860 21876
rect 1627 21845 1639 21848
rect 1581 21839 1639 21845
rect 1854 21836 1860 21848
rect 1912 21836 1918 21888
rect 2498 21836 2504 21888
rect 2556 21876 2562 21888
rect 3012 21876 3040 21975
rect 4062 21904 4068 21956
rect 4120 21904 4126 21956
rect 4157 21947 4215 21953
rect 4157 21913 4169 21947
rect 4203 21913 4215 21947
rect 4264 21944 4292 21984
rect 4341 21981 4353 22015
rect 4387 22012 4399 22015
rect 5261 22015 5319 22021
rect 5261 22012 5273 22015
rect 4387 21984 5273 22012
rect 4387 21981 4399 21984
rect 4341 21975 4399 21981
rect 5261 21981 5273 21984
rect 5307 21981 5319 22015
rect 5261 21975 5319 21981
rect 4890 21944 4896 21956
rect 4264 21916 4896 21944
rect 4157 21907 4215 21913
rect 2556 21848 3040 21876
rect 2556 21836 2562 21848
rect 3418 21836 3424 21888
rect 3476 21876 3482 21888
rect 3789 21879 3847 21885
rect 3789 21876 3801 21879
rect 3476 21848 3801 21876
rect 3476 21836 3482 21848
rect 3789 21845 3801 21848
rect 3835 21845 3847 21879
rect 3789 21839 3847 21845
rect 3970 21836 3976 21888
rect 4028 21876 4034 21888
rect 4172 21876 4200 21907
rect 4890 21904 4896 21916
rect 4948 21904 4954 21956
rect 4028 21848 4200 21876
rect 5276 21876 5304 21975
rect 5442 21972 5448 22024
rect 5500 21972 5506 22024
rect 5552 22021 5580 22052
rect 5718 22040 5724 22092
rect 5776 22080 5782 22092
rect 5776 22052 6868 22080
rect 5776 22040 5782 22052
rect 5537 22015 5595 22021
rect 5537 21981 5549 22015
rect 5583 21981 5595 22015
rect 5537 21975 5595 21981
rect 5626 21972 5632 22024
rect 5684 21972 5690 22024
rect 5902 21972 5908 22024
rect 5960 22012 5966 22024
rect 5997 22015 6055 22021
rect 5997 22012 6009 22015
rect 5960 21984 6009 22012
rect 5960 21972 5966 21984
rect 5997 21981 6009 21984
rect 6043 21981 6055 22015
rect 5997 21975 6055 21981
rect 6178 21972 6184 22024
rect 6236 21972 6242 22024
rect 6362 21972 6368 22024
rect 6420 22021 6426 22024
rect 6840 22021 6868 22052
rect 8754 22040 8760 22092
rect 8812 22080 8818 22092
rect 8941 22083 8999 22089
rect 8941 22080 8953 22083
rect 8812 22052 8953 22080
rect 8812 22040 8818 22052
rect 8941 22049 8953 22052
rect 8987 22049 8999 22083
rect 8941 22043 8999 22049
rect 6420 22015 6447 22021
rect 6435 21981 6447 22015
rect 6420 21975 6447 21981
rect 6825 22015 6883 22021
rect 6825 21981 6837 22015
rect 6871 21981 6883 22015
rect 6825 21975 6883 21981
rect 6420 21972 6426 21975
rect 6914 21972 6920 22024
rect 6972 21972 6978 22024
rect 7193 22015 7251 22021
rect 7193 21981 7205 22015
rect 7239 21981 7251 22015
rect 7193 21975 7251 21981
rect 5644 21916 5948 21944
rect 5350 21876 5356 21888
rect 5276 21848 5356 21876
rect 4028 21836 4034 21848
rect 5350 21836 5356 21848
rect 5408 21876 5414 21888
rect 5644 21876 5672 21916
rect 5408 21848 5672 21876
rect 5408 21836 5414 21848
rect 5810 21836 5816 21888
rect 5868 21836 5874 21888
rect 5920 21876 5948 21916
rect 6086 21904 6092 21956
rect 6144 21944 6150 21956
rect 6273 21947 6331 21953
rect 6273 21944 6285 21947
rect 6144 21916 6285 21944
rect 6144 21904 6150 21916
rect 6273 21913 6285 21916
rect 6319 21913 6331 21947
rect 7208 21944 7236 21975
rect 9030 21972 9036 22024
rect 9088 22012 9094 22024
rect 9404 22015 9462 22021
rect 9404 22012 9416 22015
rect 9088 21984 9416 22012
rect 9088 21972 9094 21984
rect 9404 21981 9416 21984
rect 9450 21981 9462 22015
rect 9404 21975 9462 21981
rect 6273 21907 6331 21913
rect 6380 21916 7236 21944
rect 6380 21876 6408 21916
rect 5920 21848 6408 21876
rect 6546 21836 6552 21888
rect 6604 21836 6610 21888
rect 6638 21836 6644 21888
rect 6696 21836 6702 21888
rect 8570 21836 8576 21888
rect 8628 21876 8634 21888
rect 9401 21879 9459 21885
rect 9401 21876 9413 21879
rect 8628 21848 9413 21876
rect 8628 21836 8634 21848
rect 9401 21845 9413 21848
rect 9447 21845 9459 21879
rect 9401 21839 9459 21845
rect 9490 21836 9496 21888
rect 9548 21876 9554 21888
rect 9585 21879 9643 21885
rect 9585 21876 9597 21879
rect 9548 21848 9597 21876
rect 9548 21836 9554 21848
rect 9585 21845 9597 21848
rect 9631 21845 9643 21879
rect 9585 21839 9643 21845
rect 1104 21786 28888 21808
rect 1104 21734 3658 21786
rect 3710 21734 3722 21786
rect 3774 21734 3786 21786
rect 3838 21734 3850 21786
rect 3902 21734 3914 21786
rect 3966 21734 3978 21786
rect 4030 21734 11658 21786
rect 11710 21734 11722 21786
rect 11774 21734 11786 21786
rect 11838 21734 11850 21786
rect 11902 21734 11914 21786
rect 11966 21734 11978 21786
rect 12030 21734 19658 21786
rect 19710 21734 19722 21786
rect 19774 21734 19786 21786
rect 19838 21734 19850 21786
rect 19902 21734 19914 21786
rect 19966 21734 19978 21786
rect 20030 21734 27658 21786
rect 27710 21734 27722 21786
rect 27774 21734 27786 21786
rect 27838 21734 27850 21786
rect 27902 21734 27914 21786
rect 27966 21734 27978 21786
rect 28030 21734 28888 21786
rect 1104 21712 28888 21734
rect 2130 21632 2136 21684
rect 2188 21672 2194 21684
rect 2188 21644 4844 21672
rect 2188 21632 2194 21644
rect 3234 21604 3240 21616
rect 2424 21576 3240 21604
rect 1302 21496 1308 21548
rect 1360 21536 1366 21548
rect 2424 21545 2452 21576
rect 3234 21564 3240 21576
rect 3292 21564 3298 21616
rect 4816 21604 4844 21644
rect 4890 21632 4896 21684
rect 4948 21632 4954 21684
rect 6086 21632 6092 21684
rect 6144 21672 6150 21684
rect 6914 21672 6920 21684
rect 6144 21644 6920 21672
rect 6144 21632 6150 21644
rect 6914 21632 6920 21644
rect 6972 21632 6978 21684
rect 5718 21604 5724 21616
rect 4816 21576 5724 21604
rect 5718 21564 5724 21576
rect 5776 21564 5782 21616
rect 5810 21564 5816 21616
rect 5868 21604 5874 21616
rect 5905 21607 5963 21613
rect 5905 21604 5917 21607
rect 5868 21576 5917 21604
rect 5868 21564 5874 21576
rect 5905 21573 5917 21576
rect 5951 21604 5963 21607
rect 5951 21576 7052 21604
rect 5951 21573 5963 21576
rect 5905 21567 5963 21573
rect 1397 21539 1455 21545
rect 1397 21536 1409 21539
rect 1360 21508 1409 21536
rect 1360 21496 1366 21508
rect 1397 21505 1409 21508
rect 1443 21536 1455 21539
rect 1857 21539 1915 21545
rect 1857 21536 1869 21539
rect 1443 21508 1869 21536
rect 1443 21505 1455 21508
rect 1397 21499 1455 21505
rect 1857 21505 1869 21508
rect 1903 21505 1915 21539
rect 1857 21499 1915 21505
rect 2409 21539 2467 21545
rect 2409 21505 2421 21539
rect 2455 21505 2467 21539
rect 2409 21499 2467 21505
rect 2682 21496 2688 21548
rect 2740 21496 2746 21548
rect 2777 21539 2835 21545
rect 2777 21505 2789 21539
rect 2823 21505 2835 21539
rect 2777 21499 2835 21505
rect 2590 21428 2596 21480
rect 2648 21468 2654 21480
rect 2792 21468 2820 21499
rect 3602 21496 3608 21548
rect 3660 21536 3666 21548
rect 4985 21539 5043 21545
rect 4985 21536 4997 21539
rect 3660 21508 4997 21536
rect 3660 21496 3666 21508
rect 4985 21505 4997 21508
rect 5031 21505 5043 21539
rect 4985 21499 5043 21505
rect 6089 21539 6147 21545
rect 6089 21505 6101 21539
rect 6135 21505 6147 21539
rect 6089 21499 6147 21505
rect 6181 21539 6239 21545
rect 6181 21505 6193 21539
rect 6227 21536 6239 21539
rect 6454 21536 6460 21548
rect 6227 21508 6460 21536
rect 6227 21505 6239 21508
rect 6181 21499 6239 21505
rect 2648 21440 2820 21468
rect 2648 21428 2654 21440
rect 1210 21360 1216 21412
rect 1268 21400 1274 21412
rect 1673 21403 1731 21409
rect 1673 21400 1685 21403
rect 1268 21372 1685 21400
rect 1268 21360 1274 21372
rect 1673 21369 1685 21372
rect 1719 21369 1731 21403
rect 1673 21363 1731 21369
rect 1578 21292 1584 21344
rect 1636 21292 1642 21344
rect 2406 21292 2412 21344
rect 2464 21332 2470 21344
rect 2501 21335 2559 21341
rect 2501 21332 2513 21335
rect 2464 21304 2513 21332
rect 2464 21292 2470 21304
rect 2501 21301 2513 21304
rect 2547 21301 2559 21335
rect 2501 21295 2559 21301
rect 2774 21292 2780 21344
rect 2832 21332 2838 21344
rect 2961 21335 3019 21341
rect 2961 21332 2973 21335
rect 2832 21304 2973 21332
rect 2832 21292 2838 21304
rect 2961 21301 2973 21304
rect 3007 21301 3019 21335
rect 2961 21295 3019 21301
rect 5902 21292 5908 21344
rect 5960 21292 5966 21344
rect 6104 21332 6132 21499
rect 6454 21496 6460 21508
rect 6512 21536 6518 21548
rect 7024 21545 7052 21576
rect 8478 21564 8484 21616
rect 8536 21564 8542 21616
rect 6549 21539 6607 21545
rect 6549 21536 6561 21539
rect 6512 21508 6561 21536
rect 6512 21496 6518 21508
rect 6549 21505 6561 21508
rect 6595 21505 6607 21539
rect 6549 21499 6607 21505
rect 6641 21539 6699 21545
rect 6641 21505 6653 21539
rect 6687 21505 6699 21539
rect 6641 21499 6699 21505
rect 7009 21539 7067 21545
rect 7009 21505 7021 21539
rect 7055 21505 7067 21539
rect 7009 21499 7067 21505
rect 7469 21539 7527 21545
rect 7469 21505 7481 21539
rect 7515 21505 7527 21539
rect 7469 21499 7527 21505
rect 6656 21468 6684 21499
rect 7285 21471 7343 21477
rect 7285 21468 7297 21471
rect 6656 21440 7297 21468
rect 7285 21437 7297 21440
rect 7331 21437 7343 21471
rect 7285 21431 7343 21437
rect 7484 21468 7512 21499
rect 7742 21496 7748 21548
rect 7800 21496 7806 21548
rect 7926 21496 7932 21548
rect 7984 21496 7990 21548
rect 8021 21471 8079 21477
rect 8021 21468 8033 21471
rect 7484 21440 8033 21468
rect 7006 21360 7012 21412
rect 7064 21400 7070 21412
rect 7484 21400 7512 21440
rect 8021 21437 8033 21440
rect 8067 21437 8079 21471
rect 8021 21431 8079 21437
rect 7064 21372 7512 21400
rect 8205 21403 8263 21409
rect 7064 21360 7070 21372
rect 8205 21369 8217 21403
rect 8251 21400 8263 21403
rect 8294 21400 8300 21412
rect 8251 21372 8300 21400
rect 8251 21369 8263 21372
rect 8205 21363 8263 21369
rect 8294 21360 8300 21372
rect 8352 21360 8358 21412
rect 6546 21332 6552 21344
rect 6104 21304 6552 21332
rect 6546 21292 6552 21304
rect 6604 21332 6610 21344
rect 6917 21335 6975 21341
rect 6917 21332 6929 21335
rect 6604 21304 6929 21332
rect 6604 21292 6610 21304
rect 6917 21301 6929 21304
rect 6963 21301 6975 21335
rect 6917 21295 6975 21301
rect 7190 21292 7196 21344
rect 7248 21292 7254 21344
rect 1104 21242 28888 21264
rect 1104 21190 2918 21242
rect 2970 21190 2982 21242
rect 3034 21190 3046 21242
rect 3098 21190 3110 21242
rect 3162 21190 3174 21242
rect 3226 21190 3238 21242
rect 3290 21190 10918 21242
rect 10970 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 11238 21242
rect 11290 21190 18918 21242
rect 18970 21190 18982 21242
rect 19034 21190 19046 21242
rect 19098 21190 19110 21242
rect 19162 21190 19174 21242
rect 19226 21190 19238 21242
rect 19290 21190 26918 21242
rect 26970 21190 26982 21242
rect 27034 21190 27046 21242
rect 27098 21190 27110 21242
rect 27162 21190 27174 21242
rect 27226 21190 27238 21242
rect 27290 21190 28888 21242
rect 1104 21168 28888 21190
rect 2746 21100 3372 21128
rect 2746 21060 2774 21100
rect 1688 21032 2774 21060
rect 3344 21060 3372 21100
rect 3510 21088 3516 21140
rect 3568 21128 3574 21140
rect 3881 21131 3939 21137
rect 3881 21128 3893 21131
rect 3568 21100 3893 21128
rect 3568 21088 3574 21100
rect 3881 21097 3893 21100
rect 3927 21097 3939 21131
rect 3881 21091 3939 21097
rect 5350 21088 5356 21140
rect 5408 21088 5414 21140
rect 5902 21088 5908 21140
rect 5960 21128 5966 21140
rect 7101 21131 7159 21137
rect 7101 21128 7113 21131
rect 5960 21100 7113 21128
rect 5960 21088 5966 21100
rect 7101 21097 7113 21100
rect 7147 21097 7159 21131
rect 7101 21091 7159 21097
rect 8294 21060 8300 21072
rect 3344 21032 8300 21060
rect 1688 21001 1716 21032
rect 3528 21004 3556 21032
rect 8294 21020 8300 21032
rect 8352 21020 8358 21072
rect 8938 21020 8944 21072
rect 8996 21060 9002 21072
rect 8996 21032 9536 21060
rect 8996 21020 9002 21032
rect 1673 20995 1731 21001
rect 1673 20961 1685 20995
rect 1719 20961 1731 20995
rect 1673 20955 1731 20961
rect 2774 20952 2780 21004
rect 2832 20992 2838 21004
rect 2832 20964 3188 20992
rect 2832 20952 2838 20964
rect 1302 20884 1308 20936
rect 1360 20924 1366 20936
rect 1397 20927 1455 20933
rect 1397 20924 1409 20927
rect 1360 20896 1409 20924
rect 1360 20884 1366 20896
rect 1397 20893 1409 20896
rect 1443 20893 1455 20927
rect 1397 20887 1455 20893
rect 2869 20927 2927 20933
rect 2869 20893 2881 20927
rect 2915 20893 2927 20927
rect 2869 20887 2927 20893
rect 1946 20816 1952 20868
rect 2004 20856 2010 20868
rect 2774 20856 2780 20868
rect 2004 20828 2780 20856
rect 2004 20816 2010 20828
rect 2774 20816 2780 20828
rect 2832 20816 2838 20868
rect 2884 20856 2912 20887
rect 2958 20884 2964 20936
rect 3016 20884 3022 20936
rect 3160 20933 3188 20964
rect 3510 20952 3516 21004
rect 3568 20952 3574 21004
rect 8312 20992 8340 21020
rect 9122 20992 9128 21004
rect 8312 20964 9128 20992
rect 9122 20952 9128 20964
rect 9180 20992 9186 21004
rect 9180 20964 9444 20992
rect 9180 20952 9186 20964
rect 3145 20927 3203 20933
rect 3145 20893 3157 20927
rect 3191 20893 3203 20927
rect 3145 20887 3203 20893
rect 3329 20927 3387 20933
rect 3329 20893 3341 20927
rect 3375 20924 3387 20927
rect 3789 20927 3847 20933
rect 3789 20924 3801 20927
rect 3375 20896 3801 20924
rect 3375 20893 3387 20896
rect 3329 20887 3387 20893
rect 3789 20893 3801 20896
rect 3835 20893 3847 20927
rect 3789 20887 3847 20893
rect 4246 20884 4252 20936
rect 4304 20884 4310 20936
rect 5442 20884 5448 20936
rect 5500 20884 5506 20936
rect 7006 20884 7012 20936
rect 7064 20884 7070 20936
rect 7190 20884 7196 20936
rect 7248 20924 7254 20936
rect 7285 20927 7343 20933
rect 7285 20924 7297 20927
rect 7248 20896 7297 20924
rect 7248 20884 7254 20896
rect 7285 20893 7297 20896
rect 7331 20893 7343 20927
rect 7285 20887 7343 20893
rect 7374 20884 7380 20936
rect 7432 20884 7438 20936
rect 9416 20933 9444 20964
rect 9508 20933 9536 21032
rect 9401 20927 9459 20933
rect 9401 20893 9413 20927
rect 9447 20893 9459 20927
rect 9401 20887 9459 20893
rect 9494 20927 9552 20933
rect 9494 20893 9506 20927
rect 9540 20893 9552 20927
rect 9494 20887 9552 20893
rect 3050 20856 3056 20868
rect 2884 20828 3056 20856
rect 3050 20816 3056 20828
rect 3108 20816 3114 20868
rect 7561 20859 7619 20865
rect 7561 20825 7573 20859
rect 7607 20856 7619 20859
rect 12894 20856 12900 20868
rect 7607 20828 12900 20856
rect 7607 20825 7619 20828
rect 7561 20819 7619 20825
rect 12894 20816 12900 20828
rect 12952 20816 12958 20868
rect 3326 20748 3332 20800
rect 3384 20788 3390 20800
rect 4065 20791 4123 20797
rect 4065 20788 4077 20791
rect 3384 20760 4077 20788
rect 3384 20748 3390 20760
rect 4065 20757 4077 20760
rect 4111 20757 4123 20791
rect 4065 20751 4123 20757
rect 4154 20748 4160 20800
rect 4212 20748 4218 20800
rect 4522 20748 4528 20800
rect 4580 20748 4586 20800
rect 9769 20791 9827 20797
rect 9769 20757 9781 20791
rect 9815 20788 9827 20791
rect 9858 20788 9864 20800
rect 9815 20760 9864 20788
rect 9815 20757 9827 20760
rect 9769 20751 9827 20757
rect 9858 20748 9864 20760
rect 9916 20748 9922 20800
rect 1104 20698 28888 20720
rect 1104 20646 3658 20698
rect 3710 20646 3722 20698
rect 3774 20646 3786 20698
rect 3838 20646 3850 20698
rect 3902 20646 3914 20698
rect 3966 20646 3978 20698
rect 4030 20646 11658 20698
rect 11710 20646 11722 20698
rect 11774 20646 11786 20698
rect 11838 20646 11850 20698
rect 11902 20646 11914 20698
rect 11966 20646 11978 20698
rect 12030 20646 19658 20698
rect 19710 20646 19722 20698
rect 19774 20646 19786 20698
rect 19838 20646 19850 20698
rect 19902 20646 19914 20698
rect 19966 20646 19978 20698
rect 20030 20646 27658 20698
rect 27710 20646 27722 20698
rect 27774 20646 27786 20698
rect 27838 20646 27850 20698
rect 27902 20646 27914 20698
rect 27966 20646 27978 20698
rect 28030 20646 28888 20698
rect 1104 20624 28888 20646
rect 3050 20544 3056 20596
rect 3108 20584 3114 20596
rect 3145 20587 3203 20593
rect 3145 20584 3157 20587
rect 3108 20556 3157 20584
rect 3108 20544 3114 20556
rect 3145 20553 3157 20556
rect 3191 20553 3203 20587
rect 3145 20547 3203 20553
rect 2777 20519 2835 20525
rect 2777 20485 2789 20519
rect 2823 20516 2835 20519
rect 4246 20516 4252 20528
rect 2823 20488 4252 20516
rect 2823 20485 2835 20488
rect 2777 20479 2835 20485
rect 4246 20476 4252 20488
rect 4304 20476 4310 20528
rect 5442 20476 5448 20528
rect 5500 20516 5506 20528
rect 5500 20488 9674 20516
rect 5500 20476 5506 20488
rect 1302 20408 1308 20460
rect 1360 20448 1366 20460
rect 1397 20451 1455 20457
rect 1397 20448 1409 20451
rect 1360 20420 1409 20448
rect 1360 20408 1366 20420
rect 1397 20417 1409 20420
rect 1443 20448 1455 20451
rect 1673 20451 1731 20457
rect 1673 20448 1685 20451
rect 1443 20420 1685 20448
rect 1443 20417 1455 20420
rect 1397 20411 1455 20417
rect 1673 20417 1685 20420
rect 1719 20417 1731 20451
rect 1673 20411 1731 20417
rect 2222 20408 2228 20460
rect 2280 20448 2286 20460
rect 2593 20451 2651 20457
rect 2593 20448 2605 20451
rect 2280 20420 2605 20448
rect 2280 20408 2286 20420
rect 2593 20417 2605 20420
rect 2639 20417 2651 20451
rect 2593 20411 2651 20417
rect 2682 20408 2688 20460
rect 2740 20448 2746 20460
rect 2869 20451 2927 20457
rect 2869 20448 2881 20451
rect 2740 20420 2881 20448
rect 2740 20408 2746 20420
rect 2869 20417 2881 20420
rect 2915 20417 2927 20451
rect 2869 20411 2927 20417
rect 2961 20451 3019 20457
rect 2961 20417 2973 20451
rect 3007 20417 3019 20451
rect 2961 20411 3019 20417
rect 2976 20380 3004 20411
rect 8938 20408 8944 20460
rect 8996 20448 9002 20460
rect 9033 20451 9091 20457
rect 9033 20448 9045 20451
rect 8996 20420 9045 20448
rect 8996 20408 9002 20420
rect 9033 20417 9045 20420
rect 9079 20417 9091 20451
rect 9033 20411 9091 20417
rect 9122 20408 9128 20460
rect 9180 20448 9186 20460
rect 9646 20457 9674 20488
rect 9493 20451 9551 20457
rect 9180 20420 9225 20448
rect 9180 20408 9186 20420
rect 9493 20417 9505 20451
rect 9539 20417 9551 20451
rect 9493 20411 9551 20417
rect 9631 20451 9689 20457
rect 9631 20417 9643 20451
rect 9677 20448 9689 20451
rect 9953 20451 10011 20457
rect 9953 20448 9965 20451
rect 9677 20420 9965 20448
rect 9677 20417 9689 20420
rect 9631 20411 9689 20417
rect 9953 20417 9965 20420
rect 9999 20417 10011 20451
rect 9953 20411 10011 20417
rect 10046 20451 10104 20457
rect 10046 20417 10058 20451
rect 10092 20417 10104 20451
rect 10046 20411 10104 20417
rect 1688 20352 3004 20380
rect 1688 20324 1716 20352
rect 2608 20324 2636 20352
rect 6730 20340 6736 20392
rect 6788 20380 6794 20392
rect 9508 20380 9536 20411
rect 10060 20380 10088 20411
rect 6788 20352 10088 20380
rect 6788 20340 6794 20352
rect 1670 20272 1676 20324
rect 1728 20272 1734 20324
rect 2590 20272 2596 20324
rect 2648 20272 2654 20324
rect 9401 20315 9459 20321
rect 9401 20281 9413 20315
rect 9447 20312 9459 20315
rect 9582 20312 9588 20324
rect 9447 20284 9588 20312
rect 9447 20281 9459 20284
rect 9401 20275 9459 20281
rect 9582 20272 9588 20284
rect 9640 20272 9646 20324
rect 9861 20315 9919 20321
rect 9861 20281 9873 20315
rect 9907 20312 9919 20315
rect 10042 20312 10048 20324
rect 9907 20284 10048 20312
rect 9907 20281 9919 20284
rect 9861 20275 9919 20281
rect 10042 20272 10048 20284
rect 10100 20272 10106 20324
rect 1581 20247 1639 20253
rect 1581 20213 1593 20247
rect 1627 20244 1639 20247
rect 3326 20244 3332 20256
rect 1627 20216 3332 20244
rect 1627 20213 1639 20216
rect 1581 20207 1639 20213
rect 3326 20204 3332 20216
rect 3384 20244 3390 20256
rect 5442 20244 5448 20256
rect 3384 20216 5448 20244
rect 3384 20204 3390 20216
rect 5442 20204 5448 20216
rect 5500 20204 5506 20256
rect 10137 20247 10195 20253
rect 10137 20213 10149 20247
rect 10183 20244 10195 20247
rect 10226 20244 10232 20256
rect 10183 20216 10232 20244
rect 10183 20213 10195 20216
rect 10137 20207 10195 20213
rect 10226 20204 10232 20216
rect 10284 20204 10290 20256
rect 21910 20204 21916 20256
rect 21968 20244 21974 20256
rect 24026 20244 24032 20256
rect 21968 20216 24032 20244
rect 21968 20204 21974 20216
rect 24026 20204 24032 20216
rect 24084 20204 24090 20256
rect 1104 20154 28888 20176
rect 1104 20102 2918 20154
rect 2970 20102 2982 20154
rect 3034 20102 3046 20154
rect 3098 20102 3110 20154
rect 3162 20102 3174 20154
rect 3226 20102 3238 20154
rect 3290 20102 10918 20154
rect 10970 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 11238 20154
rect 11290 20102 18918 20154
rect 18970 20102 18982 20154
rect 19034 20102 19046 20154
rect 19098 20102 19110 20154
rect 19162 20102 19174 20154
rect 19226 20102 19238 20154
rect 19290 20102 26918 20154
rect 26970 20102 26982 20154
rect 27034 20102 27046 20154
rect 27098 20102 27110 20154
rect 27162 20102 27174 20154
rect 27226 20102 27238 20154
rect 27290 20102 28888 20154
rect 1104 20080 28888 20102
rect 6457 20043 6515 20049
rect 6457 20009 6469 20043
rect 6503 20040 6515 20043
rect 6822 20040 6828 20052
rect 6503 20012 6828 20040
rect 6503 20009 6515 20012
rect 6457 20003 6515 20009
rect 6822 20000 6828 20012
rect 6880 20000 6886 20052
rect 7466 20000 7472 20052
rect 7524 20000 7530 20052
rect 9125 20043 9183 20049
rect 9125 20009 9137 20043
rect 9171 20040 9183 20043
rect 10134 20040 10140 20052
rect 9171 20012 10140 20040
rect 9171 20009 9183 20012
rect 9125 20003 9183 20009
rect 10134 20000 10140 20012
rect 10192 20000 10198 20052
rect 20796 20043 20854 20049
rect 20796 20009 20808 20043
rect 20842 20040 20854 20043
rect 22373 20043 22431 20049
rect 22373 20040 22385 20043
rect 20842 20012 22385 20040
rect 20842 20009 20854 20012
rect 20796 20003 20854 20009
rect 22373 20009 22385 20012
rect 22419 20009 22431 20043
rect 22373 20003 22431 20009
rect 23198 20000 23204 20052
rect 23256 20040 23262 20052
rect 23566 20040 23572 20052
rect 23256 20012 23572 20040
rect 23256 20000 23262 20012
rect 23566 20000 23572 20012
rect 23624 20000 23630 20052
rect 26145 20043 26203 20049
rect 26145 20009 26157 20043
rect 26191 20040 26203 20043
rect 28074 20040 28080 20052
rect 26191 20012 28080 20040
rect 26191 20009 26203 20012
rect 26145 20003 26203 20009
rect 28074 20000 28080 20012
rect 28132 20000 28138 20052
rect 3145 19975 3203 19981
rect 3145 19941 3157 19975
rect 3191 19972 3203 19975
rect 3510 19972 3516 19984
rect 3191 19944 3516 19972
rect 3191 19941 3203 19944
rect 3145 19935 3203 19941
rect 3510 19932 3516 19944
rect 3568 19932 3574 19984
rect 4522 19932 4528 19984
rect 4580 19972 4586 19984
rect 4580 19944 13124 19972
rect 4580 19932 4586 19944
rect 5810 19864 5816 19916
rect 5868 19904 5874 19916
rect 8018 19904 8024 19916
rect 5868 19876 8024 19904
rect 5868 19864 5874 19876
rect 1302 19796 1308 19848
rect 1360 19836 1366 19848
rect 1397 19839 1455 19845
rect 1397 19836 1409 19839
rect 1360 19808 1409 19836
rect 1360 19796 1366 19808
rect 1397 19805 1409 19808
rect 1443 19836 1455 19839
rect 1673 19839 1731 19845
rect 1673 19836 1685 19839
rect 1443 19808 1685 19836
rect 1443 19805 1455 19808
rect 1397 19799 1455 19805
rect 1673 19805 1685 19808
rect 1719 19805 1731 19839
rect 1673 19799 1731 19805
rect 2590 19796 2596 19848
rect 2648 19836 2654 19848
rect 5994 19836 6000 19848
rect 2648 19808 6000 19836
rect 2648 19796 2654 19808
rect 5994 19796 6000 19808
rect 6052 19836 6058 19848
rect 7392 19845 7420 19876
rect 8018 19864 8024 19876
rect 8076 19864 8082 19916
rect 8202 19864 8208 19916
rect 8260 19904 8266 19916
rect 8260 19876 9536 19904
rect 8260 19864 8266 19876
rect 9508 19845 9536 19876
rect 9858 19864 9864 19916
rect 9916 19904 9922 19916
rect 10413 19907 10471 19913
rect 10413 19904 10425 19907
rect 9916 19876 10425 19904
rect 9916 19864 9922 19876
rect 10413 19873 10425 19876
rect 10459 19873 10471 19907
rect 10413 19867 10471 19873
rect 12345 19907 12403 19913
rect 12345 19873 12357 19907
rect 12391 19904 12403 19907
rect 12434 19904 12440 19916
rect 12391 19876 12440 19904
rect 12391 19873 12403 19876
rect 12345 19867 12403 19873
rect 12434 19864 12440 19876
rect 12492 19864 12498 19916
rect 13096 19913 13124 19944
rect 22388 19944 23060 19972
rect 13081 19907 13139 19913
rect 13081 19873 13093 19907
rect 13127 19873 13139 19907
rect 13081 19867 13139 19873
rect 18785 19907 18843 19913
rect 18785 19873 18797 19907
rect 18831 19904 18843 19907
rect 20533 19907 20591 19913
rect 18831 19876 20392 19904
rect 18831 19873 18843 19876
rect 18785 19867 18843 19873
rect 6365 19839 6423 19845
rect 6365 19836 6377 19839
rect 6052 19808 6377 19836
rect 6052 19796 6058 19808
rect 6365 19805 6377 19808
rect 6411 19805 6423 19839
rect 6365 19799 6423 19805
rect 7377 19839 7435 19845
rect 7377 19805 7389 19839
rect 7423 19805 7435 19839
rect 9309 19839 9367 19845
rect 9309 19836 9321 19839
rect 7377 19799 7435 19805
rect 7484 19808 9321 19836
rect 1946 19728 1952 19780
rect 2004 19768 2010 19780
rect 2777 19771 2835 19777
rect 2777 19768 2789 19771
rect 2004 19740 2789 19768
rect 2004 19728 2010 19740
rect 2777 19737 2789 19740
rect 2823 19768 2835 19771
rect 4062 19768 4068 19780
rect 2823 19740 4068 19768
rect 2823 19737 2835 19740
rect 2777 19731 2835 19737
rect 4062 19728 4068 19740
rect 4120 19728 4126 19780
rect 6178 19728 6184 19780
rect 6236 19768 6242 19780
rect 7484 19768 7512 19808
rect 9309 19805 9321 19808
rect 9355 19805 9367 19839
rect 9309 19799 9367 19805
rect 9493 19839 9551 19845
rect 9493 19805 9505 19839
rect 9539 19805 9551 19839
rect 9493 19799 9551 19805
rect 9766 19796 9772 19848
rect 9824 19796 9830 19848
rect 10042 19796 10048 19848
rect 10100 19796 10106 19848
rect 10226 19796 10232 19848
rect 10284 19796 10290 19848
rect 13265 19839 13323 19845
rect 13265 19805 13277 19839
rect 13311 19836 13323 19839
rect 14458 19836 14464 19848
rect 13311 19808 14464 19836
rect 13311 19805 13323 19808
rect 13265 19799 13323 19805
rect 14458 19796 14464 19808
rect 14516 19796 14522 19848
rect 6236 19740 7512 19768
rect 6236 19728 6242 19740
rect 9398 19728 9404 19780
rect 9456 19728 9462 19780
rect 9582 19728 9588 19780
rect 9640 19777 9646 19780
rect 9640 19771 9669 19777
rect 9657 19768 9669 19771
rect 10137 19771 10195 19777
rect 10137 19768 10149 19771
rect 9657 19740 10149 19768
rect 9657 19737 9669 19740
rect 9640 19731 9669 19737
rect 10137 19737 10149 19740
rect 10183 19737 10195 19771
rect 10137 19731 10195 19737
rect 12437 19771 12495 19777
rect 12437 19737 12449 19771
rect 12483 19768 12495 19771
rect 12618 19768 12624 19780
rect 12483 19740 12624 19768
rect 12483 19737 12495 19740
rect 12437 19731 12495 19737
rect 9640 19728 9646 19731
rect 12618 19728 12624 19740
rect 12676 19728 12682 19780
rect 13357 19771 13415 19777
rect 13357 19768 13369 19771
rect 12912 19740 13369 19768
rect 1581 19703 1639 19709
rect 1581 19669 1593 19703
rect 1627 19700 1639 19703
rect 3050 19700 3056 19712
rect 1627 19672 3056 19700
rect 1627 19669 1639 19672
rect 1581 19663 1639 19669
rect 3050 19660 3056 19672
rect 3108 19660 3114 19712
rect 3237 19703 3295 19709
rect 3237 19669 3249 19703
rect 3283 19700 3295 19703
rect 3510 19700 3516 19712
rect 3283 19672 3516 19700
rect 3283 19669 3295 19672
rect 3237 19663 3295 19669
rect 3510 19660 3516 19672
rect 3568 19660 3574 19712
rect 9416 19700 9444 19728
rect 9861 19703 9919 19709
rect 9861 19700 9873 19703
rect 9416 19672 9873 19700
rect 9861 19669 9873 19672
rect 9907 19669 9919 19703
rect 9861 19663 9919 19669
rect 12526 19660 12532 19712
rect 12584 19660 12590 19712
rect 12912 19709 12940 19740
rect 13357 19737 13369 19740
rect 13403 19737 13415 19771
rect 18601 19771 18659 19777
rect 18601 19768 18613 19771
rect 13357 19731 13415 19737
rect 13740 19740 18613 19768
rect 13740 19709 13768 19740
rect 18601 19737 18613 19740
rect 18647 19737 18659 19771
rect 18601 19731 18659 19737
rect 12897 19703 12955 19709
rect 12897 19669 12909 19703
rect 12943 19669 12955 19703
rect 12897 19663 12955 19669
rect 13725 19703 13783 19709
rect 13725 19669 13737 19703
rect 13771 19669 13783 19703
rect 13725 19663 13783 19669
rect 18138 19660 18144 19712
rect 18196 19660 18202 19712
rect 18509 19703 18567 19709
rect 18509 19669 18521 19703
rect 18555 19700 18567 19703
rect 19061 19703 19119 19709
rect 19061 19700 19073 19703
rect 18555 19672 19073 19700
rect 18555 19669 18567 19672
rect 18509 19663 18567 19669
rect 19061 19669 19073 19672
rect 19107 19700 19119 19703
rect 19334 19700 19340 19712
rect 19107 19672 19340 19700
rect 19107 19669 19119 19672
rect 19061 19663 19119 19669
rect 19334 19660 19340 19672
rect 19392 19660 19398 19712
rect 20364 19700 20392 19876
rect 20533 19873 20545 19907
rect 20579 19904 20591 19907
rect 22388 19904 22416 19944
rect 23032 19916 23060 19944
rect 23290 19932 23296 19984
rect 23348 19932 23354 19984
rect 20579 19876 22416 19904
rect 20579 19873 20591 19876
rect 20533 19867 20591 19873
rect 22830 19864 22836 19916
rect 22888 19864 22894 19916
rect 23014 19864 23020 19916
rect 23072 19904 23078 19916
rect 24397 19907 24455 19913
rect 24397 19904 24409 19907
rect 23072 19876 24409 19904
rect 23072 19864 23078 19876
rect 24397 19873 24409 19876
rect 24443 19873 24455 19907
rect 24397 19867 24455 19873
rect 21910 19796 21916 19848
rect 21968 19796 21974 19848
rect 22186 19796 22192 19848
rect 22244 19836 22250 19848
rect 22741 19839 22799 19845
rect 22741 19836 22753 19839
rect 22244 19808 22753 19836
rect 22244 19796 22250 19808
rect 22741 19805 22753 19808
rect 22787 19805 22799 19839
rect 22741 19799 22799 19805
rect 22848 19808 23520 19836
rect 22848 19768 22876 19808
rect 22112 19740 22876 19768
rect 23293 19771 23351 19777
rect 22112 19700 22140 19740
rect 23293 19737 23305 19771
rect 23339 19768 23351 19771
rect 23382 19768 23388 19780
rect 23339 19740 23388 19768
rect 23339 19737 23351 19740
rect 23293 19731 23351 19737
rect 23382 19728 23388 19740
rect 23440 19728 23446 19780
rect 23492 19768 23520 19808
rect 23566 19796 23572 19848
rect 23624 19796 23630 19848
rect 24302 19768 24308 19780
rect 23492 19740 24308 19768
rect 24302 19728 24308 19740
rect 24360 19768 24366 19780
rect 24673 19771 24731 19777
rect 24673 19768 24685 19771
rect 24360 19740 24685 19768
rect 24360 19728 24366 19740
rect 24673 19737 24685 19740
rect 24719 19737 24731 19771
rect 24673 19731 24731 19737
rect 24780 19740 25162 19768
rect 20364 19672 22140 19700
rect 22186 19660 22192 19712
rect 22244 19700 22250 19712
rect 22281 19703 22339 19709
rect 22281 19700 22293 19703
rect 22244 19672 22293 19700
rect 22244 19660 22250 19672
rect 22281 19669 22293 19672
rect 22327 19669 22339 19703
rect 22281 19663 22339 19669
rect 23474 19660 23480 19712
rect 23532 19660 23538 19712
rect 24210 19660 24216 19712
rect 24268 19700 24274 19712
rect 24780 19700 24808 19740
rect 24268 19672 24808 19700
rect 24268 19660 24274 19672
rect 1104 19610 28888 19632
rect 1104 19558 3658 19610
rect 3710 19558 3722 19610
rect 3774 19558 3786 19610
rect 3838 19558 3850 19610
rect 3902 19558 3914 19610
rect 3966 19558 3978 19610
rect 4030 19558 11658 19610
rect 11710 19558 11722 19610
rect 11774 19558 11786 19610
rect 11838 19558 11850 19610
rect 11902 19558 11914 19610
rect 11966 19558 11978 19610
rect 12030 19558 19658 19610
rect 19710 19558 19722 19610
rect 19774 19558 19786 19610
rect 19838 19558 19850 19610
rect 19902 19558 19914 19610
rect 19966 19558 19978 19610
rect 20030 19558 27658 19610
rect 27710 19558 27722 19610
rect 27774 19558 27786 19610
rect 27838 19558 27850 19610
rect 27902 19558 27914 19610
rect 27966 19558 27978 19610
rect 28030 19558 28888 19610
rect 1104 19536 28888 19558
rect 1581 19499 1639 19505
rect 1581 19465 1593 19499
rect 1627 19465 1639 19499
rect 1581 19459 1639 19465
rect 2317 19499 2375 19505
rect 2317 19465 2329 19499
rect 2363 19496 2375 19499
rect 2682 19496 2688 19508
rect 2363 19468 2688 19496
rect 2363 19465 2375 19468
rect 2317 19459 2375 19465
rect 1596 19428 1624 19459
rect 2682 19456 2688 19468
rect 2740 19456 2746 19508
rect 3050 19456 3056 19508
rect 3108 19496 3114 19508
rect 3970 19496 3976 19508
rect 3108 19468 3976 19496
rect 3108 19456 3114 19468
rect 3970 19456 3976 19468
rect 4028 19456 4034 19508
rect 6178 19456 6184 19508
rect 6236 19456 6242 19508
rect 6730 19456 6736 19508
rect 6788 19496 6794 19508
rect 6788 19468 7604 19496
rect 6788 19456 6794 19468
rect 4522 19428 4528 19440
rect 1596 19400 4528 19428
rect 4522 19388 4528 19400
rect 4580 19428 4586 19440
rect 7466 19428 7472 19440
rect 4580 19400 6500 19428
rect 4580 19388 4586 19400
rect 1394 19320 1400 19372
rect 1452 19360 1458 19372
rect 1673 19363 1731 19369
rect 1673 19360 1685 19363
rect 1452 19332 1685 19360
rect 1452 19320 1458 19332
rect 1673 19329 1685 19332
rect 1719 19329 1731 19363
rect 1673 19323 1731 19329
rect 2225 19363 2283 19369
rect 2225 19329 2237 19363
rect 2271 19360 2283 19363
rect 2682 19360 2688 19372
rect 2271 19332 2688 19360
rect 2271 19329 2283 19332
rect 2225 19323 2283 19329
rect 2682 19320 2688 19332
rect 2740 19320 2746 19372
rect 2866 19320 2872 19372
rect 2924 19360 2930 19372
rect 2961 19363 3019 19369
rect 2961 19360 2973 19363
rect 2924 19332 2973 19360
rect 2924 19320 2930 19332
rect 2961 19329 2973 19332
rect 3007 19329 3019 19363
rect 2961 19323 3019 19329
rect 3418 19320 3424 19372
rect 3476 19360 3482 19372
rect 3881 19363 3939 19369
rect 3881 19360 3893 19363
rect 3476 19332 3893 19360
rect 3476 19320 3482 19332
rect 3881 19329 3893 19332
rect 3927 19360 3939 19363
rect 4062 19360 4068 19372
rect 3927 19332 4068 19360
rect 3927 19329 3939 19332
rect 3881 19323 3939 19329
rect 4062 19320 4068 19332
rect 4120 19320 4126 19372
rect 5353 19363 5411 19369
rect 5353 19360 5365 19363
rect 4172 19332 5365 19360
rect 3050 19252 3056 19304
rect 3108 19292 3114 19304
rect 3694 19292 3700 19304
rect 3108 19264 3700 19292
rect 3108 19252 3114 19264
rect 3694 19252 3700 19264
rect 3752 19252 3758 19304
rect 3786 19252 3792 19304
rect 3844 19252 3850 19304
rect 3970 19252 3976 19304
rect 4028 19292 4034 19304
rect 4172 19292 4200 19332
rect 5353 19329 5365 19332
rect 5399 19360 5411 19363
rect 5399 19332 5580 19360
rect 5399 19329 5411 19332
rect 5353 19323 5411 19329
rect 4028 19264 4200 19292
rect 5552 19292 5580 19332
rect 5626 19320 5632 19372
rect 5684 19320 5690 19372
rect 5810 19320 5816 19372
rect 5868 19320 5874 19372
rect 5902 19320 5908 19372
rect 5960 19320 5966 19372
rect 5994 19320 6000 19372
rect 6052 19320 6058 19372
rect 6362 19360 6368 19372
rect 6104 19332 6368 19360
rect 6104 19292 6132 19332
rect 6362 19320 6368 19332
rect 6420 19320 6426 19372
rect 6472 19334 6500 19400
rect 6656 19400 7052 19428
rect 6656 19359 6684 19400
rect 6633 19353 6691 19359
rect 6633 19334 6645 19353
rect 6472 19319 6645 19334
rect 6679 19319 6691 19353
rect 6730 19320 6736 19372
rect 6788 19320 6794 19372
rect 7024 19369 7052 19400
rect 7116 19400 7472 19428
rect 7116 19369 7144 19400
rect 7466 19388 7472 19400
rect 7524 19388 7530 19440
rect 7576 19369 7604 19468
rect 8202 19456 8208 19508
rect 8260 19456 8266 19508
rect 8297 19499 8355 19505
rect 8297 19465 8309 19499
rect 8343 19496 8355 19499
rect 9398 19496 9404 19508
rect 8343 19468 9404 19496
rect 8343 19465 8355 19468
rect 8297 19459 8355 19465
rect 9398 19456 9404 19468
rect 9456 19456 9462 19508
rect 9677 19499 9735 19505
rect 9677 19465 9689 19499
rect 9723 19496 9735 19499
rect 9766 19496 9772 19508
rect 9723 19468 9772 19496
rect 9723 19465 9735 19468
rect 9677 19459 9735 19465
rect 9766 19456 9772 19468
rect 9824 19456 9830 19508
rect 12345 19499 12403 19505
rect 12345 19465 12357 19499
rect 12391 19496 12403 19499
rect 12526 19496 12532 19508
rect 12391 19468 12532 19496
rect 12391 19465 12403 19468
rect 12345 19459 12403 19465
rect 12526 19456 12532 19468
rect 12584 19456 12590 19508
rect 23382 19456 23388 19508
rect 23440 19496 23446 19508
rect 24765 19499 24823 19505
rect 24765 19496 24777 19499
rect 23440 19468 24777 19496
rect 23440 19456 23446 19468
rect 24765 19465 24777 19468
rect 24811 19465 24823 19499
rect 24765 19459 24823 19465
rect 9858 19428 9864 19440
rect 9600 19400 9864 19428
rect 7009 19363 7067 19369
rect 7009 19329 7021 19363
rect 7055 19329 7067 19363
rect 7009 19323 7067 19329
rect 7101 19363 7159 19369
rect 7101 19329 7113 19363
rect 7147 19329 7159 19363
rect 7377 19363 7435 19369
rect 7377 19360 7389 19363
rect 7101 19323 7159 19329
rect 7208 19332 7389 19360
rect 6472 19313 6691 19319
rect 6472 19306 6684 19313
rect 5552 19264 6132 19292
rect 4028 19252 4034 19264
rect 6822 19252 6828 19304
rect 6880 19292 6886 19304
rect 7208 19292 7236 19332
rect 7377 19329 7389 19332
rect 7423 19329 7435 19363
rect 7377 19323 7435 19329
rect 7561 19363 7619 19369
rect 7561 19329 7573 19363
rect 7607 19329 7619 19363
rect 7561 19323 7619 19329
rect 8018 19320 8024 19372
rect 8076 19320 8082 19372
rect 9600 19369 9628 19400
rect 9858 19388 9864 19400
rect 9916 19388 9922 19440
rect 18138 19388 18144 19440
rect 18196 19388 18202 19440
rect 18782 19388 18788 19440
rect 18840 19388 18846 19440
rect 23290 19428 23296 19440
rect 22940 19400 23296 19428
rect 8389 19363 8447 19369
rect 8389 19329 8401 19363
rect 8435 19329 8447 19363
rect 8389 19323 8447 19329
rect 9585 19363 9643 19369
rect 9585 19329 9597 19363
rect 9631 19329 9643 19363
rect 9585 19323 9643 19329
rect 9769 19363 9827 19369
rect 9769 19329 9781 19363
rect 9815 19360 9827 19363
rect 10226 19360 10232 19372
rect 9815 19332 10232 19360
rect 9815 19329 9827 19332
rect 9769 19323 9827 19329
rect 7926 19292 7932 19304
rect 6880 19264 7236 19292
rect 7300 19264 7932 19292
rect 6880 19252 6886 19264
rect 3234 19184 3240 19236
rect 3292 19184 3298 19236
rect 3326 19184 3332 19236
rect 3384 19224 3390 19236
rect 3384 19196 3740 19224
rect 3384 19184 3390 19196
rect 2130 19116 2136 19168
rect 2188 19156 2194 19168
rect 2958 19156 2964 19168
rect 2188 19128 2964 19156
rect 2188 19116 2194 19128
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 3418 19116 3424 19168
rect 3476 19116 3482 19168
rect 3513 19159 3571 19165
rect 3513 19125 3525 19159
rect 3559 19156 3571 19159
rect 3602 19156 3608 19168
rect 3559 19128 3608 19156
rect 3559 19125 3571 19128
rect 3513 19119 3571 19125
rect 3602 19116 3608 19128
rect 3660 19116 3666 19168
rect 3712 19165 3740 19196
rect 5626 19184 5632 19236
rect 5684 19224 5690 19236
rect 6549 19227 6607 19233
rect 6549 19224 6561 19227
rect 5684 19196 6561 19224
rect 5684 19184 5690 19196
rect 6549 19193 6561 19196
rect 6595 19224 6607 19227
rect 7300 19224 7328 19264
rect 7926 19252 7932 19264
rect 7984 19252 7990 19304
rect 8404 19224 8432 19323
rect 10226 19320 10232 19332
rect 10284 19320 10290 19372
rect 12713 19363 12771 19369
rect 12713 19329 12725 19363
rect 12759 19360 12771 19363
rect 15102 19360 15108 19372
rect 12759 19332 15108 19360
rect 12759 19329 12771 19332
rect 12713 19323 12771 19329
rect 15102 19320 15108 19332
rect 15160 19320 15166 19372
rect 15286 19320 15292 19372
rect 15344 19320 15350 19372
rect 16850 19320 16856 19372
rect 16908 19360 16914 19372
rect 17865 19363 17923 19369
rect 17865 19360 17877 19363
rect 16908 19332 17877 19360
rect 16908 19320 16914 19332
rect 17865 19329 17877 19332
rect 17911 19329 17923 19363
rect 17865 19323 17923 19329
rect 22738 19320 22744 19372
rect 22796 19320 22802 19372
rect 22940 19369 22968 19400
rect 23290 19388 23296 19400
rect 23348 19388 23354 19440
rect 24026 19388 24032 19440
rect 24084 19388 24090 19440
rect 22925 19363 22983 19369
rect 22925 19329 22937 19363
rect 22971 19329 22983 19363
rect 22925 19323 22983 19329
rect 23014 19320 23020 19372
rect 23072 19320 23078 19372
rect 12802 19252 12808 19304
rect 12860 19252 12866 19304
rect 12894 19252 12900 19304
rect 12952 19252 12958 19304
rect 22833 19295 22891 19301
rect 22833 19261 22845 19295
rect 22879 19292 22891 19295
rect 23293 19295 23351 19301
rect 23293 19292 23305 19295
rect 22879 19264 23305 19292
rect 22879 19261 22891 19264
rect 22833 19255 22891 19261
rect 23293 19261 23305 19264
rect 23339 19261 23351 19295
rect 23293 19255 23351 19261
rect 6595 19196 7328 19224
rect 7392 19196 8432 19224
rect 6595 19193 6607 19196
rect 6549 19187 6607 19193
rect 3697 19159 3755 19165
rect 3697 19125 3709 19159
rect 3743 19125 3755 19159
rect 3697 19119 3755 19125
rect 5445 19159 5503 19165
rect 5445 19125 5457 19159
rect 5491 19156 5503 19159
rect 5534 19156 5540 19168
rect 5491 19128 5540 19156
rect 5491 19125 5503 19128
rect 5445 19119 5503 19125
rect 5534 19116 5540 19128
rect 5592 19156 5598 19168
rect 5902 19156 5908 19168
rect 5592 19128 5908 19156
rect 5592 19116 5598 19128
rect 5902 19116 5908 19128
rect 5960 19116 5966 19168
rect 7285 19159 7343 19165
rect 7285 19125 7297 19159
rect 7331 19156 7343 19159
rect 7392 19156 7420 19196
rect 7331 19128 7420 19156
rect 7469 19159 7527 19165
rect 7331 19125 7343 19128
rect 7285 19119 7343 19125
rect 7469 19125 7481 19159
rect 7515 19156 7527 19159
rect 8202 19156 8208 19168
rect 7515 19128 8208 19156
rect 7515 19125 7527 19128
rect 7469 19119 7527 19125
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 8665 19159 8723 19165
rect 8665 19125 8677 19159
rect 8711 19156 8723 19159
rect 9214 19156 9220 19168
rect 8711 19128 9220 19156
rect 8711 19125 8723 19128
rect 8665 19119 8723 19125
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 15470 19116 15476 19168
rect 15528 19116 15534 19168
rect 19334 19116 19340 19168
rect 19392 19156 19398 19168
rect 19613 19159 19671 19165
rect 19613 19156 19625 19159
rect 19392 19128 19625 19156
rect 19392 19116 19398 19128
rect 19613 19125 19625 19128
rect 19659 19156 19671 19159
rect 19797 19159 19855 19165
rect 19797 19156 19809 19159
rect 19659 19128 19809 19156
rect 19659 19125 19671 19128
rect 19613 19119 19671 19125
rect 19797 19125 19809 19128
rect 19843 19156 19855 19159
rect 20438 19156 20444 19168
rect 19843 19128 20444 19156
rect 19843 19125 19855 19128
rect 19797 19119 19855 19125
rect 20438 19116 20444 19128
rect 20496 19116 20502 19168
rect 1104 19066 28888 19088
rect 1104 19014 2918 19066
rect 2970 19014 2982 19066
rect 3034 19014 3046 19066
rect 3098 19014 3110 19066
rect 3162 19014 3174 19066
rect 3226 19014 3238 19066
rect 3290 19014 10918 19066
rect 10970 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 11238 19066
rect 11290 19014 18918 19066
rect 18970 19014 18982 19066
rect 19034 19014 19046 19066
rect 19098 19014 19110 19066
rect 19162 19014 19174 19066
rect 19226 19014 19238 19066
rect 19290 19014 26918 19066
rect 26970 19014 26982 19066
rect 27034 19014 27046 19066
rect 27098 19014 27110 19066
rect 27162 19014 27174 19066
rect 27226 19014 27238 19066
rect 27290 19014 28888 19066
rect 1104 18992 28888 19014
rect 2961 18955 3019 18961
rect 2961 18921 2973 18955
rect 3007 18952 3019 18955
rect 3234 18952 3240 18964
rect 3007 18924 3240 18952
rect 3007 18921 3019 18924
rect 2961 18915 3019 18921
rect 3234 18912 3240 18924
rect 3292 18912 3298 18964
rect 3418 18912 3424 18964
rect 3476 18952 3482 18964
rect 4157 18955 4215 18961
rect 4157 18952 4169 18955
rect 3476 18924 4169 18952
rect 3476 18912 3482 18924
rect 4157 18921 4169 18924
rect 4203 18921 4215 18955
rect 4157 18915 4215 18921
rect 4246 18912 4252 18964
rect 4304 18912 4310 18964
rect 12802 18912 12808 18964
rect 12860 18952 12866 18964
rect 13173 18955 13231 18961
rect 13173 18952 13185 18955
rect 12860 18924 13185 18952
rect 12860 18912 12866 18924
rect 13173 18921 13185 18924
rect 13219 18921 13231 18955
rect 13173 18915 13231 18921
rect 14458 18912 14464 18964
rect 14516 18912 14522 18964
rect 22186 18912 22192 18964
rect 22244 18912 22250 18964
rect 22738 18912 22744 18964
rect 22796 18952 22802 18964
rect 23201 18955 23259 18961
rect 23201 18952 23213 18955
rect 22796 18924 23213 18952
rect 22796 18912 22802 18924
rect 23201 18921 23213 18924
rect 23247 18921 23259 18955
rect 23201 18915 23259 18921
rect 23382 18912 23388 18964
rect 23440 18912 23446 18964
rect 24302 18912 24308 18964
rect 24360 18952 24366 18964
rect 24397 18955 24455 18961
rect 24397 18952 24409 18955
rect 24360 18924 24409 18952
rect 24360 18912 24366 18924
rect 24397 18921 24409 18924
rect 24443 18921 24455 18955
rect 24397 18915 24455 18921
rect 3602 18844 3608 18896
rect 3660 18884 3666 18896
rect 4264 18884 4292 18912
rect 3660 18856 4292 18884
rect 3660 18844 3666 18856
rect 2590 18816 2596 18828
rect 2424 18788 2596 18816
rect 1302 18708 1308 18760
rect 1360 18748 1366 18760
rect 2424 18757 2452 18788
rect 2590 18776 2596 18788
rect 2648 18776 2654 18828
rect 3142 18776 3148 18828
rect 3200 18816 3206 18828
rect 3329 18819 3387 18825
rect 3329 18816 3341 18819
rect 3200 18788 3341 18816
rect 3200 18776 3206 18788
rect 3329 18785 3341 18788
rect 3375 18816 3387 18819
rect 4249 18819 4307 18825
rect 4249 18816 4261 18819
rect 3375 18788 4261 18816
rect 3375 18785 3387 18788
rect 3329 18779 3387 18785
rect 4249 18785 4261 18788
rect 4295 18785 4307 18819
rect 4249 18779 4307 18785
rect 11241 18819 11299 18825
rect 11241 18785 11253 18819
rect 11287 18816 11299 18819
rect 11287 18788 12848 18816
rect 11287 18785 11299 18788
rect 11241 18779 11299 18785
rect 12820 18760 12848 18788
rect 14182 18776 14188 18828
rect 14240 18816 14246 18828
rect 14240 18788 16252 18816
rect 14240 18776 14246 18788
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 1360 18720 1409 18748
rect 1360 18708 1366 18720
rect 1397 18717 1409 18720
rect 1443 18748 1455 18751
rect 1673 18751 1731 18757
rect 1673 18748 1685 18751
rect 1443 18720 1685 18748
rect 1443 18717 1455 18720
rect 1397 18711 1455 18717
rect 1673 18717 1685 18720
rect 1719 18717 1731 18751
rect 1673 18711 1731 18717
rect 2409 18751 2467 18757
rect 2409 18717 2421 18751
rect 2455 18717 2467 18751
rect 2409 18711 2467 18717
rect 2777 18751 2835 18757
rect 2777 18717 2789 18751
rect 2823 18748 2835 18751
rect 2866 18748 2872 18760
rect 2823 18720 2872 18748
rect 2823 18717 2835 18720
rect 2777 18711 2835 18717
rect 2866 18708 2872 18720
rect 2924 18708 2930 18760
rect 3053 18751 3111 18757
rect 3053 18717 3065 18751
rect 3099 18748 3111 18751
rect 3234 18748 3240 18760
rect 3099 18720 3240 18748
rect 3099 18717 3111 18720
rect 3053 18711 3111 18717
rect 3234 18708 3240 18720
rect 3292 18708 3298 18760
rect 3510 18708 3516 18760
rect 3568 18748 3574 18760
rect 4065 18751 4123 18757
rect 4065 18748 4077 18751
rect 3568 18720 4077 18748
rect 3568 18708 3574 18720
rect 4065 18717 4077 18720
rect 4111 18717 4123 18751
rect 4065 18711 4123 18717
rect 4522 18708 4528 18760
rect 4580 18708 4586 18760
rect 11330 18708 11336 18760
rect 11388 18748 11394 18760
rect 11425 18751 11483 18757
rect 11425 18748 11437 18751
rect 11388 18720 11437 18748
rect 11388 18708 11394 18720
rect 11425 18717 11437 18720
rect 11471 18717 11483 18751
rect 11425 18711 11483 18717
rect 12802 18708 12808 18760
rect 12860 18708 12866 18760
rect 16224 18757 16252 18788
rect 16209 18751 16267 18757
rect 16209 18717 16221 18751
rect 16255 18748 16267 18751
rect 16850 18748 16856 18760
rect 16255 18720 16856 18748
rect 16255 18717 16267 18720
rect 16209 18711 16267 18717
rect 16850 18708 16856 18720
rect 16908 18708 16914 18760
rect 21818 18708 21824 18760
rect 21876 18708 21882 18760
rect 24578 18708 24584 18760
rect 24636 18708 24642 18760
rect 24673 18751 24731 18757
rect 24673 18717 24685 18751
rect 24719 18717 24731 18751
rect 24673 18711 24731 18717
rect 2222 18640 2228 18692
rect 2280 18680 2286 18692
rect 2593 18683 2651 18689
rect 2593 18680 2605 18683
rect 2280 18652 2605 18680
rect 2280 18640 2286 18652
rect 2593 18649 2605 18652
rect 2639 18649 2651 18683
rect 2593 18643 2651 18649
rect 2682 18640 2688 18692
rect 2740 18640 2746 18692
rect 6730 18680 6736 18692
rect 3436 18652 6736 18680
rect 1581 18615 1639 18621
rect 1581 18581 1593 18615
rect 1627 18612 1639 18615
rect 3436 18612 3464 18652
rect 6730 18640 6736 18652
rect 6788 18640 6794 18692
rect 11701 18683 11759 18689
rect 11701 18649 11713 18683
rect 11747 18649 11759 18683
rect 15502 18652 15608 18680
rect 11701 18643 11759 18649
rect 1627 18584 3464 18612
rect 1627 18581 1639 18584
rect 1581 18575 1639 18581
rect 3510 18572 3516 18624
rect 3568 18612 3574 18624
rect 3605 18615 3663 18621
rect 3605 18612 3617 18615
rect 3568 18584 3617 18612
rect 3568 18572 3574 18584
rect 3605 18581 3617 18584
rect 3651 18581 3663 18615
rect 3605 18575 3663 18581
rect 3786 18572 3792 18624
rect 3844 18572 3850 18624
rect 4430 18572 4436 18624
rect 4488 18572 4494 18624
rect 11716 18612 11744 18643
rect 15580 18624 15608 18652
rect 15930 18640 15936 18692
rect 15988 18640 15994 18692
rect 23198 18640 23204 18692
rect 23256 18680 23262 18692
rect 23353 18683 23411 18689
rect 23353 18680 23365 18683
rect 23256 18652 23365 18680
rect 23256 18640 23262 18652
rect 23353 18649 23365 18652
rect 23399 18649 23411 18683
rect 23353 18643 23411 18649
rect 23474 18640 23480 18692
rect 23532 18680 23538 18692
rect 23569 18683 23627 18689
rect 23569 18680 23581 18683
rect 23532 18652 23581 18680
rect 23532 18640 23538 18652
rect 23569 18649 23581 18652
rect 23615 18649 23627 18683
rect 23569 18643 23627 18649
rect 24486 18640 24492 18692
rect 24544 18680 24550 18692
rect 24688 18680 24716 18711
rect 24544 18652 24716 18680
rect 24544 18640 24550 18652
rect 12066 18612 12072 18624
rect 11716 18584 12072 18612
rect 12066 18572 12072 18584
rect 12124 18572 12130 18624
rect 15562 18572 15568 18624
rect 15620 18572 15626 18624
rect 22094 18572 22100 18624
rect 22152 18612 22158 18624
rect 22189 18615 22247 18621
rect 22189 18612 22201 18615
rect 22152 18584 22201 18612
rect 22152 18572 22158 18584
rect 22189 18581 22201 18584
rect 22235 18581 22247 18615
rect 22189 18575 22247 18581
rect 22370 18572 22376 18624
rect 22428 18572 22434 18624
rect 1104 18522 28888 18544
rect 1104 18470 3658 18522
rect 3710 18470 3722 18522
rect 3774 18470 3786 18522
rect 3838 18470 3850 18522
rect 3902 18470 3914 18522
rect 3966 18470 3978 18522
rect 4030 18470 11658 18522
rect 11710 18470 11722 18522
rect 11774 18470 11786 18522
rect 11838 18470 11850 18522
rect 11902 18470 11914 18522
rect 11966 18470 11978 18522
rect 12030 18470 19658 18522
rect 19710 18470 19722 18522
rect 19774 18470 19786 18522
rect 19838 18470 19850 18522
rect 19902 18470 19914 18522
rect 19966 18470 19978 18522
rect 20030 18470 27658 18522
rect 27710 18470 27722 18522
rect 27774 18470 27786 18522
rect 27838 18470 27850 18522
rect 27902 18470 27914 18522
rect 27966 18470 27978 18522
rect 28030 18470 28888 18522
rect 1104 18448 28888 18470
rect 3142 18368 3148 18420
rect 3200 18368 3206 18420
rect 4430 18408 4436 18420
rect 3344 18380 4436 18408
rect 2130 18300 2136 18352
rect 2188 18340 2194 18352
rect 2590 18340 2596 18352
rect 2188 18312 2596 18340
rect 2188 18300 2194 18312
rect 2590 18300 2596 18312
rect 2648 18300 2654 18352
rect 1302 18232 1308 18284
rect 1360 18272 1366 18284
rect 1489 18275 1547 18281
rect 1489 18272 1501 18275
rect 1360 18244 1501 18272
rect 1360 18232 1366 18244
rect 1489 18241 1501 18244
rect 1535 18272 1547 18275
rect 1765 18275 1823 18281
rect 1765 18272 1777 18275
rect 1535 18244 1777 18272
rect 1535 18241 1547 18244
rect 1489 18235 1547 18241
rect 1765 18241 1777 18244
rect 1811 18241 1823 18275
rect 1765 18235 1823 18241
rect 2314 18232 2320 18284
rect 2372 18272 2378 18284
rect 3344 18272 3372 18380
rect 4430 18368 4436 18380
rect 4488 18368 4494 18420
rect 9125 18411 9183 18417
rect 9125 18377 9137 18411
rect 9171 18408 9183 18411
rect 9171 18380 10824 18408
rect 9171 18377 9183 18380
rect 9125 18371 9183 18377
rect 3510 18300 3516 18352
rect 3568 18340 3574 18352
rect 3789 18343 3847 18349
rect 3568 18312 3740 18340
rect 3568 18300 3574 18312
rect 2372 18244 3372 18272
rect 2372 18232 2378 18244
rect 3418 18232 3424 18284
rect 3476 18272 3482 18284
rect 3605 18275 3663 18281
rect 3605 18272 3617 18275
rect 3476 18244 3617 18272
rect 3476 18232 3482 18244
rect 3605 18241 3617 18244
rect 3651 18241 3663 18275
rect 3712 18272 3740 18312
rect 3789 18309 3801 18343
rect 3835 18340 3847 18343
rect 4065 18343 4123 18349
rect 4065 18340 4077 18343
rect 3835 18312 4077 18340
rect 3835 18309 3847 18312
rect 3789 18303 3847 18309
rect 4065 18309 4077 18312
rect 4111 18309 4123 18343
rect 9490 18340 9496 18352
rect 4065 18303 4123 18309
rect 9324 18312 9496 18340
rect 3881 18275 3939 18281
rect 3881 18272 3893 18275
rect 3712 18244 3893 18272
rect 3605 18235 3663 18241
rect 3881 18241 3893 18244
rect 3927 18241 3939 18275
rect 3881 18235 3939 18241
rect 3970 18232 3976 18284
rect 4028 18232 4034 18284
rect 9324 18281 9352 18312
rect 9490 18300 9496 18312
rect 9548 18300 9554 18352
rect 9769 18343 9827 18349
rect 9769 18309 9781 18343
rect 9815 18340 9827 18343
rect 10134 18340 10140 18352
rect 9815 18312 10140 18340
rect 9815 18309 9827 18312
rect 9769 18303 9827 18309
rect 10134 18300 10140 18312
rect 10192 18300 10198 18352
rect 10796 18340 10824 18380
rect 12066 18368 12072 18420
rect 12124 18408 12130 18420
rect 12161 18411 12219 18417
rect 12161 18408 12173 18411
rect 12124 18380 12173 18408
rect 12124 18368 12130 18380
rect 12161 18377 12173 18380
rect 12207 18377 12219 18411
rect 12161 18371 12219 18377
rect 12529 18411 12587 18417
rect 12529 18377 12541 18411
rect 12575 18408 12587 18411
rect 12710 18408 12716 18420
rect 12575 18380 12716 18408
rect 12575 18377 12587 18380
rect 12529 18371 12587 18377
rect 12710 18368 12716 18380
rect 12768 18368 12774 18420
rect 15102 18368 15108 18420
rect 15160 18408 15166 18420
rect 15933 18411 15991 18417
rect 15933 18408 15945 18411
rect 15160 18380 15945 18408
rect 15160 18368 15166 18380
rect 15933 18377 15945 18380
rect 15979 18377 15991 18411
rect 15933 18371 15991 18377
rect 22094 18368 22100 18420
rect 22152 18408 22158 18420
rect 24486 18408 24492 18420
rect 22152 18380 24492 18408
rect 22152 18368 22158 18380
rect 24486 18368 24492 18380
rect 24544 18368 24550 18420
rect 12434 18340 12440 18352
rect 10796 18312 12440 18340
rect 12434 18300 12440 18312
rect 12492 18300 12498 18352
rect 23382 18300 23388 18352
rect 23440 18300 23446 18352
rect 9309 18275 9367 18281
rect 9309 18241 9321 18275
rect 9355 18241 9367 18275
rect 9309 18235 9367 18241
rect 9398 18232 9404 18284
rect 9456 18232 9462 18284
rect 9582 18232 9588 18284
rect 9640 18232 9646 18284
rect 9677 18275 9735 18281
rect 9677 18241 9689 18275
rect 9723 18241 9735 18275
rect 9677 18235 9735 18241
rect 2130 18164 2136 18216
rect 2188 18204 2194 18216
rect 2682 18204 2688 18216
rect 2188 18176 2688 18204
rect 2188 18164 2194 18176
rect 2682 18164 2688 18176
rect 2740 18164 2746 18216
rect 2866 18164 2872 18216
rect 2924 18204 2930 18216
rect 5534 18204 5540 18216
rect 2924 18176 5540 18204
rect 2924 18164 2930 18176
rect 5534 18164 5540 18176
rect 5592 18164 5598 18216
rect 9214 18164 9220 18216
rect 9272 18204 9278 18216
rect 9600 18204 9628 18232
rect 9272 18176 9628 18204
rect 9692 18204 9720 18235
rect 9858 18232 9864 18284
rect 9916 18272 9922 18284
rect 9953 18275 10011 18281
rect 9953 18272 9965 18275
rect 9916 18244 9965 18272
rect 9916 18232 9922 18244
rect 9953 18241 9965 18244
rect 9999 18241 10011 18275
rect 9953 18235 10011 18241
rect 10045 18275 10103 18281
rect 10045 18241 10057 18275
rect 10091 18241 10103 18275
rect 10045 18235 10103 18241
rect 9692 18176 9812 18204
rect 9272 18164 9278 18176
rect 3050 18096 3056 18148
rect 3108 18096 3114 18148
rect 8478 18096 8484 18148
rect 8536 18136 8542 18148
rect 9784 18145 9812 18176
rect 9769 18139 9827 18145
rect 8536 18108 9720 18136
rect 8536 18096 8542 18108
rect 1578 18028 1584 18080
rect 1636 18028 1642 18080
rect 3418 18028 3424 18080
rect 3476 18028 3482 18080
rect 9490 18028 9496 18080
rect 9548 18068 9554 18080
rect 9585 18071 9643 18077
rect 9585 18068 9597 18071
rect 9548 18040 9597 18068
rect 9548 18028 9554 18040
rect 9585 18037 9597 18040
rect 9631 18037 9643 18071
rect 9692 18068 9720 18108
rect 9769 18105 9781 18139
rect 9815 18105 9827 18139
rect 9769 18099 9827 18105
rect 10060 18068 10088 18235
rect 14182 18232 14188 18284
rect 14240 18232 14246 18284
rect 15562 18232 15568 18284
rect 15620 18272 15626 18284
rect 16209 18275 16267 18281
rect 15620 18244 16068 18272
rect 15620 18232 15626 18244
rect 12618 18164 12624 18216
rect 12676 18164 12682 18216
rect 12713 18207 12771 18213
rect 12713 18173 12725 18207
rect 12759 18173 12771 18207
rect 12713 18167 12771 18173
rect 12069 18139 12127 18145
rect 12069 18105 12081 18139
rect 12115 18136 12127 18139
rect 12158 18136 12164 18148
rect 12115 18108 12164 18136
rect 12115 18105 12127 18108
rect 12069 18099 12127 18105
rect 12158 18096 12164 18108
rect 12216 18136 12222 18148
rect 12728 18136 12756 18167
rect 14458 18164 14464 18216
rect 14516 18164 14522 18216
rect 12216 18108 12756 18136
rect 12216 18096 12222 18108
rect 16040 18077 16068 18244
rect 16209 18241 16221 18275
rect 16255 18272 16267 18275
rect 16482 18272 16488 18284
rect 16255 18244 16488 18272
rect 16255 18241 16267 18244
rect 16209 18235 16267 18241
rect 16482 18232 16488 18244
rect 16540 18232 16546 18284
rect 20898 18232 20904 18284
rect 20956 18232 20962 18284
rect 21085 18275 21143 18281
rect 21085 18241 21097 18275
rect 21131 18272 21143 18275
rect 21131 18244 22094 18272
rect 21131 18241 21143 18244
rect 21085 18235 21143 18241
rect 22066 18204 22094 18244
rect 22370 18232 22376 18284
rect 22428 18272 22434 18284
rect 23201 18275 23259 18281
rect 23201 18272 23213 18275
rect 22428 18244 23213 18272
rect 22428 18232 22434 18244
rect 23201 18241 23213 18244
rect 23247 18241 23259 18275
rect 23201 18235 23259 18241
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18272 23351 18275
rect 23400 18272 23428 18300
rect 23339 18244 23428 18272
rect 23339 18241 23351 18244
rect 23293 18235 23351 18241
rect 22066 18176 23244 18204
rect 23216 18148 23244 18176
rect 23382 18164 23388 18216
rect 23440 18164 23446 18216
rect 23477 18207 23535 18213
rect 23477 18173 23489 18207
rect 23523 18204 23535 18207
rect 24578 18204 24584 18216
rect 23523 18176 24584 18204
rect 23523 18173 23535 18176
rect 23477 18167 23535 18173
rect 24578 18164 24584 18176
rect 24636 18164 24642 18216
rect 23198 18096 23204 18148
rect 23256 18096 23262 18148
rect 9692 18040 10088 18068
rect 16025 18071 16083 18077
rect 9585 18031 9643 18037
rect 16025 18037 16037 18071
rect 16071 18068 16083 18071
rect 18230 18068 18236 18080
rect 16071 18040 18236 18068
rect 16071 18037 16083 18040
rect 16025 18031 16083 18037
rect 18230 18028 18236 18040
rect 18288 18028 18294 18080
rect 20806 18028 20812 18080
rect 20864 18068 20870 18080
rect 20901 18071 20959 18077
rect 20901 18068 20913 18071
rect 20864 18040 20913 18068
rect 20864 18028 20870 18040
rect 20901 18037 20913 18040
rect 20947 18037 20959 18071
rect 20901 18031 20959 18037
rect 23017 18071 23075 18077
rect 23017 18037 23029 18071
rect 23063 18068 23075 18071
rect 23106 18068 23112 18080
rect 23063 18040 23112 18068
rect 23063 18037 23075 18040
rect 23017 18031 23075 18037
rect 23106 18028 23112 18040
rect 23164 18028 23170 18080
rect 1104 17978 28888 18000
rect 1104 17926 2918 17978
rect 2970 17926 2982 17978
rect 3034 17926 3046 17978
rect 3098 17926 3110 17978
rect 3162 17926 3174 17978
rect 3226 17926 3238 17978
rect 3290 17926 10918 17978
rect 10970 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 11238 17978
rect 11290 17926 18918 17978
rect 18970 17926 18982 17978
rect 19034 17926 19046 17978
rect 19098 17926 19110 17978
rect 19162 17926 19174 17978
rect 19226 17926 19238 17978
rect 19290 17926 26918 17978
rect 26970 17926 26982 17978
rect 27034 17926 27046 17978
rect 27098 17926 27110 17978
rect 27162 17926 27174 17978
rect 27226 17926 27238 17978
rect 27290 17926 28888 17978
rect 1104 17904 28888 17926
rect 2314 17824 2320 17876
rect 2372 17824 2378 17876
rect 3329 17867 3387 17873
rect 3329 17833 3341 17867
rect 3375 17864 3387 17867
rect 4154 17864 4160 17876
rect 3375 17836 4160 17864
rect 3375 17833 3387 17836
rect 3329 17827 3387 17833
rect 4154 17824 4160 17836
rect 4212 17824 4218 17876
rect 7285 17867 7343 17873
rect 7285 17833 7297 17867
rect 7331 17864 7343 17867
rect 7374 17864 7380 17876
rect 7331 17836 7380 17864
rect 7331 17833 7343 17836
rect 7285 17827 7343 17833
rect 7374 17824 7380 17836
rect 7432 17824 7438 17876
rect 14458 17824 14464 17876
rect 14516 17864 14522 17876
rect 14737 17867 14795 17873
rect 14737 17864 14749 17867
rect 14516 17836 14749 17864
rect 14516 17824 14522 17836
rect 14737 17833 14749 17836
rect 14783 17833 14795 17867
rect 14737 17827 14795 17833
rect 15930 17824 15936 17876
rect 15988 17864 15994 17876
rect 16301 17867 16359 17873
rect 16301 17864 16313 17867
rect 15988 17836 16313 17864
rect 15988 17824 15994 17836
rect 16301 17833 16313 17836
rect 16347 17833 16359 17867
rect 16301 17827 16359 17833
rect 16482 17824 16488 17876
rect 16540 17864 16546 17876
rect 16540 17836 21128 17864
rect 16540 17824 16546 17836
rect 1673 17799 1731 17805
rect 1673 17765 1685 17799
rect 1719 17796 1731 17799
rect 1719 17768 5856 17796
rect 1719 17765 1731 17768
rect 1673 17759 1731 17765
rect 2685 17731 2743 17737
rect 2685 17697 2697 17731
rect 2731 17728 2743 17731
rect 3418 17728 3424 17740
rect 2731 17700 3424 17728
rect 2731 17697 2743 17700
rect 2685 17691 2743 17697
rect 3418 17688 3424 17700
rect 3476 17688 3482 17740
rect 5828 17672 5856 17768
rect 6822 17688 6828 17740
rect 6880 17688 6886 17740
rect 14734 17688 14740 17740
rect 14792 17728 14798 17740
rect 15289 17731 15347 17737
rect 15289 17728 15301 17731
rect 14792 17700 15301 17728
rect 14792 17688 14798 17700
rect 15289 17697 15301 17700
rect 15335 17697 15347 17731
rect 15289 17691 15347 17697
rect 15470 17688 15476 17740
rect 15528 17728 15534 17740
rect 15657 17731 15715 17737
rect 15657 17728 15669 17731
rect 15528 17700 15669 17728
rect 15528 17688 15534 17700
rect 15657 17697 15669 17700
rect 15703 17728 15715 17731
rect 18233 17731 18291 17737
rect 18233 17728 18245 17731
rect 15703 17700 18245 17728
rect 15703 17697 15715 17700
rect 15657 17691 15715 17697
rect 18233 17697 18245 17700
rect 18279 17728 18291 17731
rect 18874 17728 18880 17740
rect 18279 17700 18880 17728
rect 18279 17697 18291 17700
rect 18233 17691 18291 17697
rect 18874 17688 18880 17700
rect 18932 17688 18938 17740
rect 19797 17731 19855 17737
rect 19797 17697 19809 17731
rect 19843 17728 19855 17731
rect 20714 17728 20720 17740
rect 19843 17700 20720 17728
rect 19843 17697 19855 17700
rect 19797 17691 19855 17697
rect 20714 17688 20720 17700
rect 20772 17688 20778 17740
rect 21100 17728 21128 17836
rect 21174 17824 21180 17876
rect 21232 17864 21238 17876
rect 21545 17867 21603 17873
rect 21545 17864 21557 17867
rect 21232 17836 21557 17864
rect 21232 17824 21238 17836
rect 21545 17833 21557 17836
rect 21591 17864 21603 17867
rect 21818 17864 21824 17876
rect 21591 17836 21824 17864
rect 21591 17833 21603 17836
rect 21545 17827 21603 17833
rect 21818 17824 21824 17836
rect 21876 17824 21882 17876
rect 21637 17731 21695 17737
rect 21637 17728 21649 17731
rect 21100 17700 21649 17728
rect 21637 17697 21649 17700
rect 21683 17697 21695 17731
rect 24118 17728 24124 17740
rect 21637 17691 21695 17697
rect 22066 17700 24124 17728
rect 2222 17620 2228 17672
rect 2280 17620 2286 17672
rect 3050 17620 3056 17672
rect 3108 17620 3114 17672
rect 3145 17663 3203 17669
rect 3145 17629 3157 17663
rect 3191 17660 3203 17663
rect 4154 17660 4160 17672
rect 3191 17632 4160 17660
rect 3191 17629 3203 17632
rect 3145 17623 3203 17629
rect 4154 17620 4160 17632
rect 4212 17620 4218 17672
rect 5810 17620 5816 17672
rect 5868 17620 5874 17672
rect 5906 17663 5964 17669
rect 5906 17629 5918 17663
rect 5952 17629 5964 17663
rect 5906 17623 5964 17629
rect 1210 17552 1216 17604
rect 1268 17592 1274 17604
rect 1489 17595 1547 17601
rect 1489 17592 1501 17595
rect 1268 17564 1501 17592
rect 1268 17552 1274 17564
rect 1489 17561 1501 17564
rect 1535 17592 1547 17595
rect 1765 17595 1823 17601
rect 1765 17592 1777 17595
rect 1535 17564 1777 17592
rect 1535 17561 1547 17564
rect 1489 17555 1547 17561
rect 1765 17561 1777 17564
rect 1811 17561 1823 17595
rect 1765 17555 1823 17561
rect 2777 17595 2835 17601
rect 2777 17561 2789 17595
rect 2823 17592 2835 17595
rect 4522 17592 4528 17604
rect 2823 17564 4528 17592
rect 2823 17561 2835 17564
rect 2777 17555 2835 17561
rect 4522 17552 4528 17564
rect 4580 17552 4586 17604
rect 5718 17552 5724 17604
rect 5776 17592 5782 17604
rect 5920 17592 5948 17623
rect 6730 17620 6736 17672
rect 6788 17660 6794 17672
rect 6914 17660 6920 17672
rect 6788 17632 6920 17660
rect 6788 17620 6794 17632
rect 6914 17620 6920 17632
rect 6972 17620 6978 17672
rect 7009 17663 7067 17669
rect 7009 17629 7021 17663
rect 7055 17629 7067 17663
rect 7009 17623 7067 17629
rect 5776 17564 5948 17592
rect 7024 17592 7052 17623
rect 7098 17620 7104 17672
rect 7156 17620 7162 17672
rect 14550 17620 14556 17672
rect 14608 17660 14614 17672
rect 15933 17663 15991 17669
rect 15933 17660 15945 17663
rect 14608 17632 15945 17660
rect 14608 17620 14614 17632
rect 15933 17629 15945 17632
rect 15979 17629 15991 17663
rect 15933 17623 15991 17629
rect 21913 17663 21971 17669
rect 21913 17629 21925 17663
rect 21959 17660 21971 17663
rect 22066 17660 22094 17700
rect 24118 17688 24124 17700
rect 24176 17688 24182 17740
rect 21959 17632 22094 17660
rect 21959 17629 21971 17632
rect 21913 17623 21971 17629
rect 7742 17592 7748 17604
rect 7024 17564 7748 17592
rect 5776 17552 5782 17564
rect 7742 17552 7748 17564
rect 7800 17552 7806 17604
rect 15102 17552 15108 17604
rect 15160 17552 15166 17604
rect 15197 17595 15255 17601
rect 15197 17561 15209 17595
rect 15243 17592 15255 17595
rect 16206 17592 16212 17604
rect 15243 17564 16212 17592
rect 15243 17561 15255 17564
rect 15197 17555 15255 17561
rect 16206 17552 16212 17564
rect 16264 17552 16270 17604
rect 18049 17595 18107 17601
rect 18049 17561 18061 17595
rect 18095 17592 18107 17595
rect 18690 17592 18696 17604
rect 18095 17564 18696 17592
rect 18095 17561 18107 17564
rect 18049 17555 18107 17561
rect 18690 17552 18696 17564
rect 18748 17552 18754 17604
rect 20073 17595 20131 17601
rect 20073 17561 20085 17595
rect 20119 17561 20131 17595
rect 22066 17592 22094 17632
rect 21298 17564 22094 17592
rect 20073 17555 20131 17561
rect 6181 17527 6239 17533
rect 6181 17493 6193 17527
rect 6227 17524 6239 17527
rect 6362 17524 6368 17536
rect 6227 17496 6368 17524
rect 6227 17493 6239 17496
rect 6181 17487 6239 17493
rect 6362 17484 6368 17496
rect 6420 17484 6426 17536
rect 15838 17484 15844 17536
rect 15896 17484 15902 17536
rect 17678 17484 17684 17536
rect 17736 17484 17742 17536
rect 18141 17527 18199 17533
rect 18141 17493 18153 17527
rect 18187 17524 18199 17527
rect 18598 17524 18604 17536
rect 18187 17496 18604 17524
rect 18187 17493 18199 17496
rect 18141 17487 18199 17493
rect 18598 17484 18604 17496
rect 18656 17484 18662 17536
rect 20088 17524 20116 17555
rect 20806 17524 20812 17536
rect 20088 17496 20812 17524
rect 20806 17484 20812 17496
rect 20864 17484 20870 17536
rect 1104 17434 28888 17456
rect 1104 17382 3658 17434
rect 3710 17382 3722 17434
rect 3774 17382 3786 17434
rect 3838 17382 3850 17434
rect 3902 17382 3914 17434
rect 3966 17382 3978 17434
rect 4030 17382 11658 17434
rect 11710 17382 11722 17434
rect 11774 17382 11786 17434
rect 11838 17382 11850 17434
rect 11902 17382 11914 17434
rect 11966 17382 11978 17434
rect 12030 17382 19658 17434
rect 19710 17382 19722 17434
rect 19774 17382 19786 17434
rect 19838 17382 19850 17434
rect 19902 17382 19914 17434
rect 19966 17382 19978 17434
rect 20030 17382 27658 17434
rect 27710 17382 27722 17434
rect 27774 17382 27786 17434
rect 27838 17382 27850 17434
rect 27902 17382 27914 17434
rect 27966 17382 27978 17434
rect 28030 17382 28888 17434
rect 1104 17360 28888 17382
rect 7098 17280 7104 17332
rect 7156 17280 7162 17332
rect 7742 17280 7748 17332
rect 7800 17280 7806 17332
rect 9309 17323 9367 17329
rect 9309 17289 9321 17323
rect 9355 17320 9367 17323
rect 9398 17320 9404 17332
rect 9355 17292 9404 17320
rect 9355 17289 9367 17292
rect 9309 17283 9367 17289
rect 9398 17280 9404 17292
rect 9456 17280 9462 17332
rect 18598 17280 18604 17332
rect 18656 17320 18662 17332
rect 18656 17292 18736 17320
rect 18656 17280 18662 17292
rect 1578 17212 1584 17264
rect 1636 17252 1642 17264
rect 6270 17252 6276 17264
rect 1636 17224 6276 17252
rect 1636 17212 1642 17224
rect 6270 17212 6276 17224
rect 6328 17252 6334 17264
rect 6328 17224 6676 17252
rect 6328 17212 6334 17224
rect 1302 17144 1308 17196
rect 1360 17184 1366 17196
rect 1489 17187 1547 17193
rect 1489 17184 1501 17187
rect 1360 17156 1501 17184
rect 1360 17144 1366 17156
rect 1489 17153 1501 17156
rect 1535 17184 1547 17187
rect 1765 17187 1823 17193
rect 1765 17184 1777 17187
rect 1535 17156 1777 17184
rect 1535 17153 1547 17156
rect 1489 17147 1547 17153
rect 1765 17153 1777 17156
rect 1811 17153 1823 17187
rect 1765 17147 1823 17153
rect 5442 17144 5448 17196
rect 5500 17144 5506 17196
rect 6362 17144 6368 17196
rect 6420 17144 6426 17196
rect 6549 17187 6607 17193
rect 6549 17153 6561 17187
rect 6595 17153 6607 17187
rect 6648 17184 6676 17224
rect 6822 17212 6828 17264
rect 6880 17252 6886 17264
rect 8941 17255 8999 17261
rect 6880 17224 7604 17252
rect 6880 17212 6886 17224
rect 6917 17187 6975 17193
rect 6917 17184 6929 17187
rect 6648 17156 6929 17184
rect 6549 17147 6607 17153
rect 6917 17153 6929 17156
rect 6963 17184 6975 17187
rect 7193 17187 7251 17193
rect 7193 17184 7205 17187
rect 6963 17156 7205 17184
rect 6963 17153 6975 17156
rect 6917 17147 6975 17153
rect 7193 17153 7205 17156
rect 7239 17153 7251 17187
rect 7193 17147 7251 17153
rect 7377 17187 7435 17193
rect 7377 17153 7389 17187
rect 7423 17153 7435 17187
rect 7377 17147 7435 17153
rect 5718 17076 5724 17128
rect 5776 17076 5782 17128
rect 6181 17119 6239 17125
rect 6181 17085 6193 17119
rect 6227 17116 6239 17119
rect 6564 17116 6592 17147
rect 6227 17088 6592 17116
rect 6227 17085 6239 17088
rect 6181 17079 6239 17085
rect 6638 17076 6644 17128
rect 6696 17076 6702 17128
rect 6730 17076 6736 17128
rect 6788 17116 6794 17128
rect 7392 17116 7420 17147
rect 7466 17144 7472 17196
rect 7524 17144 7530 17196
rect 7576 17193 7604 17224
rect 8941 17221 8953 17255
rect 8987 17252 8999 17255
rect 9030 17252 9036 17264
rect 8987 17224 9036 17252
rect 8987 17221 8999 17224
rect 8941 17215 8999 17221
rect 9030 17212 9036 17224
rect 9088 17212 9094 17264
rect 9157 17255 9215 17261
rect 9157 17221 9169 17255
rect 9203 17252 9215 17255
rect 9858 17252 9864 17264
rect 9203 17224 9864 17252
rect 9203 17221 9215 17224
rect 9157 17215 9215 17221
rect 9858 17212 9864 17224
rect 9916 17212 9922 17264
rect 18708 17261 18736 17292
rect 20898 17280 20904 17332
rect 20956 17320 20962 17332
rect 20993 17323 21051 17329
rect 20993 17320 21005 17323
rect 20956 17292 21005 17320
rect 20956 17280 20962 17292
rect 20993 17289 21005 17292
rect 21039 17289 21051 17323
rect 24578 17320 24584 17332
rect 20993 17283 21051 17289
rect 21468 17292 24584 17320
rect 18693 17255 18751 17261
rect 18693 17221 18705 17255
rect 18739 17221 18751 17255
rect 18693 17215 18751 17221
rect 18874 17212 18880 17264
rect 18932 17212 18938 17264
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17184 7619 17187
rect 8386 17184 8392 17196
rect 7607 17156 8392 17184
rect 7607 17153 7619 17156
rect 7561 17147 7619 17153
rect 8386 17144 8392 17156
rect 8444 17144 8450 17196
rect 18230 17144 18236 17196
rect 18288 17144 18294 17196
rect 21174 17144 21180 17196
rect 21232 17144 21238 17196
rect 21468 17193 21496 17292
rect 21818 17212 21824 17264
rect 21876 17252 21882 17264
rect 22005 17255 22063 17261
rect 22005 17252 22017 17255
rect 21876 17224 22017 17252
rect 21876 17212 21882 17224
rect 22005 17221 22017 17224
rect 22051 17221 22063 17255
rect 22005 17215 22063 17221
rect 22388 17193 22416 17292
rect 24578 17280 24584 17292
rect 24636 17280 24642 17332
rect 23014 17252 23020 17264
rect 22848 17224 23020 17252
rect 22848 17193 22876 17224
rect 23014 17212 23020 17224
rect 23072 17212 23078 17264
rect 23106 17212 23112 17264
rect 23164 17212 23170 17264
rect 21453 17187 21511 17193
rect 21453 17153 21465 17187
rect 21499 17153 21511 17187
rect 21453 17147 21511 17153
rect 21637 17187 21695 17193
rect 21637 17153 21649 17187
rect 21683 17153 21695 17187
rect 21637 17147 21695 17153
rect 22373 17187 22431 17193
rect 22373 17153 22385 17187
rect 22419 17153 22431 17187
rect 22373 17147 22431 17153
rect 22833 17187 22891 17193
rect 22833 17153 22845 17187
rect 22879 17153 22891 17187
rect 22833 17147 22891 17153
rect 6788 17088 7420 17116
rect 6788 17076 6794 17088
rect 16850 17076 16856 17128
rect 16908 17076 16914 17128
rect 17129 17119 17187 17125
rect 17129 17085 17141 17119
rect 17175 17116 17187 17119
rect 19061 17119 19119 17125
rect 19061 17116 19073 17119
rect 17175 17088 19073 17116
rect 17175 17085 17187 17088
rect 17129 17079 17187 17085
rect 19061 17085 19073 17088
rect 19107 17085 19119 17119
rect 19061 17079 19119 17085
rect 19886 17076 19892 17128
rect 19944 17116 19950 17128
rect 20622 17116 20628 17128
rect 19944 17088 20628 17116
rect 19944 17076 19950 17088
rect 20622 17076 20628 17088
rect 20680 17116 20686 17128
rect 21652 17116 21680 17147
rect 24210 17144 24216 17196
rect 24268 17144 24274 17196
rect 20680 17088 21680 17116
rect 20680 17076 20686 17088
rect 5810 17008 5816 17060
rect 5868 17048 5874 17060
rect 5997 17051 6055 17057
rect 5997 17048 6009 17051
rect 5868 17020 6009 17048
rect 5868 17008 5874 17020
rect 5997 17017 6009 17020
rect 6043 17048 6055 17051
rect 7834 17048 7840 17060
rect 6043 17020 7840 17048
rect 6043 17017 6055 17020
rect 5997 17011 6055 17017
rect 7834 17008 7840 17020
rect 7892 17008 7898 17060
rect 21821 17051 21879 17057
rect 21821 17017 21833 17051
rect 21867 17048 21879 17051
rect 21867 17020 22692 17048
rect 21867 17017 21879 17020
rect 21821 17011 21879 17017
rect 1581 16983 1639 16989
rect 1581 16949 1593 16983
rect 1627 16980 1639 16983
rect 2590 16980 2596 16992
rect 1627 16952 2596 16980
rect 1627 16949 1639 16952
rect 1581 16943 1639 16949
rect 2590 16940 2596 16952
rect 2648 16940 2654 16992
rect 3602 16940 3608 16992
rect 3660 16980 3666 16992
rect 5537 16983 5595 16989
rect 5537 16980 5549 16983
rect 3660 16952 5549 16980
rect 3660 16940 3666 16952
rect 5537 16949 5549 16952
rect 5583 16980 5595 16983
rect 6822 16980 6828 16992
rect 5583 16952 6828 16980
rect 5583 16949 5595 16952
rect 5537 16943 5595 16949
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 9122 16940 9128 16992
rect 9180 16940 9186 16992
rect 21174 16940 21180 16992
rect 21232 16980 21238 16992
rect 22005 16983 22063 16989
rect 22005 16980 22017 16983
rect 21232 16952 22017 16980
rect 21232 16940 21238 16952
rect 22005 16949 22017 16952
rect 22051 16949 22063 16983
rect 22664 16980 22692 17020
rect 23198 16980 23204 16992
rect 22664 16952 23204 16980
rect 22005 16943 22063 16949
rect 23198 16940 23204 16952
rect 23256 16940 23262 16992
rect 1104 16890 28888 16912
rect 1104 16838 2918 16890
rect 2970 16838 2982 16890
rect 3034 16838 3046 16890
rect 3098 16838 3110 16890
rect 3162 16838 3174 16890
rect 3226 16838 3238 16890
rect 3290 16838 10918 16890
rect 10970 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 11238 16890
rect 11290 16838 18918 16890
rect 18970 16838 18982 16890
rect 19034 16838 19046 16890
rect 19098 16838 19110 16890
rect 19162 16838 19174 16890
rect 19226 16838 19238 16890
rect 19290 16838 26918 16890
rect 26970 16838 26982 16890
rect 27034 16838 27046 16890
rect 27098 16838 27110 16890
rect 27162 16838 27174 16890
rect 27226 16838 27238 16890
rect 27290 16838 28888 16890
rect 1104 16816 28888 16838
rect 2498 16736 2504 16788
rect 2556 16776 2562 16788
rect 2685 16779 2743 16785
rect 2685 16776 2697 16779
rect 2556 16748 2697 16776
rect 2556 16736 2562 16748
rect 2685 16745 2697 16748
rect 2731 16745 2743 16779
rect 2685 16739 2743 16745
rect 6365 16779 6423 16785
rect 6365 16745 6377 16779
rect 6411 16776 6423 16779
rect 6638 16776 6644 16788
rect 6411 16748 6644 16776
rect 6411 16745 6423 16748
rect 6365 16739 6423 16745
rect 6638 16736 6644 16748
rect 6696 16736 6702 16788
rect 6825 16779 6883 16785
rect 6825 16745 6837 16779
rect 6871 16776 6883 16779
rect 7466 16776 7472 16788
rect 6871 16748 7472 16776
rect 6871 16745 6883 16748
rect 6825 16739 6883 16745
rect 1673 16711 1731 16717
rect 1673 16677 1685 16711
rect 1719 16708 1731 16711
rect 1762 16708 1768 16720
rect 1719 16680 1768 16708
rect 1719 16677 1731 16680
rect 1673 16671 1731 16677
rect 1762 16668 1768 16680
rect 1820 16668 1826 16720
rect 2590 16668 2596 16720
rect 2648 16708 2654 16720
rect 6178 16708 6184 16720
rect 2648 16680 6184 16708
rect 2648 16668 2654 16680
rect 6178 16668 6184 16680
rect 6236 16668 6242 16720
rect 6549 16711 6607 16717
rect 6549 16677 6561 16711
rect 6595 16708 6607 16711
rect 6730 16708 6736 16720
rect 6595 16680 6736 16708
rect 6595 16677 6607 16680
rect 6549 16671 6607 16677
rect 6730 16668 6736 16680
rect 6788 16668 6794 16720
rect 6840 16640 6868 16739
rect 7466 16736 7472 16748
rect 7524 16736 7530 16788
rect 8570 16736 8576 16788
rect 8628 16736 8634 16788
rect 11241 16779 11299 16785
rect 11241 16745 11253 16779
rect 11287 16776 11299 16779
rect 12710 16776 12716 16788
rect 11287 16748 12716 16776
rect 11287 16745 11299 16748
rect 11241 16739 11299 16745
rect 12710 16736 12716 16748
rect 12768 16736 12774 16788
rect 17208 16779 17266 16785
rect 17208 16745 17220 16779
rect 17254 16776 17266 16779
rect 17678 16776 17684 16788
rect 17254 16748 17684 16776
rect 17254 16745 17266 16748
rect 17208 16739 17266 16745
rect 17678 16736 17684 16748
rect 17736 16736 17742 16788
rect 18690 16736 18696 16788
rect 18748 16736 18754 16788
rect 23845 16779 23903 16785
rect 23845 16745 23857 16779
rect 23891 16776 23903 16779
rect 23891 16748 24532 16776
rect 23891 16745 23903 16748
rect 23845 16739 23903 16745
rect 20714 16668 20720 16720
rect 20772 16708 20778 16720
rect 23014 16708 23020 16720
rect 20772 16680 23020 16708
rect 20772 16668 20778 16680
rect 23014 16668 23020 16680
rect 23072 16708 23078 16720
rect 23072 16680 24440 16708
rect 23072 16668 23078 16680
rect 6564 16612 6868 16640
rect 6564 16584 6592 16612
rect 8294 16600 8300 16652
rect 8352 16640 8358 16652
rect 9122 16640 9128 16652
rect 8352 16612 9128 16640
rect 8352 16600 8358 16612
rect 9122 16600 9128 16612
rect 9180 16600 9186 16652
rect 11330 16600 11336 16652
rect 11388 16600 11394 16652
rect 11609 16643 11667 16649
rect 11609 16609 11621 16643
rect 11655 16640 11667 16643
rect 12066 16640 12072 16652
rect 11655 16612 12072 16640
rect 11655 16609 11667 16612
rect 11609 16603 11667 16609
rect 12066 16600 12072 16612
rect 12124 16600 12130 16652
rect 16850 16600 16856 16652
rect 16908 16640 16914 16652
rect 16945 16643 17003 16649
rect 16945 16640 16957 16643
rect 16908 16612 16957 16640
rect 16908 16600 16914 16612
rect 16945 16609 16957 16612
rect 16991 16640 17003 16643
rect 17310 16640 17316 16652
rect 16991 16612 17316 16640
rect 16991 16609 17003 16612
rect 16945 16603 17003 16609
rect 17310 16600 17316 16612
rect 17368 16600 17374 16652
rect 22002 16640 22008 16652
rect 19996 16612 22008 16640
rect 2774 16532 2780 16584
rect 2832 16581 2838 16584
rect 2832 16575 2881 16581
rect 2832 16541 2835 16575
rect 2869 16541 2881 16575
rect 2832 16535 2881 16541
rect 3236 16575 3294 16581
rect 3236 16541 3248 16575
rect 3282 16541 3294 16575
rect 3236 16535 3294 16541
rect 3329 16575 3387 16581
rect 3329 16541 3341 16575
rect 3375 16541 3387 16575
rect 3329 16535 3387 16541
rect 2832 16532 2838 16535
rect 1486 16464 1492 16516
rect 1544 16504 1550 16516
rect 1765 16507 1823 16513
rect 1765 16504 1777 16507
rect 1544 16476 1777 16504
rect 1544 16464 1550 16476
rect 1765 16473 1777 16476
rect 1811 16473 1823 16507
rect 1765 16467 1823 16473
rect 2314 16464 2320 16516
rect 2372 16504 2378 16516
rect 2961 16507 3019 16513
rect 2961 16504 2973 16507
rect 2372 16476 2973 16504
rect 2372 16464 2378 16476
rect 2961 16473 2973 16476
rect 3007 16473 3019 16507
rect 2961 16467 3019 16473
rect 3050 16464 3056 16516
rect 3108 16464 3114 16516
rect 3252 16436 3280 16535
rect 3344 16504 3372 16535
rect 3418 16532 3424 16584
rect 3476 16532 3482 16584
rect 3602 16532 3608 16584
rect 3660 16532 3666 16584
rect 5902 16532 5908 16584
rect 5960 16532 5966 16584
rect 6454 16532 6460 16584
rect 6512 16532 6518 16584
rect 6546 16532 6552 16584
rect 6604 16532 6610 16584
rect 6914 16532 6920 16584
rect 6972 16532 6978 16584
rect 7098 16532 7104 16584
rect 7156 16572 7162 16584
rect 7929 16575 7987 16581
rect 7929 16572 7941 16575
rect 7156 16544 7941 16572
rect 7156 16532 7162 16544
rect 7929 16541 7941 16544
rect 7975 16541 7987 16575
rect 7929 16535 7987 16541
rect 8077 16575 8135 16581
rect 8077 16541 8089 16575
rect 8123 16572 8135 16575
rect 8312 16572 8340 16600
rect 8123 16544 8340 16572
rect 8123 16541 8135 16544
rect 8077 16535 8135 16541
rect 8386 16532 8392 16584
rect 8444 16581 8450 16584
rect 8444 16572 8452 16581
rect 8444 16544 8489 16572
rect 8444 16535 8452 16544
rect 8444 16532 8450 16535
rect 12710 16532 12716 16584
rect 12768 16532 12774 16584
rect 19886 16532 19892 16584
rect 19944 16532 19950 16584
rect 19996 16581 20024 16612
rect 22002 16600 22008 16612
rect 22060 16600 22066 16652
rect 23198 16600 23204 16652
rect 23256 16640 23262 16652
rect 24412 16649 24440 16680
rect 23569 16643 23627 16649
rect 23569 16640 23581 16643
rect 23256 16612 23581 16640
rect 23256 16600 23262 16612
rect 23569 16609 23581 16612
rect 23615 16609 23627 16643
rect 23569 16603 23627 16609
rect 24397 16643 24455 16649
rect 24397 16609 24409 16643
rect 24443 16609 24455 16643
rect 24504 16640 24532 16748
rect 24673 16643 24731 16649
rect 24673 16640 24685 16643
rect 24504 16612 24685 16640
rect 24397 16603 24455 16609
rect 24673 16609 24685 16612
rect 24719 16609 24731 16643
rect 24673 16603 24731 16609
rect 19981 16575 20039 16581
rect 19981 16541 19993 16575
rect 20027 16541 20039 16575
rect 19981 16535 20039 16541
rect 23474 16532 23480 16584
rect 23532 16532 23538 16584
rect 3513 16507 3571 16513
rect 3513 16504 3525 16507
rect 3344 16476 3525 16504
rect 3513 16473 3525 16476
rect 3559 16473 3571 16507
rect 3513 16467 3571 16473
rect 6638 16464 6644 16516
rect 6696 16504 6702 16516
rect 6696 16476 6960 16504
rect 6696 16464 6702 16476
rect 3326 16436 3332 16448
rect 3252 16408 3332 16436
rect 3326 16396 3332 16408
rect 3384 16396 3390 16448
rect 6932 16436 6960 16476
rect 8202 16464 8208 16516
rect 8260 16464 8266 16516
rect 8297 16507 8355 16513
rect 8297 16473 8309 16507
rect 8343 16473 8355 16507
rect 8297 16467 8355 16473
rect 8312 16436 8340 16467
rect 18230 16464 18236 16516
rect 18288 16464 18294 16516
rect 6932 16408 8340 16436
rect 12526 16396 12532 16448
rect 12584 16436 12590 16448
rect 13081 16439 13139 16445
rect 13081 16436 13093 16439
rect 12584 16408 13093 16436
rect 12584 16396 12590 16408
rect 13081 16405 13093 16408
rect 13127 16405 13139 16439
rect 23492 16436 23520 16532
rect 24118 16464 24124 16516
rect 24176 16504 24182 16516
rect 24176 16476 25162 16504
rect 24176 16464 24182 16476
rect 26145 16439 26203 16445
rect 26145 16436 26157 16439
rect 23492 16408 26157 16436
rect 13081 16399 13139 16405
rect 26145 16405 26157 16408
rect 26191 16405 26203 16439
rect 26145 16399 26203 16405
rect 1104 16346 28888 16368
rect 1104 16294 3658 16346
rect 3710 16294 3722 16346
rect 3774 16294 3786 16346
rect 3838 16294 3850 16346
rect 3902 16294 3914 16346
rect 3966 16294 3978 16346
rect 4030 16294 11658 16346
rect 11710 16294 11722 16346
rect 11774 16294 11786 16346
rect 11838 16294 11850 16346
rect 11902 16294 11914 16346
rect 11966 16294 11978 16346
rect 12030 16294 19658 16346
rect 19710 16294 19722 16346
rect 19774 16294 19786 16346
rect 19838 16294 19850 16346
rect 19902 16294 19914 16346
rect 19966 16294 19978 16346
rect 20030 16294 27658 16346
rect 27710 16294 27722 16346
rect 27774 16294 27786 16346
rect 27838 16294 27850 16346
rect 27902 16294 27914 16346
rect 27966 16294 27978 16346
rect 28030 16294 28888 16346
rect 1104 16272 28888 16294
rect 1578 16192 1584 16244
rect 1636 16192 1642 16244
rect 2038 16192 2044 16244
rect 2096 16232 2102 16244
rect 2590 16232 2596 16244
rect 2096 16204 2596 16232
rect 2096 16192 2102 16204
rect 2590 16192 2596 16204
rect 2648 16192 2654 16244
rect 2777 16235 2835 16241
rect 2777 16201 2789 16235
rect 2823 16232 2835 16235
rect 3050 16232 3056 16244
rect 2823 16204 3056 16232
rect 2823 16201 2835 16204
rect 2777 16195 2835 16201
rect 3050 16192 3056 16204
rect 3108 16192 3114 16244
rect 3418 16192 3424 16244
rect 3476 16232 3482 16244
rect 3602 16232 3608 16244
rect 3476 16204 3608 16232
rect 3476 16192 3482 16204
rect 3602 16192 3608 16204
rect 3660 16192 3666 16244
rect 6181 16235 6239 16241
rect 6181 16201 6193 16235
rect 6227 16232 6239 16235
rect 6933 16235 6991 16241
rect 6933 16232 6945 16235
rect 6227 16204 6945 16232
rect 6227 16201 6239 16204
rect 6181 16195 6239 16201
rect 6933 16201 6945 16204
rect 6979 16232 6991 16235
rect 6979 16204 7052 16232
rect 6979 16201 6991 16204
rect 6933 16195 6991 16201
rect 2314 16124 2320 16176
rect 2372 16164 2378 16176
rect 5994 16164 6000 16176
rect 2372 16136 3372 16164
rect 2372 16124 2378 16136
rect 1302 16056 1308 16108
rect 1360 16096 1366 16108
rect 1489 16099 1547 16105
rect 1489 16096 1501 16099
rect 1360 16068 1501 16096
rect 1360 16056 1366 16068
rect 1489 16065 1501 16068
rect 1535 16096 1547 16099
rect 1765 16099 1823 16105
rect 1765 16096 1777 16099
rect 1535 16068 1777 16096
rect 1535 16065 1547 16068
rect 1489 16059 1547 16065
rect 1765 16065 1777 16068
rect 1811 16065 1823 16099
rect 1765 16059 1823 16065
rect 2225 16099 2283 16105
rect 2225 16065 2237 16099
rect 2271 16065 2283 16099
rect 2225 16059 2283 16065
rect 2240 16028 2268 16059
rect 2498 16056 2504 16108
rect 2556 16056 2562 16108
rect 2590 16056 2596 16108
rect 2648 16056 2654 16108
rect 2682 16056 2688 16108
rect 2740 16096 2746 16108
rect 3344 16105 3372 16136
rect 5828 16136 6000 16164
rect 2869 16099 2927 16105
rect 2869 16096 2881 16099
rect 2740 16068 2881 16096
rect 2740 16056 2746 16068
rect 2869 16065 2881 16068
rect 2915 16065 2927 16099
rect 2869 16059 2927 16065
rect 3053 16099 3111 16105
rect 3053 16065 3065 16099
rect 3099 16065 3111 16099
rect 3053 16059 3111 16065
rect 3329 16099 3387 16105
rect 3329 16065 3341 16099
rect 3375 16065 3387 16099
rect 3329 16059 3387 16065
rect 3421 16099 3479 16105
rect 3421 16065 3433 16099
rect 3467 16096 3479 16099
rect 3510 16096 3516 16108
rect 3467 16068 3516 16096
rect 3467 16065 3479 16068
rect 3421 16059 3479 16065
rect 3068 16028 3096 16059
rect 3510 16056 3516 16068
rect 3568 16056 3574 16108
rect 3605 16099 3663 16105
rect 3605 16065 3617 16099
rect 3651 16096 3663 16099
rect 4246 16096 4252 16108
rect 3651 16068 4252 16096
rect 3651 16065 3663 16068
rect 3605 16059 3663 16065
rect 4246 16056 4252 16068
rect 4304 16056 4310 16108
rect 5828 16105 5856 16136
rect 5994 16124 6000 16136
rect 6052 16124 6058 16176
rect 6086 16124 6092 16176
rect 6144 16164 6150 16176
rect 6733 16167 6791 16173
rect 6733 16164 6745 16167
rect 6144 16136 6745 16164
rect 6144 16124 6150 16136
rect 6733 16133 6745 16136
rect 6779 16133 6791 16167
rect 6733 16127 6791 16133
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16065 5871 16099
rect 5813 16059 5871 16065
rect 5906 16099 5964 16105
rect 5906 16065 5918 16099
rect 5952 16065 5964 16099
rect 5906 16059 5964 16065
rect 2240 16000 3096 16028
rect 2317 15963 2375 15969
rect 2317 15929 2329 15963
rect 2363 15960 2375 15963
rect 2406 15960 2412 15972
rect 2363 15932 2412 15960
rect 2363 15929 2375 15932
rect 2317 15923 2375 15929
rect 2406 15920 2412 15932
rect 2464 15920 2470 15972
rect 3068 15960 3096 16000
rect 3237 16031 3295 16037
rect 3237 15997 3249 16031
rect 3283 16028 3295 16031
rect 4062 16028 4068 16040
rect 3283 16000 4068 16028
rect 3283 15997 3295 16000
rect 3237 15991 3295 15997
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 3418 15960 3424 15972
rect 3068 15932 3424 15960
rect 3418 15920 3424 15932
rect 3476 15960 3482 15972
rect 3878 15960 3884 15972
rect 3476 15932 3884 15960
rect 3476 15920 3482 15932
rect 3878 15920 3884 15932
rect 3936 15920 3942 15972
rect 2424 15892 2452 15920
rect 5442 15892 5448 15904
rect 2424 15864 5448 15892
rect 5442 15852 5448 15864
rect 5500 15892 5506 15904
rect 5920 15892 5948 16059
rect 5500 15864 5948 15892
rect 5500 15852 5506 15864
rect 6730 15852 6736 15904
rect 6788 15892 6794 15904
rect 6917 15895 6975 15901
rect 6917 15892 6929 15895
rect 6788 15864 6929 15892
rect 6788 15852 6794 15864
rect 6917 15861 6929 15864
rect 6963 15861 6975 15895
rect 7024 15892 7052 16204
rect 7098 16192 7104 16244
rect 7156 16192 7162 16244
rect 8202 16192 8208 16244
rect 8260 16232 8266 16244
rect 9309 16235 9367 16241
rect 9309 16232 9321 16235
rect 8260 16204 9321 16232
rect 8260 16192 8266 16204
rect 9309 16201 9321 16204
rect 9355 16201 9367 16235
rect 9309 16195 9367 16201
rect 9858 16192 9864 16244
rect 9916 16192 9922 16244
rect 9968 16204 10272 16232
rect 7190 16124 7196 16176
rect 7248 16124 7254 16176
rect 7282 16124 7288 16176
rect 7340 16164 7346 16176
rect 7393 16167 7451 16173
rect 7393 16164 7405 16167
rect 7340 16136 7405 16164
rect 7340 16124 7346 16136
rect 7393 16133 7405 16136
rect 7439 16133 7451 16167
rect 7393 16127 7451 16133
rect 9217 16167 9275 16173
rect 9217 16133 9229 16167
rect 9263 16164 9275 16167
rect 9677 16167 9735 16173
rect 9677 16164 9689 16167
rect 9263 16136 9689 16164
rect 9263 16133 9275 16136
rect 9217 16127 9275 16133
rect 9677 16133 9689 16136
rect 9723 16164 9735 16167
rect 9968 16164 9996 16204
rect 9723 16136 9996 16164
rect 10029 16167 10087 16173
rect 9723 16133 9735 16136
rect 9677 16127 9735 16133
rect 10029 16133 10041 16167
rect 10075 16164 10087 16167
rect 10134 16164 10140 16176
rect 10075 16136 10140 16164
rect 10075 16133 10087 16136
rect 10029 16127 10087 16133
rect 10134 16124 10140 16136
rect 10192 16124 10198 16176
rect 10244 16173 10272 16204
rect 12066 16192 12072 16244
rect 12124 16192 12130 16244
rect 12437 16235 12495 16241
rect 12437 16201 12449 16235
rect 12483 16232 12495 16235
rect 12526 16232 12532 16244
rect 12483 16204 12532 16232
rect 12483 16201 12495 16204
rect 12437 16195 12495 16201
rect 12526 16192 12532 16204
rect 12584 16192 12590 16244
rect 16022 16232 16028 16244
rect 12728 16204 16028 16232
rect 10229 16167 10287 16173
rect 10229 16133 10241 16167
rect 10275 16133 10287 16167
rect 10229 16127 10287 16133
rect 8846 16056 8852 16108
rect 8904 16056 8910 16108
rect 8938 16056 8944 16108
rect 8996 16096 9002 16108
rect 9493 16099 9551 16105
rect 8996 16068 9041 16096
rect 8996 16056 9002 16068
rect 9493 16065 9505 16099
rect 9539 16096 9551 16099
rect 9582 16096 9588 16108
rect 9539 16068 9588 16096
rect 9539 16065 9551 16068
rect 9493 16059 9551 16065
rect 9582 16056 9588 16068
rect 9640 16056 9646 16108
rect 9769 16099 9827 16105
rect 9769 16065 9781 16099
rect 9815 16096 9827 16099
rect 11977 16099 12035 16105
rect 9815 16068 10088 16096
rect 9815 16065 9827 16068
rect 9769 16059 9827 16065
rect 7561 15963 7619 15969
rect 7561 15929 7573 15963
rect 7607 15960 7619 15963
rect 8294 15960 8300 15972
rect 7607 15932 8300 15960
rect 7607 15929 7619 15932
rect 7561 15923 7619 15929
rect 8294 15920 8300 15932
rect 8352 15920 8358 15972
rect 10060 15901 10088 16068
rect 11977 16065 11989 16099
rect 12023 16096 12035 16099
rect 12728 16096 12756 16204
rect 16022 16192 16028 16204
rect 16080 16192 16086 16244
rect 14550 16124 14556 16176
rect 14608 16124 14614 16176
rect 14734 16124 14740 16176
rect 14792 16164 14798 16176
rect 14792 16136 18460 16164
rect 14792 16124 14798 16136
rect 18432 16105 18460 16136
rect 12023 16068 12756 16096
rect 12023 16065 12035 16068
rect 11977 16059 12035 16065
rect 12526 15988 12532 16040
rect 12584 15988 12590 16040
rect 12728 16037 12756 16068
rect 18417 16099 18475 16105
rect 18417 16065 18429 16099
rect 18463 16065 18475 16099
rect 18417 16059 18475 16065
rect 18601 16099 18659 16105
rect 18601 16065 18613 16099
rect 18647 16096 18659 16099
rect 18690 16096 18696 16108
rect 18647 16068 18696 16096
rect 18647 16065 18659 16068
rect 18601 16059 18659 16065
rect 18690 16056 18696 16068
rect 18748 16056 18754 16108
rect 12713 16031 12771 16037
rect 12713 15997 12725 16031
rect 12759 15997 12771 16031
rect 12713 15991 12771 15997
rect 15010 15988 15016 16040
rect 15068 15988 15074 16040
rect 15289 16031 15347 16037
rect 15289 16028 15301 16031
rect 15212 16000 15301 16028
rect 15212 15904 15240 16000
rect 15289 15997 15301 16000
rect 15335 15997 15347 16031
rect 15289 15991 15347 15997
rect 7377 15895 7435 15901
rect 7377 15892 7389 15895
rect 7024 15864 7389 15892
rect 6917 15855 6975 15861
rect 7377 15861 7389 15864
rect 7423 15861 7435 15895
rect 7377 15855 7435 15861
rect 10045 15895 10103 15901
rect 10045 15861 10057 15895
rect 10091 15892 10103 15895
rect 10594 15892 10600 15904
rect 10091 15864 10600 15892
rect 10091 15861 10103 15864
rect 10045 15855 10103 15861
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 13538 15852 13544 15904
rect 13596 15852 13602 15904
rect 15194 15852 15200 15904
rect 15252 15852 15258 15904
rect 18782 15852 18788 15904
rect 18840 15852 18846 15904
rect 1104 15802 28888 15824
rect 1104 15750 2918 15802
rect 2970 15750 2982 15802
rect 3034 15750 3046 15802
rect 3098 15750 3110 15802
rect 3162 15750 3174 15802
rect 3226 15750 3238 15802
rect 3290 15750 10918 15802
rect 10970 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 11238 15802
rect 11290 15750 18918 15802
rect 18970 15750 18982 15802
rect 19034 15750 19046 15802
rect 19098 15750 19110 15802
rect 19162 15750 19174 15802
rect 19226 15750 19238 15802
rect 19290 15750 26918 15802
rect 26970 15750 26982 15802
rect 27034 15750 27046 15802
rect 27098 15750 27110 15802
rect 27162 15750 27174 15802
rect 27226 15750 27238 15802
rect 27290 15750 28888 15802
rect 1104 15728 28888 15750
rect 2961 15691 3019 15697
rect 2961 15657 2973 15691
rect 3007 15688 3019 15691
rect 3326 15688 3332 15700
rect 3007 15660 3332 15688
rect 3007 15657 3019 15660
rect 2961 15651 3019 15657
rect 3326 15648 3332 15660
rect 3384 15648 3390 15700
rect 3878 15648 3884 15700
rect 3936 15648 3942 15700
rect 5718 15648 5724 15700
rect 5776 15688 5782 15700
rect 6089 15691 6147 15697
rect 5776 15660 6040 15688
rect 5776 15648 5782 15660
rect 2590 15580 2596 15632
rect 2648 15620 2654 15632
rect 6012 15620 6040 15660
rect 6089 15657 6101 15691
rect 6135 15688 6147 15691
rect 7190 15688 7196 15700
rect 6135 15660 7196 15688
rect 6135 15657 6147 15660
rect 6089 15651 6147 15657
rect 7190 15648 7196 15660
rect 7248 15648 7254 15700
rect 9582 15648 9588 15700
rect 9640 15648 9646 15700
rect 10134 15648 10140 15700
rect 10192 15688 10198 15700
rect 10321 15691 10379 15697
rect 10321 15688 10333 15691
rect 10192 15660 10333 15688
rect 10192 15648 10198 15660
rect 10321 15657 10333 15660
rect 10367 15657 10379 15691
rect 10321 15651 10379 15657
rect 10594 15648 10600 15700
rect 10652 15648 10658 15700
rect 12526 15648 12532 15700
rect 12584 15688 12590 15700
rect 12713 15691 12771 15697
rect 12713 15688 12725 15691
rect 12584 15660 12725 15688
rect 12584 15648 12590 15660
rect 12713 15657 12725 15660
rect 12759 15657 12771 15691
rect 12713 15651 12771 15657
rect 14829 15691 14887 15697
rect 14829 15657 14841 15691
rect 14875 15688 14887 15691
rect 15010 15688 15016 15700
rect 14875 15660 15016 15688
rect 14875 15657 14887 15660
rect 14829 15651 14887 15657
rect 15010 15648 15016 15660
rect 15068 15648 15074 15700
rect 6917 15623 6975 15629
rect 2648 15592 5948 15620
rect 6012 15592 6868 15620
rect 2648 15580 2654 15592
rect 1670 15512 1676 15564
rect 1728 15512 1734 15564
rect 3053 15555 3111 15561
rect 3053 15552 3065 15555
rect 2608 15524 3065 15552
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 2314 15444 2320 15496
rect 2372 15444 2378 15496
rect 2406 15444 2412 15496
rect 2464 15444 2470 15496
rect 2608 15493 2636 15524
rect 3053 15521 3065 15524
rect 3099 15521 3111 15555
rect 3053 15515 3111 15521
rect 2593 15487 2651 15493
rect 2593 15453 2605 15487
rect 2639 15453 2651 15487
rect 2593 15447 2651 15453
rect 2823 15487 2881 15493
rect 2823 15453 2835 15487
rect 2869 15484 2881 15487
rect 3160 15484 3188 15592
rect 5718 15552 5724 15564
rect 2869 15456 3188 15484
rect 3252 15524 5724 15552
rect 2869 15453 2881 15456
rect 2823 15447 2881 15453
rect 2498 15376 2504 15428
rect 2556 15416 2562 15428
rect 2682 15416 2688 15428
rect 2556 15388 2688 15416
rect 2556 15376 2562 15388
rect 2682 15376 2688 15388
rect 2740 15376 2746 15428
rect 1854 15308 1860 15360
rect 1912 15348 1918 15360
rect 3252 15348 3280 15524
rect 3326 15444 3332 15496
rect 3384 15444 3390 15496
rect 3436 15493 3464 15524
rect 5718 15512 5724 15524
rect 5776 15512 5782 15564
rect 5920 15561 5948 15592
rect 5905 15555 5963 15561
rect 5905 15521 5917 15555
rect 5951 15552 5963 15555
rect 6454 15552 6460 15564
rect 5951 15524 6460 15552
rect 5951 15521 5963 15524
rect 5905 15515 5963 15521
rect 6454 15512 6460 15524
rect 6512 15512 6518 15564
rect 6840 15552 6868 15592
rect 6917 15589 6929 15623
rect 6963 15620 6975 15623
rect 7282 15620 7288 15632
rect 6963 15592 7288 15620
rect 6963 15589 6975 15592
rect 6917 15583 6975 15589
rect 7282 15580 7288 15592
rect 7340 15580 7346 15632
rect 8386 15580 8392 15632
rect 8444 15620 8450 15632
rect 8846 15620 8852 15632
rect 8444 15592 8852 15620
rect 8444 15580 8450 15592
rect 8846 15580 8852 15592
rect 8904 15620 8910 15632
rect 9401 15623 9459 15629
rect 9401 15620 9413 15623
rect 8904 15592 9413 15620
rect 8904 15580 8910 15592
rect 9401 15589 9413 15592
rect 9447 15589 9459 15623
rect 9401 15583 9459 15589
rect 8938 15552 8944 15564
rect 6840 15524 8944 15552
rect 8938 15512 8944 15524
rect 8996 15552 9002 15564
rect 9125 15555 9183 15561
rect 9125 15552 9137 15555
rect 8996 15524 9137 15552
rect 8996 15512 9002 15524
rect 9125 15521 9137 15524
rect 9171 15521 9183 15555
rect 9600 15552 9628 15648
rect 14550 15580 14556 15632
rect 14608 15620 14614 15632
rect 15562 15620 15568 15632
rect 14608 15592 15568 15620
rect 14608 15580 14614 15592
rect 15562 15580 15568 15592
rect 15620 15580 15626 15632
rect 13357 15555 13415 15561
rect 9600 15524 10180 15552
rect 9125 15515 9183 15521
rect 3421 15487 3479 15493
rect 3421 15453 3433 15487
rect 3467 15453 3479 15487
rect 3421 15447 3479 15453
rect 3789 15487 3847 15493
rect 3789 15453 3801 15487
rect 3835 15453 3847 15487
rect 3789 15447 3847 15453
rect 5813 15487 5871 15493
rect 5813 15453 5825 15487
rect 5859 15484 5871 15487
rect 6086 15484 6092 15496
rect 5859 15456 6092 15484
rect 5859 15453 5871 15456
rect 5813 15447 5871 15453
rect 3602 15416 3608 15428
rect 3344 15388 3608 15416
rect 3344 15360 3372 15388
rect 3602 15376 3608 15388
rect 3660 15416 3666 15428
rect 3804 15416 3832 15447
rect 6086 15444 6092 15456
rect 6144 15444 6150 15496
rect 6549 15487 6607 15493
rect 6549 15453 6561 15487
rect 6595 15453 6607 15487
rect 6549 15447 6607 15453
rect 3660 15388 3832 15416
rect 3660 15376 3666 15388
rect 5442 15376 5448 15428
rect 5500 15416 5506 15428
rect 6564 15416 6592 15447
rect 6638 15444 6644 15496
rect 6696 15484 6702 15496
rect 9677 15487 9735 15493
rect 6696 15456 6741 15484
rect 6696 15444 6702 15456
rect 9677 15453 9689 15487
rect 9723 15484 9735 15487
rect 9766 15484 9772 15496
rect 9723 15456 9772 15484
rect 9723 15453 9735 15456
rect 9677 15447 9735 15453
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 10152 15493 10180 15524
rect 13357 15521 13369 15555
rect 13403 15552 13415 15555
rect 13630 15552 13636 15564
rect 13403 15524 13636 15552
rect 13403 15521 13415 15524
rect 13357 15515 13415 15521
rect 13630 15512 13636 15524
rect 13688 15512 13694 15564
rect 14277 15555 14335 15561
rect 14277 15521 14289 15555
rect 14323 15552 14335 15555
rect 14734 15552 14740 15564
rect 14323 15524 14740 15552
rect 14323 15521 14335 15524
rect 14277 15515 14335 15521
rect 14734 15512 14740 15524
rect 14792 15512 14798 15564
rect 15194 15512 15200 15564
rect 15252 15552 15258 15564
rect 17037 15555 17095 15561
rect 17037 15552 17049 15555
rect 15252 15524 17049 15552
rect 15252 15512 15258 15524
rect 17037 15521 17049 15524
rect 17083 15552 17095 15555
rect 17310 15552 17316 15564
rect 17083 15524 17316 15552
rect 17083 15521 17095 15524
rect 17037 15515 17095 15521
rect 17310 15512 17316 15524
rect 17368 15512 17374 15564
rect 9861 15487 9919 15493
rect 9861 15453 9873 15487
rect 9907 15453 9919 15487
rect 9861 15447 9919 15453
rect 10137 15487 10195 15493
rect 10137 15453 10149 15487
rect 10183 15453 10195 15487
rect 10137 15447 10195 15453
rect 9876 15416 9904 15447
rect 10410 15444 10416 15496
rect 10468 15444 10474 15496
rect 10506 15487 10564 15493
rect 10506 15453 10518 15487
rect 10552 15453 10564 15487
rect 10506 15447 10564 15453
rect 10520 15416 10548 15447
rect 13078 15444 13084 15496
rect 13136 15484 13142 15496
rect 13538 15484 13544 15496
rect 13136 15456 13544 15484
rect 13136 15444 13142 15456
rect 13538 15444 13544 15456
rect 13596 15484 13602 15496
rect 14461 15487 14519 15493
rect 14461 15484 14473 15487
rect 13596 15456 14473 15484
rect 13596 15444 13602 15456
rect 14461 15453 14473 15456
rect 14507 15453 14519 15487
rect 14461 15447 14519 15453
rect 16945 15487 17003 15493
rect 16945 15453 16957 15487
rect 16991 15484 17003 15487
rect 18785 15487 18843 15493
rect 18785 15484 18797 15487
rect 16991 15456 18797 15484
rect 16991 15453 17003 15456
rect 16945 15447 17003 15453
rect 18785 15453 18797 15456
rect 18831 15484 18843 15487
rect 19334 15484 19340 15496
rect 18831 15456 19340 15484
rect 18831 15453 18843 15456
rect 18785 15447 18843 15453
rect 19334 15444 19340 15456
rect 19392 15484 19398 15496
rect 19981 15487 20039 15493
rect 19981 15484 19993 15487
rect 19392 15456 19993 15484
rect 19392 15444 19398 15456
rect 19981 15453 19993 15456
rect 20027 15484 20039 15487
rect 20165 15487 20223 15493
rect 20165 15484 20177 15487
rect 20027 15456 20177 15484
rect 20027 15453 20039 15456
rect 19981 15447 20039 15453
rect 20165 15453 20177 15456
rect 20211 15453 20223 15487
rect 20165 15447 20223 15453
rect 5500 15388 6592 15416
rect 9646 15388 10548 15416
rect 5500 15376 5506 15388
rect 1912 15320 3280 15348
rect 1912 15308 1918 15320
rect 3326 15308 3332 15360
rect 3384 15308 3390 15360
rect 5902 15308 5908 15360
rect 5960 15348 5966 15360
rect 9646 15348 9674 15388
rect 5960 15320 9674 15348
rect 13173 15351 13231 15357
rect 5960 15308 5966 15320
rect 13173 15317 13185 15351
rect 13219 15348 13231 15351
rect 13262 15348 13268 15360
rect 13219 15320 13268 15348
rect 13219 15317 13231 15320
rect 13173 15311 13231 15317
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 14366 15308 14372 15360
rect 14424 15308 14430 15360
rect 20714 15308 20720 15360
rect 20772 15348 20778 15360
rect 21358 15348 21364 15360
rect 20772 15320 21364 15348
rect 20772 15308 20778 15320
rect 21358 15308 21364 15320
rect 21416 15348 21422 15360
rect 21453 15351 21511 15357
rect 21453 15348 21465 15351
rect 21416 15320 21465 15348
rect 21416 15308 21422 15320
rect 21453 15317 21465 15320
rect 21499 15317 21511 15351
rect 21453 15311 21511 15317
rect 1104 15258 28888 15280
rect 1104 15206 3658 15258
rect 3710 15206 3722 15258
rect 3774 15206 3786 15258
rect 3838 15206 3850 15258
rect 3902 15206 3914 15258
rect 3966 15206 3978 15258
rect 4030 15206 11658 15258
rect 11710 15206 11722 15258
rect 11774 15206 11786 15258
rect 11838 15206 11850 15258
rect 11902 15206 11914 15258
rect 11966 15206 11978 15258
rect 12030 15206 19658 15258
rect 19710 15206 19722 15258
rect 19774 15206 19786 15258
rect 19838 15206 19850 15258
rect 19902 15206 19914 15258
rect 19966 15206 19978 15258
rect 20030 15206 27658 15258
rect 27710 15206 27722 15258
rect 27774 15206 27786 15258
rect 27838 15206 27850 15258
rect 27902 15206 27914 15258
rect 27966 15206 27978 15258
rect 28030 15206 28888 15258
rect 1104 15184 28888 15206
rect 1394 15104 1400 15156
rect 1452 15144 1458 15156
rect 1765 15147 1823 15153
rect 1765 15144 1777 15147
rect 1452 15116 1777 15144
rect 1452 15104 1458 15116
rect 1765 15113 1777 15116
rect 1811 15113 1823 15147
rect 1765 15107 1823 15113
rect 2314 15104 2320 15156
rect 2372 15144 2378 15156
rect 2501 15147 2559 15153
rect 2501 15144 2513 15147
rect 2372 15116 2513 15144
rect 2372 15104 2378 15116
rect 2501 15113 2513 15116
rect 2547 15113 2559 15147
rect 3510 15144 3516 15156
rect 2501 15107 2559 15113
rect 2792 15116 3516 15144
rect 2406 15036 2412 15088
rect 2464 15076 2470 15088
rect 2593 15079 2651 15085
rect 2593 15076 2605 15079
rect 2464 15048 2605 15076
rect 2464 15036 2470 15048
rect 2593 15045 2605 15048
rect 2639 15045 2651 15079
rect 2593 15039 2651 15045
rect 1302 14968 1308 15020
rect 1360 15008 1366 15020
rect 1489 15011 1547 15017
rect 1489 15008 1501 15011
rect 1360 14980 1501 15008
rect 1360 14968 1366 14980
rect 1489 14977 1501 14980
rect 1535 14977 1547 15011
rect 1489 14971 1547 14977
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 2792 15008 2820 15116
rect 3510 15104 3516 15116
rect 3568 15104 3574 15156
rect 9214 15104 9220 15156
rect 9272 15144 9278 15156
rect 9309 15147 9367 15153
rect 9309 15144 9321 15147
rect 9272 15116 9321 15144
rect 9272 15104 9278 15116
rect 9309 15113 9321 15116
rect 9355 15113 9367 15147
rect 9309 15107 9367 15113
rect 9674 15104 9680 15156
rect 9732 15144 9738 15156
rect 9769 15147 9827 15153
rect 9769 15144 9781 15147
rect 9732 15116 9781 15144
rect 9732 15104 9738 15116
rect 9769 15113 9781 15116
rect 9815 15113 9827 15147
rect 9769 15107 9827 15113
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 12713 15147 12771 15153
rect 12713 15144 12725 15147
rect 12676 15116 12725 15144
rect 12676 15104 12682 15116
rect 12713 15113 12725 15116
rect 12759 15113 12771 15147
rect 12713 15107 12771 15113
rect 13078 15104 13084 15156
rect 13136 15104 13142 15156
rect 18782 15104 18788 15156
rect 18840 15144 18846 15156
rect 21545 15147 21603 15153
rect 18840 15116 19196 15144
rect 18840 15104 18846 15116
rect 4430 15076 4436 15088
rect 2884 15048 4436 15076
rect 2884 15017 2912 15048
rect 4430 15036 4436 15048
rect 4488 15036 4494 15088
rect 8018 15036 8024 15088
rect 8076 15076 8082 15088
rect 9401 15079 9459 15085
rect 9401 15076 9413 15079
rect 8076 15048 9413 15076
rect 8076 15036 8082 15048
rect 9401 15045 9413 15048
rect 9447 15045 9459 15079
rect 9401 15039 9459 15045
rect 18414 15036 18420 15088
rect 18472 15076 18478 15088
rect 18969 15079 19027 15085
rect 18969 15076 18981 15079
rect 18472 15048 18981 15076
rect 18472 15036 18478 15048
rect 18969 15045 18981 15048
rect 19015 15045 19027 15079
rect 18969 15039 19027 15045
rect 1719 14980 2820 15008
rect 2868 15011 2926 15017
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 2868 14977 2880 15011
rect 2914 14977 2926 15011
rect 2868 14971 2926 14977
rect 2958 14968 2964 15020
rect 3016 14968 3022 15020
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 15008 3479 15011
rect 6638 15008 6644 15020
rect 3467 14980 6644 15008
rect 3467 14977 3479 14980
rect 3421 14971 3479 14977
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14940 2099 14943
rect 2498 14940 2504 14952
rect 2087 14912 2504 14940
rect 2087 14909 2099 14912
rect 2041 14903 2099 14909
rect 2498 14900 2504 14912
rect 2556 14900 2562 14952
rect 2590 14900 2596 14952
rect 2648 14940 2654 14952
rect 3436 14940 3464 14971
rect 6638 14968 6644 14980
rect 6696 14968 6702 15020
rect 9493 15011 9551 15017
rect 9493 14977 9505 15011
rect 9539 15008 9551 15011
rect 9582 15008 9588 15020
rect 9539 14980 9588 15008
rect 9539 14977 9551 14980
rect 9493 14971 9551 14977
rect 9582 14968 9588 14980
rect 9640 14968 9646 15020
rect 9861 15011 9919 15017
rect 9861 14977 9873 15011
rect 9907 15008 9919 15011
rect 10042 15008 10048 15020
rect 9907 14980 10048 15008
rect 9907 14977 9919 14980
rect 9861 14971 9919 14977
rect 10042 14968 10048 14980
rect 10100 15008 10106 15020
rect 10410 15008 10416 15020
rect 10100 14980 10416 15008
rect 10100 14968 10106 14980
rect 10410 14968 10416 14980
rect 10468 14968 10474 15020
rect 18782 14968 18788 15020
rect 18840 14968 18846 15020
rect 19168 15017 19196 15116
rect 21545 15113 21557 15147
rect 21591 15144 21603 15147
rect 21591 15116 22140 15144
rect 21591 15113 21603 15116
rect 21545 15107 21603 15113
rect 20257 15079 20315 15085
rect 20257 15045 20269 15079
rect 20303 15076 20315 15079
rect 20714 15076 20720 15088
rect 20303 15048 20720 15076
rect 20303 15045 20315 15048
rect 20257 15039 20315 15045
rect 20714 15036 20720 15048
rect 20772 15076 20778 15088
rect 22112 15085 22140 15116
rect 22097 15079 22155 15085
rect 20772 15048 21864 15076
rect 20772 15036 20778 15048
rect 18877 15011 18935 15017
rect 18877 14977 18889 15011
rect 18923 14977 18935 15011
rect 18877 14971 18935 14977
rect 19153 15011 19211 15017
rect 19153 14977 19165 15011
rect 19199 15008 19211 15011
rect 19610 15008 19616 15020
rect 19199 14980 19616 15008
rect 19199 14977 19211 14980
rect 19153 14971 19211 14977
rect 2648 14912 3464 14940
rect 2648 14900 2654 14912
rect 3694 14900 3700 14952
rect 3752 14940 3758 14952
rect 4062 14940 4068 14952
rect 3752 14912 4068 14940
rect 3752 14900 3758 14912
rect 4062 14900 4068 14912
rect 4120 14940 4126 14952
rect 5994 14940 6000 14952
rect 4120 14912 6000 14940
rect 4120 14900 4126 14912
rect 5994 14900 6000 14912
rect 6052 14900 6058 14952
rect 6178 14900 6184 14952
rect 6236 14940 6242 14952
rect 9033 14943 9091 14949
rect 9033 14940 9045 14943
rect 6236 14912 9045 14940
rect 6236 14900 6242 14912
rect 9033 14909 9045 14912
rect 9079 14909 9091 14943
rect 9033 14903 9091 14909
rect 9125 14943 9183 14949
rect 9125 14909 9137 14943
rect 9171 14940 9183 14943
rect 9766 14940 9772 14952
rect 9171 14912 9772 14940
rect 9171 14909 9183 14912
rect 9125 14903 9183 14909
rect 1854 14832 1860 14884
rect 1912 14872 1918 14884
rect 2317 14875 2375 14881
rect 2317 14872 2329 14875
rect 1912 14844 2329 14872
rect 1912 14832 1918 14844
rect 2317 14841 2329 14844
rect 2363 14841 2375 14875
rect 2516 14872 2544 14900
rect 3234 14872 3240 14884
rect 2516 14844 3240 14872
rect 2317 14835 2375 14841
rect 3234 14832 3240 14844
rect 3292 14832 3298 14884
rect 5718 14832 5724 14884
rect 5776 14872 5782 14884
rect 6196 14872 6224 14900
rect 5776 14844 6224 14872
rect 9048 14872 9076 14903
rect 9766 14900 9772 14912
rect 9824 14940 9830 14952
rect 9953 14943 10011 14949
rect 9953 14940 9965 14943
rect 9824 14912 9965 14940
rect 9824 14900 9830 14912
rect 9953 14909 9965 14912
rect 9999 14909 10011 14943
rect 9953 14903 10011 14909
rect 13173 14943 13231 14949
rect 13173 14909 13185 14943
rect 13219 14940 13231 14943
rect 13262 14940 13268 14952
rect 13219 14912 13268 14940
rect 13219 14909 13231 14912
rect 13173 14903 13231 14909
rect 13262 14900 13268 14912
rect 13320 14900 13326 14952
rect 13354 14900 13360 14952
rect 13412 14900 13418 14952
rect 18892 14940 18920 14971
rect 19610 14968 19616 14980
rect 19668 15008 19674 15020
rect 20993 15011 21051 15017
rect 20993 15008 21005 15011
rect 19668 14980 21005 15008
rect 19668 14968 19674 14980
rect 20993 14977 21005 14980
rect 21039 14977 21051 15011
rect 20993 14971 21051 14977
rect 21174 14968 21180 15020
rect 21232 14968 21238 15020
rect 21836 15017 21864 15048
rect 22097 15045 22109 15079
rect 22143 15045 22155 15079
rect 23474 15076 23480 15088
rect 23322 15048 23480 15076
rect 22097 15039 22155 15045
rect 23474 15036 23480 15048
rect 23532 15076 23538 15088
rect 24210 15076 24216 15088
rect 23532 15048 24216 15076
rect 23532 15036 23538 15048
rect 24210 15036 24216 15048
rect 24268 15036 24274 15088
rect 21269 15011 21327 15017
rect 21269 14977 21281 15011
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 21361 15011 21419 15017
rect 21361 14977 21373 15011
rect 21407 14977 21419 15011
rect 21361 14971 21419 14977
rect 21821 15011 21879 15017
rect 21821 14977 21833 15011
rect 21867 14977 21879 15011
rect 21821 14971 21879 14977
rect 20622 14940 20628 14952
rect 18892 14912 20628 14940
rect 20622 14900 20628 14912
rect 20680 14940 20686 14952
rect 21284 14940 21312 14971
rect 20680 14912 21312 14940
rect 20680 14900 20686 14912
rect 9858 14872 9864 14884
rect 9048 14844 9864 14872
rect 5776 14832 5782 14844
rect 9858 14832 9864 14844
rect 9916 14832 9922 14884
rect 17954 14764 17960 14816
rect 18012 14804 18018 14816
rect 18601 14807 18659 14813
rect 18601 14804 18613 14807
rect 18012 14776 18613 14804
rect 18012 14764 18018 14776
rect 18601 14773 18613 14776
rect 18647 14773 18659 14807
rect 21376 14804 21404 14971
rect 21910 14804 21916 14816
rect 21376 14776 21916 14804
rect 18601 14767 18659 14773
rect 21910 14764 21916 14776
rect 21968 14804 21974 14816
rect 23569 14807 23627 14813
rect 23569 14804 23581 14807
rect 21968 14776 23581 14804
rect 21968 14764 21974 14776
rect 23569 14773 23581 14776
rect 23615 14773 23627 14807
rect 23569 14767 23627 14773
rect 1104 14714 28888 14736
rect 1104 14662 2918 14714
rect 2970 14662 2982 14714
rect 3034 14662 3046 14714
rect 3098 14662 3110 14714
rect 3162 14662 3174 14714
rect 3226 14662 3238 14714
rect 3290 14662 10918 14714
rect 10970 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 11238 14714
rect 11290 14662 18918 14714
rect 18970 14662 18982 14714
rect 19034 14662 19046 14714
rect 19098 14662 19110 14714
rect 19162 14662 19174 14714
rect 19226 14662 19238 14714
rect 19290 14662 26918 14714
rect 26970 14662 26982 14714
rect 27034 14662 27046 14714
rect 27098 14662 27110 14714
rect 27162 14662 27174 14714
rect 27226 14662 27238 14714
rect 27290 14662 28888 14714
rect 1104 14640 28888 14662
rect 1302 14560 1308 14612
rect 1360 14600 1366 14612
rect 1673 14603 1731 14609
rect 1673 14600 1685 14603
rect 1360 14572 1685 14600
rect 1360 14560 1366 14572
rect 1673 14569 1685 14572
rect 1719 14569 1731 14603
rect 1673 14563 1731 14569
rect 4246 14560 4252 14612
rect 4304 14560 4310 14612
rect 15838 14560 15844 14612
rect 15896 14600 15902 14612
rect 16117 14603 16175 14609
rect 16117 14600 16129 14603
rect 15896 14572 16129 14600
rect 15896 14560 15902 14572
rect 16117 14569 16129 14572
rect 16163 14569 16175 14603
rect 16117 14563 16175 14569
rect 16206 14560 16212 14612
rect 16264 14560 16270 14612
rect 1581 14535 1639 14541
rect 1581 14501 1593 14535
rect 1627 14532 1639 14535
rect 2590 14532 2596 14544
rect 1627 14504 2596 14532
rect 1627 14501 1639 14504
rect 1581 14495 1639 14501
rect 2590 14492 2596 14504
rect 2648 14492 2654 14544
rect 19245 14535 19303 14541
rect 19245 14501 19257 14535
rect 19291 14501 19303 14535
rect 19245 14495 19303 14501
rect 20916 14504 21496 14532
rect 3694 14464 3700 14476
rect 3344 14436 3700 14464
rect 1302 14356 1308 14408
rect 1360 14396 1366 14408
rect 1397 14399 1455 14405
rect 1397 14396 1409 14399
rect 1360 14368 1409 14396
rect 1360 14356 1366 14368
rect 1397 14365 1409 14368
rect 1443 14396 1455 14399
rect 1857 14399 1915 14405
rect 1857 14396 1869 14399
rect 1443 14368 1869 14396
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 1857 14365 1869 14368
rect 1903 14365 1915 14399
rect 1857 14359 1915 14365
rect 2406 14356 2412 14408
rect 2464 14396 2470 14408
rect 2682 14396 2688 14408
rect 2464 14368 2688 14396
rect 2464 14356 2470 14368
rect 2682 14356 2688 14368
rect 2740 14396 2746 14408
rect 3344 14405 3372 14436
rect 3694 14424 3700 14436
rect 3752 14424 3758 14476
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 15473 14467 15531 14473
rect 15473 14464 15485 14467
rect 15252 14436 15485 14464
rect 15252 14424 15258 14436
rect 15473 14433 15485 14436
rect 15519 14433 15531 14467
rect 15473 14427 15531 14433
rect 16114 14424 16120 14476
rect 16172 14464 16178 14476
rect 16761 14467 16819 14473
rect 16761 14464 16773 14467
rect 16172 14436 16773 14464
rect 16172 14424 16178 14436
rect 16761 14433 16773 14436
rect 16807 14433 16819 14467
rect 16761 14427 16819 14433
rect 17310 14424 17316 14476
rect 17368 14424 17374 14476
rect 17589 14467 17647 14473
rect 17589 14433 17601 14467
rect 17635 14464 17647 14467
rect 19260 14464 19288 14495
rect 17635 14436 19288 14464
rect 17635 14433 17647 14436
rect 17589 14427 17647 14433
rect 19518 14424 19524 14476
rect 19576 14464 19582 14476
rect 19576 14436 19840 14464
rect 19576 14424 19582 14436
rect 2961 14399 3019 14405
rect 2961 14396 2973 14399
rect 2740 14368 2973 14396
rect 2740 14356 2746 14368
rect 2961 14365 2973 14368
rect 3007 14365 3019 14399
rect 2961 14359 3019 14365
rect 3329 14399 3387 14405
rect 3329 14365 3341 14399
rect 3375 14365 3387 14399
rect 3329 14359 3387 14365
rect 3510 14356 3516 14408
rect 3568 14396 3574 14408
rect 3789 14399 3847 14405
rect 3789 14396 3801 14399
rect 3568 14368 3801 14396
rect 3568 14356 3574 14368
rect 3789 14365 3801 14368
rect 3835 14365 3847 14399
rect 3789 14359 3847 14365
rect 4065 14399 4123 14405
rect 4065 14365 4077 14399
rect 4111 14365 4123 14399
rect 4065 14359 4123 14365
rect 3142 14288 3148 14340
rect 3200 14288 3206 14340
rect 3237 14331 3295 14337
rect 3237 14297 3249 14331
rect 3283 14328 3295 14331
rect 3418 14328 3424 14340
rect 3283 14300 3424 14328
rect 3283 14297 3295 14300
rect 3237 14291 3295 14297
rect 3418 14288 3424 14300
rect 3476 14288 3482 14340
rect 4080 14328 4108 14359
rect 18690 14356 18696 14408
rect 18748 14356 18754 14408
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14365 19487 14399
rect 19429 14359 19487 14365
rect 3528 14300 4108 14328
rect 15657 14331 15715 14337
rect 3528 14269 3556 14300
rect 15657 14297 15669 14331
rect 15703 14328 15715 14331
rect 15930 14328 15936 14340
rect 15703 14300 15936 14328
rect 15703 14297 15715 14300
rect 15657 14291 15715 14297
rect 15930 14288 15936 14300
rect 15988 14328 15994 14340
rect 16669 14331 16727 14337
rect 16669 14328 16681 14331
rect 15988 14300 16681 14328
rect 15988 14288 15994 14300
rect 16669 14297 16681 14300
rect 16715 14297 16727 14331
rect 16669 14291 16727 14297
rect 3513 14263 3571 14269
rect 3513 14229 3525 14263
rect 3559 14229 3571 14263
rect 3513 14223 3571 14229
rect 3881 14263 3939 14269
rect 3881 14229 3893 14263
rect 3927 14260 3939 14263
rect 4062 14260 4068 14272
rect 3927 14232 4068 14260
rect 3927 14229 3939 14232
rect 3881 14223 3939 14229
rect 4062 14220 4068 14232
rect 4120 14220 4126 14272
rect 15194 14220 15200 14272
rect 15252 14220 15258 14272
rect 15749 14263 15807 14269
rect 15749 14229 15761 14263
rect 15795 14260 15807 14263
rect 16574 14260 16580 14272
rect 15795 14232 16580 14260
rect 15795 14229 15807 14232
rect 15749 14223 15807 14229
rect 16574 14220 16580 14232
rect 16632 14220 16638 14272
rect 18874 14220 18880 14272
rect 18932 14260 18938 14272
rect 19061 14263 19119 14269
rect 19061 14260 19073 14263
rect 18932 14232 19073 14260
rect 18932 14220 18938 14232
rect 19061 14229 19073 14232
rect 19107 14260 19119 14263
rect 19444 14260 19472 14359
rect 19610 14356 19616 14408
rect 19668 14356 19674 14408
rect 19812 14405 19840 14436
rect 20916 14405 20944 14504
rect 21358 14424 21364 14476
rect 21416 14424 21422 14476
rect 21468 14464 21496 14504
rect 23198 14464 23204 14476
rect 21468 14436 23204 14464
rect 23198 14424 23204 14436
rect 23256 14424 23262 14476
rect 19797 14399 19855 14405
rect 19797 14365 19809 14399
rect 19843 14365 19855 14399
rect 19797 14359 19855 14365
rect 20717 14399 20775 14405
rect 20717 14365 20729 14399
rect 20763 14365 20775 14399
rect 20717 14359 20775 14365
rect 20901 14399 20959 14405
rect 20901 14365 20913 14399
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 19521 14331 19579 14337
rect 19521 14297 19533 14331
rect 19567 14297 19579 14331
rect 19628 14328 19656 14356
rect 20732 14328 20760 14359
rect 21082 14356 21088 14408
rect 21140 14356 21146 14408
rect 19628 14300 20760 14328
rect 20993 14331 21051 14337
rect 19521 14291 19579 14297
rect 20993 14297 21005 14331
rect 21039 14297 21051 14331
rect 20993 14291 21051 14297
rect 21637 14331 21695 14337
rect 21637 14297 21649 14331
rect 21683 14297 21695 14331
rect 23474 14328 23480 14340
rect 22862 14300 23480 14328
rect 21637 14291 21695 14297
rect 19107 14232 19472 14260
rect 19536 14260 19564 14291
rect 20622 14260 20628 14272
rect 19536 14232 20628 14260
rect 19107 14229 19119 14232
rect 19061 14223 19119 14229
rect 20622 14220 20628 14232
rect 20680 14260 20686 14272
rect 21008 14260 21036 14291
rect 20680 14232 21036 14260
rect 21269 14263 21327 14269
rect 20680 14220 20686 14232
rect 21269 14229 21281 14263
rect 21315 14260 21327 14263
rect 21652 14260 21680 14291
rect 23474 14288 23480 14300
rect 23532 14288 23538 14340
rect 21315 14232 21680 14260
rect 21315 14229 21327 14232
rect 21269 14223 21327 14229
rect 23106 14220 23112 14272
rect 23164 14220 23170 14272
rect 1104 14170 28888 14192
rect 1104 14118 3658 14170
rect 3710 14118 3722 14170
rect 3774 14118 3786 14170
rect 3838 14118 3850 14170
rect 3902 14118 3914 14170
rect 3966 14118 3978 14170
rect 4030 14118 11658 14170
rect 11710 14118 11722 14170
rect 11774 14118 11786 14170
rect 11838 14118 11850 14170
rect 11902 14118 11914 14170
rect 11966 14118 11978 14170
rect 12030 14118 19658 14170
rect 19710 14118 19722 14170
rect 19774 14118 19786 14170
rect 19838 14118 19850 14170
rect 19902 14118 19914 14170
rect 19966 14118 19978 14170
rect 20030 14118 27658 14170
rect 27710 14118 27722 14170
rect 27774 14118 27786 14170
rect 27838 14118 27850 14170
rect 27902 14118 27914 14170
rect 27966 14118 27978 14170
rect 28030 14118 28888 14170
rect 1104 14096 28888 14118
rect 3510 14016 3516 14068
rect 3568 14016 3574 14068
rect 3605 14059 3663 14065
rect 3605 14025 3617 14059
rect 3651 14056 3663 14059
rect 4062 14056 4068 14068
rect 3651 14028 4068 14056
rect 3651 14025 3663 14028
rect 3605 14019 3663 14025
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 8389 14059 8447 14065
rect 6656 14028 8248 14056
rect 1673 13991 1731 13997
rect 1673 13957 1685 13991
rect 1719 13988 1731 13991
rect 3142 13988 3148 14000
rect 1719 13960 3148 13988
rect 1719 13957 1731 13960
rect 1673 13951 1731 13957
rect 3142 13948 3148 13960
rect 3200 13988 3206 14000
rect 3200 13960 3372 13988
rect 3200 13948 3206 13960
rect 1302 13880 1308 13932
rect 1360 13920 1366 13932
rect 1489 13923 1547 13929
rect 1489 13920 1501 13923
rect 1360 13892 1501 13920
rect 1360 13880 1366 13892
rect 1489 13889 1501 13892
rect 1535 13920 1547 13923
rect 1765 13923 1823 13929
rect 1765 13920 1777 13923
rect 1535 13892 1777 13920
rect 1535 13889 1547 13892
rect 1489 13883 1547 13889
rect 1765 13889 1777 13892
rect 1811 13889 1823 13923
rect 1765 13883 1823 13889
rect 2958 13880 2964 13932
rect 3016 13880 3022 13932
rect 3344 13929 3372 13960
rect 4080 13960 5948 13988
rect 3237 13923 3295 13929
rect 3237 13889 3249 13923
rect 3283 13889 3295 13923
rect 3237 13883 3295 13889
rect 3329 13923 3387 13929
rect 3329 13889 3341 13923
rect 3375 13889 3387 13923
rect 3329 13883 3387 13889
rect 3252 13852 3280 13883
rect 2746 13824 3280 13852
rect 3344 13852 3372 13883
rect 3786 13880 3792 13932
rect 3844 13880 3850 13932
rect 3878 13880 3884 13932
rect 3936 13880 3942 13932
rect 3970 13880 3976 13932
rect 4028 13920 4034 13932
rect 4080 13929 4108 13960
rect 4065 13923 4123 13929
rect 4065 13920 4077 13923
rect 4028 13892 4077 13920
rect 4028 13880 4034 13892
rect 4065 13889 4077 13892
rect 4111 13889 4123 13923
rect 4065 13883 4123 13889
rect 4154 13880 4160 13932
rect 4212 13880 4218 13932
rect 5920 13920 5948 13960
rect 5994 13948 6000 14000
rect 6052 13988 6058 14000
rect 6656 13988 6684 14028
rect 6052 13960 6684 13988
rect 6052 13948 6058 13960
rect 5920 13892 6408 13920
rect 6086 13852 6092 13864
rect 3344 13824 6092 13852
rect 2406 13744 2412 13796
rect 2464 13784 2470 13796
rect 2746 13784 2774 13824
rect 6086 13812 6092 13824
rect 6144 13812 6150 13864
rect 6380 13852 6408 13892
rect 6454 13880 6460 13932
rect 6512 13880 6518 13932
rect 6656 13929 6684 13960
rect 8018 13948 8024 14000
rect 8076 13948 8082 14000
rect 6611 13923 6684 13929
rect 6611 13889 6623 13923
rect 6657 13892 6684 13923
rect 6657 13889 6669 13892
rect 6611 13883 6669 13889
rect 7006 13880 7012 13932
rect 7064 13920 7070 13932
rect 7745 13923 7803 13929
rect 7745 13920 7757 13923
rect 7064 13892 7757 13920
rect 7064 13880 7070 13892
rect 7745 13889 7757 13892
rect 7791 13889 7803 13923
rect 7745 13883 7803 13889
rect 7893 13923 7951 13929
rect 7893 13889 7905 13923
rect 7939 13920 7951 13923
rect 7939 13889 7972 13920
rect 7893 13883 7972 13889
rect 7944 13852 7972 13883
rect 8110 13880 8116 13932
rect 8168 13880 8174 13932
rect 8220 13929 8248 14028
rect 8389 14025 8401 14059
rect 8435 14056 8447 14059
rect 8478 14056 8484 14068
rect 8435 14028 8484 14056
rect 8435 14025 8447 14028
rect 8389 14019 8447 14025
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 9582 14016 9588 14068
rect 9640 14016 9646 14068
rect 11977 14059 12035 14065
rect 11977 14025 11989 14059
rect 12023 14056 12035 14059
rect 12158 14056 12164 14068
rect 12023 14028 12164 14056
rect 12023 14025 12035 14028
rect 11977 14019 12035 14025
rect 12158 14016 12164 14028
rect 12216 14016 12222 14068
rect 15102 14056 15108 14068
rect 14752 14028 15108 14056
rect 14752 14000 14780 14028
rect 15102 14016 15108 14028
rect 15160 14016 15166 14068
rect 18782 14016 18788 14068
rect 18840 14056 18846 14068
rect 19429 14059 19487 14065
rect 19429 14056 19441 14059
rect 18840 14028 19441 14056
rect 18840 14016 18846 14028
rect 19429 14025 19441 14028
rect 19475 14025 19487 14059
rect 19429 14019 19487 14025
rect 21913 14059 21971 14065
rect 21913 14025 21925 14059
rect 21959 14056 21971 14059
rect 22278 14056 22284 14068
rect 21959 14028 22284 14056
rect 21959 14025 21971 14028
rect 21913 14019 21971 14025
rect 22278 14016 22284 14028
rect 22336 14016 22342 14068
rect 22370 14016 22376 14068
rect 22428 14056 22434 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 22428 14028 23397 14056
rect 22428 14016 22434 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 23385 14019 23443 14025
rect 9214 13948 9220 14000
rect 9272 13948 9278 14000
rect 9490 13997 9496 14000
rect 9433 13991 9496 13997
rect 9433 13957 9445 13991
rect 9479 13957 9496 13991
rect 9433 13951 9496 13957
rect 9490 13948 9496 13951
rect 9548 13948 9554 14000
rect 14734 13988 14740 14000
rect 14200 13960 14740 13988
rect 8210 13923 8268 13929
rect 8210 13889 8222 13923
rect 8256 13889 8268 13923
rect 8210 13883 8268 13889
rect 12437 13923 12495 13929
rect 12437 13889 12449 13923
rect 12483 13920 12495 13923
rect 13262 13920 13268 13932
rect 12483 13892 13268 13920
rect 12483 13889 12495 13892
rect 12437 13883 12495 13889
rect 13262 13880 13268 13892
rect 13320 13880 13326 13932
rect 14200 13929 14228 13960
rect 14734 13948 14740 13960
rect 14792 13948 14798 14000
rect 17954 13948 17960 14000
rect 18012 13948 18018 14000
rect 18506 13948 18512 14000
rect 18564 13948 18570 14000
rect 21358 13948 21364 14000
rect 21416 13988 21422 14000
rect 21416 13960 23980 13988
rect 21416 13948 21422 13960
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 15562 13880 15568 13932
rect 15620 13920 15626 13932
rect 15620 13892 16988 13920
rect 15620 13880 15626 13892
rect 8938 13852 8944 13864
rect 6380 13824 7880 13852
rect 7944 13824 8944 13852
rect 3326 13784 3332 13796
rect 2464 13756 2774 13784
rect 2976 13756 3332 13784
rect 2464 13744 2470 13756
rect 2590 13676 2596 13728
rect 2648 13716 2654 13728
rect 2976 13716 3004 13756
rect 3326 13744 3332 13756
rect 3384 13744 3390 13796
rect 6825 13787 6883 13793
rect 6825 13753 6837 13787
rect 6871 13784 6883 13787
rect 7098 13784 7104 13796
rect 6871 13756 7104 13784
rect 6871 13753 6883 13756
rect 6825 13747 6883 13753
rect 7098 13744 7104 13756
rect 7156 13744 7162 13796
rect 7852 13784 7880 13824
rect 8938 13812 8944 13824
rect 8996 13812 9002 13864
rect 10042 13852 10048 13864
rect 9048 13824 10048 13852
rect 9048 13784 9076 13824
rect 10042 13812 10048 13824
rect 10100 13812 10106 13864
rect 12526 13812 12532 13864
rect 12584 13812 12590 13864
rect 12621 13855 12679 13861
rect 12621 13821 12633 13855
rect 12667 13821 12679 13855
rect 12621 13815 12679 13821
rect 7852 13756 9076 13784
rect 12158 13744 12164 13796
rect 12216 13784 12222 13796
rect 12636 13784 12664 13815
rect 14458 13812 14464 13864
rect 14516 13812 14522 13864
rect 15930 13812 15936 13864
rect 15988 13812 15994 13864
rect 16114 13812 16120 13864
rect 16172 13812 16178 13864
rect 16960 13852 16988 13892
rect 17310 13880 17316 13932
rect 17368 13920 17374 13932
rect 17681 13923 17739 13929
rect 17681 13920 17693 13923
rect 17368 13892 17693 13920
rect 17368 13880 17374 13892
rect 17681 13889 17693 13892
rect 17727 13889 17739 13923
rect 17681 13883 17739 13889
rect 21082 13880 21088 13932
rect 21140 13920 21146 13932
rect 22281 13923 22339 13929
rect 22281 13920 22293 13923
rect 21140 13892 22293 13920
rect 21140 13880 21146 13892
rect 22281 13889 22293 13892
rect 22327 13920 22339 13923
rect 23106 13920 23112 13932
rect 22327 13892 23112 13920
rect 22327 13889 22339 13892
rect 22281 13883 22339 13889
rect 23106 13880 23112 13892
rect 23164 13920 23170 13932
rect 23952 13929 23980 13960
rect 24210 13948 24216 14000
rect 24268 13988 24274 14000
rect 24670 13988 24676 14000
rect 24268 13960 24676 13988
rect 24268 13948 24274 13960
rect 24670 13948 24676 13960
rect 24728 13948 24734 14000
rect 23477 13923 23535 13929
rect 23477 13920 23489 13923
rect 23164 13892 23489 13920
rect 23164 13880 23170 13892
rect 23477 13889 23489 13892
rect 23523 13889 23535 13923
rect 23477 13883 23535 13889
rect 23937 13923 23995 13929
rect 23937 13889 23949 13923
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 18506 13852 18512 13864
rect 16960 13824 18512 13852
rect 18506 13812 18512 13824
rect 18564 13812 18570 13864
rect 21910 13812 21916 13864
rect 21968 13852 21974 13864
rect 22370 13852 22376 13864
rect 21968 13824 22376 13852
rect 21968 13812 21974 13824
rect 22370 13812 22376 13824
rect 22428 13812 22434 13864
rect 22465 13855 22523 13861
rect 22465 13821 22477 13855
rect 22511 13821 22523 13855
rect 22465 13815 22523 13821
rect 12216 13756 12664 13784
rect 12216 13744 12222 13756
rect 2648 13688 3004 13716
rect 2648 13676 2654 13688
rect 3050 13676 3056 13728
rect 3108 13716 3114 13728
rect 3786 13716 3792 13728
rect 3108 13688 3792 13716
rect 3108 13676 3114 13688
rect 3786 13676 3792 13688
rect 3844 13716 3850 13728
rect 8386 13716 8392 13728
rect 3844 13688 8392 13716
rect 3844 13676 3850 13688
rect 8386 13676 8392 13688
rect 8444 13676 8450 13728
rect 9398 13676 9404 13728
rect 9456 13676 9462 13728
rect 12066 13676 12072 13728
rect 12124 13676 12130 13728
rect 22480 13716 22508 13815
rect 23198 13812 23204 13864
rect 23256 13812 23262 13864
rect 24210 13812 24216 13864
rect 24268 13812 24274 13864
rect 24762 13812 24768 13864
rect 24820 13852 24826 13864
rect 25685 13855 25743 13861
rect 25685 13852 25697 13855
rect 24820 13824 25697 13852
rect 24820 13812 24826 13824
rect 25685 13821 25697 13824
rect 25731 13821 25743 13855
rect 25685 13815 25743 13821
rect 23658 13716 23664 13728
rect 22480 13688 23664 13716
rect 23658 13676 23664 13688
rect 23716 13676 23722 13728
rect 23842 13676 23848 13728
rect 23900 13676 23906 13728
rect 1104 13626 28888 13648
rect 1104 13574 2918 13626
rect 2970 13574 2982 13626
rect 3034 13574 3046 13626
rect 3098 13574 3110 13626
rect 3162 13574 3174 13626
rect 3226 13574 3238 13626
rect 3290 13574 10918 13626
rect 10970 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 11238 13626
rect 11290 13574 18918 13626
rect 18970 13574 18982 13626
rect 19034 13574 19046 13626
rect 19098 13574 19110 13626
rect 19162 13574 19174 13626
rect 19226 13574 19238 13626
rect 19290 13574 26918 13626
rect 26970 13574 26982 13626
rect 27034 13574 27046 13626
rect 27098 13574 27110 13626
rect 27162 13574 27174 13626
rect 27226 13574 27238 13626
rect 27290 13574 28888 13626
rect 1104 13552 28888 13574
rect 3510 13472 3516 13524
rect 3568 13472 3574 13524
rect 4154 13472 4160 13524
rect 4212 13512 4218 13524
rect 4525 13515 4583 13521
rect 4525 13512 4537 13515
rect 4212 13484 4537 13512
rect 4212 13472 4218 13484
rect 4525 13481 4537 13484
rect 4571 13481 4583 13515
rect 4525 13475 4583 13481
rect 6086 13472 6092 13524
rect 6144 13512 6150 13524
rect 6454 13512 6460 13524
rect 6144 13484 6460 13512
rect 6144 13472 6150 13484
rect 6454 13472 6460 13484
rect 6512 13512 6518 13524
rect 6825 13515 6883 13521
rect 6825 13512 6837 13515
rect 6512 13484 6837 13512
rect 6512 13472 6518 13484
rect 6825 13481 6837 13484
rect 6871 13481 6883 13515
rect 6825 13475 6883 13481
rect 7006 13472 7012 13524
rect 7064 13472 7070 13524
rect 7285 13515 7343 13521
rect 7285 13481 7297 13515
rect 7331 13481 7343 13515
rect 7285 13475 7343 13481
rect 7653 13515 7711 13521
rect 7653 13481 7665 13515
rect 7699 13512 7711 13515
rect 8110 13512 8116 13524
rect 7699 13484 8116 13512
rect 7699 13481 7711 13484
rect 7653 13475 7711 13481
rect 2866 13404 2872 13456
rect 2924 13444 2930 13456
rect 3970 13444 3976 13456
rect 2924 13416 3976 13444
rect 2924 13404 2930 13416
rect 3970 13404 3976 13416
rect 4028 13404 4034 13456
rect 7300 13444 7328 13475
rect 8110 13472 8116 13484
rect 8168 13472 8174 13524
rect 8938 13472 8944 13524
rect 8996 13472 9002 13524
rect 14458 13472 14464 13524
rect 14516 13472 14522 13524
rect 24210 13472 24216 13524
rect 24268 13512 24274 13524
rect 24397 13515 24455 13521
rect 24397 13512 24409 13515
rect 24268 13484 24409 13512
rect 24268 13472 24274 13484
rect 24397 13481 24409 13484
rect 24443 13481 24455 13515
rect 24397 13475 24455 13481
rect 6840 13416 7328 13444
rect 7469 13447 7527 13453
rect 1673 13379 1731 13385
rect 1673 13345 1685 13379
rect 1719 13376 1731 13379
rect 2774 13376 2780 13388
rect 1719 13348 2780 13376
rect 1719 13345 1731 13348
rect 1673 13339 1731 13345
rect 2774 13336 2780 13348
rect 2832 13336 2838 13388
rect 3510 13336 3516 13388
rect 3568 13376 3574 13388
rect 4065 13379 4123 13385
rect 4065 13376 4077 13379
rect 3568 13348 4077 13376
rect 3568 13336 3574 13348
rect 4065 13345 4077 13348
rect 4111 13345 4123 13379
rect 4065 13339 4123 13345
rect 4246 13336 4252 13388
rect 4304 13336 4310 13388
rect 6270 13336 6276 13388
rect 6328 13376 6334 13388
rect 6457 13379 6515 13385
rect 6457 13376 6469 13379
rect 6328 13348 6469 13376
rect 6328 13336 6334 13348
rect 6457 13345 6469 13348
rect 6503 13345 6515 13379
rect 6457 13339 6515 13345
rect 1210 13268 1216 13320
rect 1268 13308 1274 13320
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 1268 13280 1409 13308
rect 1268 13268 1274 13280
rect 1397 13277 1409 13280
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 2498 13268 2504 13320
rect 2556 13308 2562 13320
rect 3234 13308 3240 13320
rect 2556 13280 3240 13308
rect 2556 13268 2562 13280
rect 3234 13268 3240 13280
rect 3292 13308 3298 13320
rect 3605 13311 3663 13317
rect 3605 13308 3617 13311
rect 3292 13280 3617 13308
rect 3292 13268 3298 13280
rect 3605 13277 3617 13280
rect 3651 13277 3663 13311
rect 3605 13271 3663 13277
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13277 4031 13311
rect 3973 13271 4031 13277
rect 4157 13311 4215 13317
rect 4157 13277 4169 13311
rect 4203 13277 4215 13311
rect 4157 13271 4215 13277
rect 3418 13200 3424 13252
rect 3476 13240 3482 13252
rect 3988 13240 4016 13271
rect 3476 13212 4016 13240
rect 3476 13200 3482 13212
rect 4062 13200 4068 13252
rect 4120 13240 4126 13252
rect 4172 13240 4200 13271
rect 4430 13268 4436 13320
rect 4488 13268 4494 13320
rect 5994 13268 6000 13320
rect 6052 13268 6058 13320
rect 6151 13311 6209 13317
rect 6151 13277 6163 13311
rect 6197 13308 6209 13311
rect 6546 13308 6552 13320
rect 6197 13280 6552 13308
rect 6197 13277 6209 13280
rect 6151 13271 6209 13277
rect 6546 13268 6552 13280
rect 6604 13268 6610 13320
rect 6840 13249 6868 13416
rect 7469 13413 7481 13447
rect 7515 13444 7527 13447
rect 8018 13444 8024 13456
rect 7515 13416 8024 13444
rect 7515 13413 7527 13416
rect 7469 13407 7527 13413
rect 8018 13404 8024 13416
rect 8076 13404 8082 13456
rect 14826 13404 14832 13456
rect 14884 13444 14890 13456
rect 14884 13416 15056 13444
rect 14884 13404 14890 13416
rect 6914 13336 6920 13388
rect 6972 13376 6978 13388
rect 7834 13376 7840 13388
rect 6972 13348 7840 13376
rect 6972 13336 6978 13348
rect 7834 13336 7840 13348
rect 7892 13376 7898 13388
rect 8757 13379 8815 13385
rect 7892 13348 8524 13376
rect 7892 13336 7898 13348
rect 7561 13311 7619 13317
rect 7561 13308 7573 13311
rect 6932 13280 7573 13308
rect 4120 13212 4200 13240
rect 6365 13243 6423 13249
rect 4120 13200 4126 13212
rect 6365 13209 6377 13243
rect 6411 13240 6423 13243
rect 6825 13243 6883 13249
rect 6825 13240 6837 13243
rect 6411 13212 6837 13240
rect 6411 13209 6423 13212
rect 6365 13203 6423 13209
rect 6825 13209 6837 13212
rect 6871 13209 6883 13243
rect 6825 13203 6883 13209
rect 3789 13175 3847 13181
rect 3789 13141 3801 13175
rect 3835 13172 3847 13175
rect 4522 13172 4528 13184
rect 3835 13144 4528 13172
rect 3835 13141 3847 13144
rect 3789 13135 3847 13141
rect 4522 13132 4528 13144
rect 4580 13132 4586 13184
rect 6546 13132 6552 13184
rect 6604 13172 6610 13184
rect 6932 13172 6960 13280
rect 7561 13277 7573 13280
rect 7607 13277 7619 13311
rect 7561 13271 7619 13277
rect 8386 13268 8392 13320
rect 8444 13268 8450 13320
rect 8496 13317 8524 13348
rect 8757 13345 8769 13379
rect 8803 13376 8815 13379
rect 9217 13379 9275 13385
rect 9217 13376 9229 13379
rect 8803 13348 9229 13376
rect 8803 13345 8815 13348
rect 8757 13339 8815 13345
rect 9217 13345 9229 13348
rect 9263 13376 9275 13379
rect 9398 13376 9404 13388
rect 9263 13348 9404 13376
rect 9263 13345 9275 13348
rect 9217 13339 9275 13345
rect 9398 13336 9404 13348
rect 9456 13336 9462 13388
rect 15028 13385 15056 13416
rect 24486 13404 24492 13456
rect 24544 13444 24550 13456
rect 24544 13416 24992 13444
rect 24544 13404 24550 13416
rect 15013 13379 15071 13385
rect 15013 13345 15025 13379
rect 15059 13345 15071 13379
rect 15013 13339 15071 13345
rect 23842 13336 23848 13388
rect 23900 13376 23906 13388
rect 24964 13385 24992 13416
rect 24857 13379 24915 13385
rect 24857 13376 24869 13379
rect 23900 13348 24869 13376
rect 23900 13336 23906 13348
rect 24857 13345 24869 13348
rect 24903 13345 24915 13379
rect 24857 13339 24915 13345
rect 24949 13379 25007 13385
rect 24949 13345 24961 13379
rect 24995 13345 25007 13379
rect 24949 13339 25007 13345
rect 8482 13311 8540 13317
rect 8482 13277 8494 13311
rect 8528 13308 8540 13311
rect 8846 13308 8852 13320
rect 8528 13280 8852 13308
rect 8528 13277 8540 13280
rect 8482 13271 8540 13277
rect 8846 13268 8852 13280
rect 8904 13268 8910 13320
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13308 9183 13311
rect 9490 13308 9496 13320
rect 9171 13280 9496 13308
rect 9171 13277 9183 13280
rect 9125 13271 9183 13277
rect 9490 13268 9496 13280
rect 9548 13308 9554 13320
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 9548 13280 9689 13308
rect 9548 13268 9554 13280
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 9858 13268 9864 13320
rect 9916 13317 9922 13320
rect 9916 13311 9949 13317
rect 9937 13277 9949 13311
rect 9916 13271 9949 13277
rect 9916 13268 9922 13271
rect 10042 13268 10048 13320
rect 10100 13268 10106 13320
rect 11330 13268 11336 13320
rect 11388 13308 11394 13320
rect 12989 13311 13047 13317
rect 12989 13308 13001 13311
rect 11388 13280 13001 13308
rect 11388 13268 11394 13280
rect 12989 13277 13001 13280
rect 13035 13277 13047 13311
rect 12989 13271 13047 13277
rect 14829 13311 14887 13317
rect 14829 13277 14841 13311
rect 14875 13308 14887 13311
rect 15930 13308 15936 13320
rect 14875 13280 15936 13308
rect 14875 13277 14887 13280
rect 14829 13271 14887 13277
rect 15930 13268 15936 13280
rect 15988 13268 15994 13320
rect 24762 13268 24768 13320
rect 24820 13268 24826 13320
rect 7098 13200 7104 13252
rect 7156 13200 7162 13252
rect 11425 13243 11483 13249
rect 11425 13209 11437 13243
rect 11471 13240 11483 13243
rect 11514 13240 11520 13252
rect 11471 13212 11520 13240
rect 11471 13209 11483 13212
rect 11425 13203 11483 13209
rect 11514 13200 11520 13212
rect 11572 13240 11578 13252
rect 13265 13243 13323 13249
rect 13265 13240 13277 13243
rect 11572 13212 13277 13240
rect 11572 13200 11578 13212
rect 13265 13209 13277 13212
rect 13311 13209 13323 13243
rect 13265 13203 13323 13209
rect 13814 13200 13820 13252
rect 13872 13240 13878 13252
rect 14921 13243 14979 13249
rect 14921 13240 14933 13243
rect 13872 13212 14933 13240
rect 13872 13200 13878 13212
rect 14921 13209 14933 13212
rect 14967 13209 14979 13243
rect 14921 13203 14979 13209
rect 6604 13144 6960 13172
rect 6604 13132 6610 13144
rect 7190 13132 7196 13184
rect 7248 13172 7254 13184
rect 7301 13175 7359 13181
rect 7301 13172 7313 13175
rect 7248 13144 7313 13172
rect 7248 13132 7254 13144
rect 7301 13141 7313 13144
rect 7347 13141 7359 13175
rect 7301 13135 7359 13141
rect 9214 13132 9220 13184
rect 9272 13172 9278 13184
rect 9585 13175 9643 13181
rect 9585 13172 9597 13175
rect 9272 13144 9597 13172
rect 9272 13132 9278 13144
rect 9585 13141 9597 13144
rect 9631 13141 9643 13175
rect 9585 13135 9643 13141
rect 13446 13132 13452 13184
rect 13504 13132 13510 13184
rect 1104 13082 28888 13104
rect 1104 13030 3658 13082
rect 3710 13030 3722 13082
rect 3774 13030 3786 13082
rect 3838 13030 3850 13082
rect 3902 13030 3914 13082
rect 3966 13030 3978 13082
rect 4030 13030 11658 13082
rect 11710 13030 11722 13082
rect 11774 13030 11786 13082
rect 11838 13030 11850 13082
rect 11902 13030 11914 13082
rect 11966 13030 11978 13082
rect 12030 13030 19658 13082
rect 19710 13030 19722 13082
rect 19774 13030 19786 13082
rect 19838 13030 19850 13082
rect 19902 13030 19914 13082
rect 19966 13030 19978 13082
rect 20030 13030 27658 13082
rect 27710 13030 27722 13082
rect 27774 13030 27786 13082
rect 27838 13030 27850 13082
rect 27902 13030 27914 13082
rect 27966 13030 27978 13082
rect 28030 13030 28888 13082
rect 1104 13008 28888 13030
rect 1210 12928 1216 12980
rect 1268 12968 1274 12980
rect 1673 12971 1731 12977
rect 1673 12968 1685 12971
rect 1268 12940 1685 12968
rect 1268 12928 1274 12940
rect 1673 12937 1685 12940
rect 1719 12937 1731 12971
rect 1673 12931 1731 12937
rect 2774 12928 2780 12980
rect 2832 12928 2838 12980
rect 3418 12928 3424 12980
rect 3476 12928 3482 12980
rect 3602 12928 3608 12980
rect 3660 12968 3666 12980
rect 6546 12968 6552 12980
rect 3660 12940 6552 12968
rect 3660 12928 3666 12940
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 6917 12971 6975 12977
rect 6917 12937 6929 12971
rect 6963 12968 6975 12971
rect 7190 12968 7196 12980
rect 6963 12940 7196 12968
rect 6963 12937 6975 12940
rect 6917 12931 6975 12937
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 9214 12928 9220 12980
rect 9272 12928 9278 12980
rect 11422 12928 11428 12980
rect 11480 12968 11486 12980
rect 12710 12968 12716 12980
rect 11480 12940 12716 12968
rect 11480 12928 11486 12940
rect 2409 12903 2467 12909
rect 2409 12869 2421 12903
rect 2455 12900 2467 12903
rect 2792 12900 2820 12928
rect 4062 12900 4068 12912
rect 2455 12872 4068 12900
rect 2455 12869 2467 12872
rect 2409 12863 2467 12869
rect 4062 12860 4068 12872
rect 4120 12860 4126 12912
rect 8386 12860 8392 12912
rect 8444 12900 8450 12912
rect 11793 12903 11851 12909
rect 8444 12872 8984 12900
rect 8444 12860 8450 12872
rect 1302 12792 1308 12844
rect 1360 12832 1366 12844
rect 1397 12835 1455 12841
rect 1397 12832 1409 12835
rect 1360 12804 1409 12832
rect 1360 12792 1366 12804
rect 1397 12801 1409 12804
rect 1443 12832 1455 12835
rect 1857 12835 1915 12841
rect 1857 12832 1869 12835
rect 1443 12804 1869 12832
rect 1443 12801 1455 12804
rect 1397 12795 1455 12801
rect 1857 12801 1869 12804
rect 1903 12801 1915 12835
rect 1857 12795 1915 12801
rect 2590 12792 2596 12844
rect 2648 12841 2654 12844
rect 2648 12835 2681 12841
rect 2669 12801 2681 12835
rect 2648 12795 2681 12801
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12832 2835 12835
rect 2958 12832 2964 12844
rect 2823 12804 2964 12832
rect 2823 12801 2835 12804
rect 2777 12795 2835 12801
rect 2648 12792 2654 12795
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 3053 12835 3111 12841
rect 3053 12801 3065 12835
rect 3099 12832 3111 12835
rect 3326 12832 3332 12844
rect 3099 12804 3332 12832
rect 3099 12801 3111 12804
rect 3053 12795 3111 12801
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 6270 12792 6276 12844
rect 6328 12832 6334 12844
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6328 12804 6561 12832
rect 6328 12792 6334 12804
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 8846 12792 8852 12844
rect 8904 12792 8910 12844
rect 8956 12841 8984 12872
rect 11793 12869 11805 12903
rect 11839 12900 11851 12903
rect 12066 12900 12072 12912
rect 11839 12872 12072 12900
rect 11839 12869 11851 12872
rect 11793 12863 11851 12869
rect 12066 12860 12072 12872
rect 12124 12860 12130 12912
rect 12176 12900 12204 12940
rect 12710 12928 12716 12940
rect 12768 12928 12774 12980
rect 13262 12928 13268 12980
rect 13320 12928 13326 12980
rect 14826 12928 14832 12980
rect 14884 12968 14890 12980
rect 15838 12968 15844 12980
rect 14884 12940 15844 12968
rect 14884 12928 14890 12940
rect 15838 12928 15844 12940
rect 15896 12928 15902 12980
rect 18782 12928 18788 12980
rect 18840 12968 18846 12980
rect 19153 12971 19211 12977
rect 19153 12968 19165 12971
rect 18840 12940 19165 12968
rect 18840 12928 18846 12940
rect 19153 12937 19165 12940
rect 19199 12968 19211 12971
rect 19797 12971 19855 12977
rect 19797 12968 19809 12971
rect 19199 12940 19809 12968
rect 19199 12937 19211 12940
rect 19153 12931 19211 12937
rect 19797 12937 19809 12940
rect 19843 12937 19855 12971
rect 19797 12931 19855 12937
rect 12176 12872 12282 12900
rect 15286 12860 15292 12912
rect 15344 12900 15350 12912
rect 15749 12903 15807 12909
rect 15749 12900 15761 12903
rect 15344 12872 15761 12900
rect 15344 12860 15350 12872
rect 15749 12869 15761 12872
rect 15795 12900 15807 12903
rect 16942 12900 16948 12912
rect 15795 12872 16948 12900
rect 15795 12869 15807 12872
rect 15749 12863 15807 12869
rect 16942 12860 16948 12872
rect 17000 12860 17006 12912
rect 18690 12860 18696 12912
rect 18748 12900 18754 12912
rect 19061 12903 19119 12909
rect 19061 12900 19073 12903
rect 18748 12872 19073 12900
rect 18748 12860 18754 12872
rect 19061 12869 19073 12872
rect 19107 12900 19119 12903
rect 19889 12903 19947 12909
rect 19889 12900 19901 12903
rect 19107 12872 19901 12900
rect 19107 12869 19119 12872
rect 19061 12863 19119 12869
rect 19889 12869 19901 12872
rect 19935 12869 19947 12903
rect 19889 12863 19947 12869
rect 8942 12835 9000 12841
rect 8942 12801 8954 12835
rect 8988 12801 9000 12835
rect 8942 12795 9000 12801
rect 11330 12792 11336 12844
rect 11388 12832 11394 12844
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 11388 12804 11529 12832
rect 11388 12792 11394 12804
rect 11517 12801 11529 12804
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 13357 12835 13415 12841
rect 13357 12801 13369 12835
rect 13403 12832 13415 12835
rect 13446 12832 13452 12844
rect 13403 12804 13452 12832
rect 13403 12801 13415 12804
rect 13357 12795 13415 12801
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 13630 12792 13636 12844
rect 13688 12792 13694 12844
rect 2406 12724 2412 12776
rect 2464 12764 2470 12776
rect 3145 12767 3203 12773
rect 3145 12764 3157 12767
rect 2464 12736 3157 12764
rect 2464 12724 2470 12736
rect 3145 12733 3157 12736
rect 3191 12733 3203 12767
rect 3145 12727 3203 12733
rect 3234 12724 3240 12776
rect 3292 12764 3298 12776
rect 3418 12764 3424 12776
rect 3292 12736 3424 12764
rect 3292 12724 3298 12736
rect 3418 12724 3424 12736
rect 3476 12724 3482 12776
rect 6454 12724 6460 12776
rect 6512 12724 6518 12776
rect 18782 12724 18788 12776
rect 18840 12764 18846 12776
rect 19245 12767 19303 12773
rect 19245 12764 19257 12767
rect 18840 12736 19257 12764
rect 18840 12724 18846 12736
rect 19245 12733 19257 12736
rect 19291 12764 19303 12767
rect 19518 12764 19524 12776
rect 19291 12736 19524 12764
rect 19291 12733 19303 12736
rect 19245 12727 19303 12733
rect 19518 12724 19524 12736
rect 19576 12724 19582 12776
rect 19705 12767 19763 12773
rect 19705 12733 19717 12767
rect 19751 12764 19763 12767
rect 20530 12764 20536 12776
rect 19751 12736 20536 12764
rect 19751 12733 19763 12736
rect 19705 12727 19763 12733
rect 20530 12724 20536 12736
rect 20588 12764 20594 12776
rect 21174 12764 21180 12776
rect 20588 12736 21180 12764
rect 20588 12724 20594 12736
rect 21174 12724 21180 12736
rect 21232 12724 21238 12776
rect 1581 12699 1639 12705
rect 1581 12665 1593 12699
rect 1627 12696 1639 12699
rect 2866 12696 2872 12708
rect 1627 12668 2872 12696
rect 1627 12665 1639 12668
rect 1581 12659 1639 12665
rect 2866 12656 2872 12668
rect 2924 12656 2930 12708
rect 2958 12656 2964 12708
rect 3016 12696 3022 12708
rect 3602 12696 3608 12708
rect 3016 12668 3608 12696
rect 3016 12656 3022 12668
rect 3602 12656 3608 12668
rect 3660 12656 3666 12708
rect 2038 12588 2044 12640
rect 2096 12628 2102 12640
rect 3237 12631 3295 12637
rect 3237 12628 3249 12631
rect 2096 12600 3249 12628
rect 2096 12588 2102 12600
rect 3237 12597 3249 12600
rect 3283 12628 3295 12631
rect 6270 12628 6276 12640
rect 3283 12600 6276 12628
rect 3283 12597 3295 12600
rect 3237 12591 3295 12597
rect 6270 12588 6276 12600
rect 6328 12588 6334 12640
rect 11333 12631 11391 12637
rect 11333 12597 11345 12631
rect 11379 12628 11391 12631
rect 11422 12628 11428 12640
rect 11379 12600 11428 12628
rect 11379 12597 11391 12600
rect 11333 12591 11391 12597
rect 11422 12588 11428 12600
rect 11480 12588 11486 12640
rect 16758 12588 16764 12640
rect 16816 12588 16822 12640
rect 18690 12588 18696 12640
rect 18748 12588 18754 12640
rect 20257 12631 20315 12637
rect 20257 12597 20269 12631
rect 20303 12628 20315 12631
rect 22002 12628 22008 12640
rect 20303 12600 22008 12628
rect 20303 12597 20315 12600
rect 20257 12591 20315 12597
rect 22002 12588 22008 12600
rect 22060 12588 22066 12640
rect 1104 12538 28888 12560
rect 1104 12486 2918 12538
rect 2970 12486 2982 12538
rect 3034 12486 3046 12538
rect 3098 12486 3110 12538
rect 3162 12486 3174 12538
rect 3226 12486 3238 12538
rect 3290 12486 10918 12538
rect 10970 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 11238 12538
rect 11290 12486 18918 12538
rect 18970 12486 18982 12538
rect 19034 12486 19046 12538
rect 19098 12486 19110 12538
rect 19162 12486 19174 12538
rect 19226 12486 19238 12538
rect 19290 12486 26918 12538
rect 26970 12486 26982 12538
rect 27034 12486 27046 12538
rect 27098 12486 27110 12538
rect 27162 12486 27174 12538
rect 27226 12486 27238 12538
rect 27290 12486 28888 12538
rect 1104 12464 28888 12486
rect 3053 12427 3111 12433
rect 3053 12393 3065 12427
rect 3099 12424 3111 12427
rect 3326 12424 3332 12436
rect 3099 12396 3332 12424
rect 3099 12393 3111 12396
rect 3053 12387 3111 12393
rect 3326 12384 3332 12396
rect 3384 12384 3390 12436
rect 12526 12384 12532 12436
rect 12584 12424 12590 12436
rect 12805 12427 12863 12433
rect 12805 12424 12817 12427
rect 12584 12396 12817 12424
rect 12584 12384 12590 12396
rect 12805 12393 12817 12396
rect 12851 12393 12863 12427
rect 12805 12387 12863 12393
rect 13630 12384 13636 12436
rect 13688 12424 13694 12436
rect 20806 12424 20812 12436
rect 13688 12396 20812 12424
rect 13688 12384 13694 12396
rect 20806 12384 20812 12396
rect 20864 12384 20870 12436
rect 2961 12359 3019 12365
rect 2961 12325 2973 12359
rect 3007 12356 3019 12359
rect 3602 12356 3608 12368
rect 3007 12328 3608 12356
rect 3007 12325 3019 12328
rect 2961 12319 3019 12325
rect 3602 12316 3608 12328
rect 3660 12316 3666 12368
rect 11885 12359 11943 12365
rect 11885 12325 11897 12359
rect 11931 12356 11943 12359
rect 12713 12359 12771 12365
rect 11931 12328 12664 12356
rect 11931 12325 11943 12328
rect 11885 12319 11943 12325
rect 1946 12248 1952 12300
rect 2004 12248 2010 12300
rect 12161 12291 12219 12297
rect 12161 12257 12173 12291
rect 12207 12288 12219 12291
rect 12526 12288 12532 12300
rect 12207 12260 12532 12288
rect 12207 12257 12219 12260
rect 12161 12251 12219 12257
rect 12526 12248 12532 12260
rect 12584 12248 12590 12300
rect 12636 12288 12664 12328
rect 12713 12325 12725 12359
rect 12759 12356 12771 12359
rect 13814 12356 13820 12368
rect 12759 12328 13820 12356
rect 12759 12325 12771 12328
rect 12713 12319 12771 12325
rect 13814 12316 13820 12328
rect 13872 12316 13878 12368
rect 21910 12316 21916 12368
rect 21968 12356 21974 12368
rect 21968 12328 23888 12356
rect 21968 12316 21974 12328
rect 13354 12288 13360 12300
rect 12636 12260 13360 12288
rect 13354 12248 13360 12260
rect 13412 12288 13418 12300
rect 13449 12291 13507 12297
rect 13449 12288 13461 12291
rect 13412 12260 13461 12288
rect 13412 12248 13418 12260
rect 13449 12257 13461 12260
rect 13495 12288 13507 12291
rect 13722 12288 13728 12300
rect 13495 12260 13728 12288
rect 13495 12257 13507 12260
rect 13449 12251 13507 12257
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 14734 12248 14740 12300
rect 14792 12288 14798 12300
rect 14921 12291 14979 12297
rect 14921 12288 14933 12291
rect 14792 12260 14933 12288
rect 14792 12248 14798 12260
rect 14921 12257 14933 12260
rect 14967 12257 14979 12291
rect 14921 12251 14979 12257
rect 22002 12248 22008 12300
rect 22060 12288 22066 12300
rect 23860 12297 23888 12328
rect 24486 12316 24492 12368
rect 24544 12316 24550 12368
rect 24670 12316 24676 12368
rect 24728 12316 24734 12368
rect 23661 12291 23719 12297
rect 23661 12288 23673 12291
rect 22060 12260 23673 12288
rect 22060 12248 22066 12260
rect 23661 12257 23673 12260
rect 23707 12257 23719 12291
rect 23661 12251 23719 12257
rect 23845 12291 23903 12297
rect 23845 12257 23857 12291
rect 23891 12288 23903 12291
rect 24504 12288 24532 12316
rect 23891 12260 24532 12288
rect 23891 12257 23903 12260
rect 23845 12251 23903 12257
rect 1302 12180 1308 12232
rect 1360 12220 1366 12232
rect 2225 12223 2283 12229
rect 2225 12220 2237 12223
rect 1360 12192 2237 12220
rect 1360 12180 1366 12192
rect 2225 12189 2237 12192
rect 2271 12220 2283 12223
rect 2317 12223 2375 12229
rect 2317 12220 2329 12223
rect 2271 12192 2329 12220
rect 2271 12189 2283 12192
rect 2225 12183 2283 12189
rect 2317 12189 2329 12192
rect 2363 12189 2375 12223
rect 2317 12183 2375 12189
rect 4249 12223 4307 12229
rect 4249 12189 4261 12223
rect 4295 12220 4307 12223
rect 5718 12220 5724 12232
rect 4295 12192 5724 12220
rect 4295 12189 4307 12192
rect 4249 12183 4307 12189
rect 5718 12180 5724 12192
rect 5776 12180 5782 12232
rect 10686 12180 10692 12232
rect 10744 12220 10750 12232
rect 11701 12223 11759 12229
rect 11701 12220 11713 12223
rect 10744 12192 11713 12220
rect 10744 12180 10750 12192
rect 11701 12189 11713 12192
rect 11747 12189 11759 12223
rect 13265 12223 13323 12229
rect 13265 12220 13277 12223
rect 11701 12183 11759 12189
rect 12268 12192 13277 12220
rect 2590 12112 2596 12164
rect 2648 12112 2654 12164
rect 4154 12044 4160 12096
rect 4212 12044 4218 12096
rect 11146 12044 11152 12096
rect 11204 12084 11210 12096
rect 12268 12093 12296 12192
rect 13265 12189 13277 12192
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 16758 12180 16764 12232
rect 16816 12180 16822 12232
rect 17037 12223 17095 12229
rect 17037 12220 17049 12223
rect 16868 12192 17049 12220
rect 12526 12112 12532 12164
rect 12584 12152 12590 12164
rect 13630 12152 13636 12164
rect 12584 12124 13636 12152
rect 12584 12112 12590 12124
rect 13630 12112 13636 12124
rect 13688 12112 13694 12164
rect 15197 12155 15255 12161
rect 15197 12121 15209 12155
rect 15243 12152 15255 12155
rect 15286 12152 15292 12164
rect 15243 12124 15292 12152
rect 15243 12121 15255 12124
rect 15197 12115 15255 12121
rect 15286 12112 15292 12124
rect 15344 12112 15350 12164
rect 16206 12112 16212 12164
rect 16264 12112 16270 12164
rect 16482 12112 16488 12164
rect 16540 12152 16546 12164
rect 16868 12152 16896 12192
rect 17037 12189 17049 12192
rect 17083 12220 17095 12223
rect 24489 12223 24547 12229
rect 24489 12220 24501 12223
rect 17083 12192 24501 12220
rect 17083 12189 17095 12192
rect 17037 12183 17095 12189
rect 24489 12189 24501 12192
rect 24535 12189 24547 12223
rect 24489 12183 24547 12189
rect 16540 12124 16896 12152
rect 16540 12112 16546 12124
rect 16942 12112 16948 12164
rect 17000 12152 17006 12164
rect 21729 12155 21787 12161
rect 21729 12152 21741 12155
rect 17000 12124 21741 12152
rect 17000 12112 17006 12124
rect 21729 12121 21741 12124
rect 21775 12152 21787 12155
rect 21818 12152 21824 12164
rect 21775 12124 21824 12152
rect 21775 12121 21787 12124
rect 21729 12115 21787 12121
rect 21818 12112 21824 12124
rect 21876 12112 21882 12164
rect 12253 12087 12311 12093
rect 12253 12084 12265 12087
rect 11204 12056 12265 12084
rect 11204 12044 11210 12056
rect 12253 12053 12265 12056
rect 12299 12053 12311 12087
rect 12253 12047 12311 12053
rect 12345 12087 12403 12093
rect 12345 12053 12357 12087
rect 12391 12084 12403 12087
rect 13173 12087 13231 12093
rect 13173 12084 13185 12087
rect 12391 12056 13185 12084
rect 12391 12053 12403 12056
rect 12345 12047 12403 12053
rect 13173 12053 13185 12056
rect 13219 12084 13231 12087
rect 13262 12084 13268 12096
rect 13219 12056 13268 12084
rect 13219 12053 13231 12056
rect 13173 12047 13231 12053
rect 13262 12044 13268 12056
rect 13320 12044 13326 12096
rect 16666 12044 16672 12096
rect 16724 12044 16730 12096
rect 23201 12087 23259 12093
rect 23201 12053 23213 12087
rect 23247 12084 23259 12087
rect 23290 12084 23296 12096
rect 23247 12056 23296 12084
rect 23247 12053 23259 12056
rect 23201 12047 23259 12053
rect 23290 12044 23296 12056
rect 23348 12044 23354 12096
rect 23566 12044 23572 12096
rect 23624 12044 23630 12096
rect 1104 11994 28888 12016
rect 1104 11942 3658 11994
rect 3710 11942 3722 11994
rect 3774 11942 3786 11994
rect 3838 11942 3850 11994
rect 3902 11942 3914 11994
rect 3966 11942 3978 11994
rect 4030 11942 11658 11994
rect 11710 11942 11722 11994
rect 11774 11942 11786 11994
rect 11838 11942 11850 11994
rect 11902 11942 11914 11994
rect 11966 11942 11978 11994
rect 12030 11942 19658 11994
rect 19710 11942 19722 11994
rect 19774 11942 19786 11994
rect 19838 11942 19850 11994
rect 19902 11942 19914 11994
rect 19966 11942 19978 11994
rect 20030 11942 27658 11994
rect 27710 11942 27722 11994
rect 27774 11942 27786 11994
rect 27838 11942 27850 11994
rect 27902 11942 27914 11994
rect 27966 11942 27978 11994
rect 28030 11942 28888 11994
rect 1104 11920 28888 11942
rect 2406 11840 2412 11892
rect 2464 11840 2470 11892
rect 8846 11840 8852 11892
rect 8904 11880 8910 11892
rect 9309 11883 9367 11889
rect 9309 11880 9321 11883
rect 8904 11852 9321 11880
rect 8904 11840 8910 11852
rect 9309 11849 9321 11852
rect 9355 11880 9367 11883
rect 9355 11852 11008 11880
rect 9355 11849 9367 11852
rect 9309 11843 9367 11849
rect 10980 11812 11008 11852
rect 15286 11840 15292 11892
rect 15344 11840 15350 11892
rect 15562 11840 15568 11892
rect 15620 11880 15626 11892
rect 16206 11880 16212 11892
rect 15620 11852 16212 11880
rect 15620 11840 15626 11852
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 18690 11840 18696 11892
rect 18748 11880 18754 11892
rect 18785 11883 18843 11889
rect 18785 11880 18797 11883
rect 18748 11852 18797 11880
rect 18748 11840 18754 11852
rect 18785 11849 18797 11852
rect 18831 11849 18843 11883
rect 18785 11843 18843 11849
rect 22278 11840 22284 11892
rect 22336 11840 22342 11892
rect 23566 11840 23572 11892
rect 23624 11880 23630 11892
rect 24762 11880 24768 11892
rect 23624 11852 24768 11880
rect 23624 11840 23630 11852
rect 24762 11840 24768 11852
rect 24820 11840 24826 11892
rect 11422 11812 11428 11824
rect 10902 11784 11428 11812
rect 11422 11772 11428 11784
rect 11480 11772 11486 11824
rect 15657 11815 15715 11821
rect 15657 11781 15669 11815
rect 15703 11812 15715 11815
rect 16666 11812 16672 11824
rect 15703 11784 16672 11812
rect 15703 11781 15715 11784
rect 15657 11775 15715 11781
rect 16666 11772 16672 11784
rect 16724 11772 16730 11824
rect 23290 11772 23296 11824
rect 23348 11772 23354 11824
rect 24578 11812 24584 11824
rect 24518 11784 24584 11812
rect 24578 11772 24584 11784
rect 24636 11772 24642 11824
rect 1946 11704 1952 11756
rect 2004 11704 2010 11756
rect 2314 11704 2320 11756
rect 2372 11704 2378 11756
rect 2774 11704 2780 11756
rect 2832 11744 2838 11756
rect 2869 11747 2927 11753
rect 2869 11744 2881 11747
rect 2832 11716 2881 11744
rect 2832 11704 2838 11716
rect 2869 11713 2881 11716
rect 2915 11713 2927 11747
rect 13265 11747 13323 11753
rect 13265 11744 13277 11747
rect 2869 11707 2927 11713
rect 13096 11716 13277 11744
rect 1302 11636 1308 11688
rect 1360 11676 1366 11688
rect 2225 11679 2283 11685
rect 2225 11676 2237 11679
rect 1360 11648 2237 11676
rect 1360 11636 1366 11648
rect 2225 11645 2237 11648
rect 2271 11676 2283 11679
rect 2593 11679 2651 11685
rect 2593 11676 2605 11679
rect 2271 11648 2605 11676
rect 2271 11645 2283 11648
rect 2225 11639 2283 11645
rect 2593 11645 2605 11648
rect 2639 11645 2651 11679
rect 2593 11639 2651 11645
rect 2682 11636 2688 11688
rect 2740 11676 2746 11688
rect 3145 11679 3203 11685
rect 3145 11676 3157 11679
rect 2740 11648 3157 11676
rect 2740 11636 2746 11648
rect 3145 11645 3157 11648
rect 3191 11645 3203 11679
rect 3145 11639 3203 11645
rect 9398 11636 9404 11688
rect 9456 11636 9462 11688
rect 9674 11636 9680 11688
rect 9732 11636 9738 11688
rect 1026 11568 1032 11620
rect 1084 11608 1090 11620
rect 13096 11617 13124 11716
rect 13265 11713 13277 11716
rect 13311 11713 13323 11747
rect 13265 11707 13323 11713
rect 15010 11704 15016 11756
rect 15068 11744 15074 11756
rect 16114 11744 16120 11756
rect 15068 11716 16120 11744
rect 15068 11704 15074 11716
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11744 16359 11747
rect 16482 11744 16488 11756
rect 16347 11716 16488 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 16482 11704 16488 11716
rect 16540 11704 16546 11756
rect 16592 11716 16804 11744
rect 15746 11636 15752 11688
rect 15804 11636 15810 11688
rect 15838 11636 15844 11688
rect 15896 11676 15902 11688
rect 15933 11679 15991 11685
rect 15933 11676 15945 11679
rect 15896 11648 15945 11676
rect 15896 11636 15902 11648
rect 15933 11645 15945 11648
rect 15979 11676 15991 11679
rect 16592 11676 16620 11716
rect 15979 11648 16620 11676
rect 15979 11645 15991 11648
rect 15933 11639 15991 11645
rect 16666 11636 16672 11688
rect 16724 11636 16730 11688
rect 16776 11676 16804 11716
rect 16942 11704 16948 11756
rect 17000 11704 17006 11756
rect 18693 11747 18751 11753
rect 18693 11713 18705 11747
rect 18739 11744 18751 11747
rect 19426 11744 19432 11756
rect 18739 11716 19432 11744
rect 18739 11713 18751 11716
rect 18693 11707 18751 11713
rect 19426 11704 19432 11716
rect 19484 11704 19490 11756
rect 20714 11704 20720 11756
rect 20772 11744 20778 11756
rect 22189 11747 22247 11753
rect 22189 11744 22201 11747
rect 20772 11716 22201 11744
rect 20772 11704 20778 11716
rect 22189 11713 22201 11716
rect 22235 11713 22247 11747
rect 22189 11707 22247 11713
rect 18877 11679 18935 11685
rect 18877 11676 18889 11679
rect 16776 11648 18889 11676
rect 18877 11645 18889 11648
rect 18923 11645 18935 11679
rect 18877 11639 18935 11645
rect 21910 11636 21916 11688
rect 21968 11676 21974 11688
rect 22373 11679 22431 11685
rect 22373 11676 22385 11679
rect 21968 11648 22385 11676
rect 21968 11636 21974 11648
rect 22373 11645 22385 11648
rect 22419 11645 22431 11679
rect 22373 11639 22431 11645
rect 23017 11679 23075 11685
rect 23017 11645 23029 11679
rect 23063 11645 23075 11679
rect 23017 11639 23075 11645
rect 13081 11611 13139 11617
rect 13081 11608 13093 11611
rect 1084 11580 9352 11608
rect 1084 11568 1090 11580
rect 3237 11543 3295 11549
rect 3237 11509 3249 11543
rect 3283 11540 3295 11543
rect 3326 11540 3332 11552
rect 3283 11512 3332 11540
rect 3283 11509 3295 11512
rect 3237 11503 3295 11509
rect 3326 11500 3332 11512
rect 3384 11500 3390 11552
rect 3421 11543 3479 11549
rect 3421 11509 3433 11543
rect 3467 11540 3479 11543
rect 3602 11540 3608 11552
rect 3467 11512 3608 11540
rect 3467 11509 3479 11512
rect 3421 11503 3479 11509
rect 3602 11500 3608 11512
rect 3660 11540 3666 11552
rect 4246 11540 4252 11552
rect 3660 11512 4252 11540
rect 3660 11500 3666 11512
rect 4246 11500 4252 11512
rect 4304 11500 4310 11552
rect 9324 11540 9352 11580
rect 10704 11580 13093 11608
rect 10704 11540 10732 11580
rect 13081 11577 13093 11580
rect 13127 11577 13139 11611
rect 19334 11608 19340 11620
rect 13081 11571 13139 11577
rect 15120 11580 19340 11608
rect 9324 11512 10732 11540
rect 10778 11500 10784 11552
rect 10836 11540 10842 11552
rect 11146 11540 11152 11552
rect 10836 11512 11152 11540
rect 10836 11500 10842 11512
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 11422 11500 11428 11552
rect 11480 11540 11486 11552
rect 15120 11549 15148 11580
rect 19334 11568 19340 11580
rect 19392 11568 19398 11620
rect 22002 11568 22008 11620
rect 22060 11608 22066 11620
rect 23032 11608 23060 11639
rect 22060 11580 23060 11608
rect 22060 11568 22066 11580
rect 14553 11543 14611 11549
rect 14553 11540 14565 11543
rect 11480 11512 14565 11540
rect 11480 11500 11486 11512
rect 14553 11509 14565 11512
rect 14599 11540 14611 11543
rect 15105 11543 15163 11549
rect 15105 11540 15117 11543
rect 14599 11512 15117 11540
rect 14599 11509 14611 11512
rect 14553 11503 14611 11509
rect 15105 11509 15117 11512
rect 15151 11509 15163 11543
rect 15105 11503 15163 11509
rect 17586 11500 17592 11552
rect 17644 11540 17650 11552
rect 18325 11543 18383 11549
rect 18325 11540 18337 11543
rect 17644 11512 18337 11540
rect 17644 11500 17650 11512
rect 18325 11509 18337 11512
rect 18371 11509 18383 11543
rect 18325 11503 18383 11509
rect 21821 11543 21879 11549
rect 21821 11509 21833 11543
rect 21867 11540 21879 11543
rect 22094 11540 22100 11552
rect 21867 11512 22100 11540
rect 21867 11509 21879 11512
rect 21821 11503 21879 11509
rect 22094 11500 22100 11512
rect 22152 11500 22158 11552
rect 1104 11450 28888 11472
rect 1104 11398 2918 11450
rect 2970 11398 2982 11450
rect 3034 11398 3046 11450
rect 3098 11398 3110 11450
rect 3162 11398 3174 11450
rect 3226 11398 3238 11450
rect 3290 11398 10918 11450
rect 10970 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 11238 11450
rect 11290 11398 18918 11450
rect 18970 11398 18982 11450
rect 19034 11398 19046 11450
rect 19098 11398 19110 11450
rect 19162 11398 19174 11450
rect 19226 11398 19238 11450
rect 19290 11398 26918 11450
rect 26970 11398 26982 11450
rect 27034 11398 27046 11450
rect 27098 11398 27110 11450
rect 27162 11398 27174 11450
rect 27226 11398 27238 11450
rect 27290 11398 28888 11450
rect 1104 11376 28888 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 2130 11336 2136 11348
rect 1627 11308 2136 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 2317 11339 2375 11345
rect 2317 11305 2329 11339
rect 2363 11336 2375 11339
rect 2682 11336 2688 11348
rect 2363 11308 2688 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 3145 11339 3203 11345
rect 3145 11305 3157 11339
rect 3191 11336 3203 11339
rect 3694 11336 3700 11348
rect 3191 11308 3700 11336
rect 3191 11305 3203 11308
rect 3145 11299 3203 11305
rect 3694 11296 3700 11308
rect 3752 11296 3758 11348
rect 3786 11296 3792 11348
rect 3844 11296 3850 11348
rect 3878 11296 3884 11348
rect 3936 11336 3942 11348
rect 3936 11308 4752 11336
rect 3936 11296 3942 11308
rect 4338 11268 4344 11280
rect 3620 11240 4344 11268
rect 2038 11160 2044 11212
rect 2096 11160 2102 11212
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 1949 11135 2007 11141
rect 1949 11132 1961 11135
rect 1636 11104 1961 11132
rect 1636 11092 1642 11104
rect 1949 11101 1961 11104
rect 1995 11132 2007 11135
rect 2314 11132 2320 11144
rect 1995 11104 2320 11132
rect 1995 11101 2007 11104
rect 1949 11095 2007 11101
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 3329 11135 3387 11141
rect 3329 11101 3341 11135
rect 3375 11132 3387 11135
rect 3510 11132 3516 11144
rect 3375 11104 3516 11132
rect 3375 11101 3387 11104
rect 3329 11095 3387 11101
rect 3510 11092 3516 11104
rect 3568 11092 3574 11144
rect 3620 11141 3648 11240
rect 4338 11228 4344 11240
rect 4396 11268 4402 11280
rect 4617 11271 4675 11277
rect 4617 11268 4629 11271
rect 4396 11240 4629 11268
rect 4396 11228 4402 11240
rect 4617 11237 4629 11240
rect 4663 11237 4675 11271
rect 4617 11231 4675 11237
rect 4154 11200 4160 11212
rect 3988 11172 4160 11200
rect 3988 11141 4016 11172
rect 4154 11160 4160 11172
rect 4212 11200 4218 11212
rect 4724 11209 4752 11308
rect 14366 11296 14372 11348
rect 14424 11336 14430 11348
rect 14461 11339 14519 11345
rect 14461 11336 14473 11339
rect 14424 11308 14473 11336
rect 14424 11296 14430 11308
rect 14461 11305 14473 11308
rect 14507 11305 14519 11339
rect 14461 11299 14519 11305
rect 15746 11296 15752 11348
rect 15804 11336 15810 11348
rect 16025 11339 16083 11345
rect 16025 11336 16037 11339
rect 15804 11308 16037 11336
rect 15804 11296 15810 11308
rect 16025 11305 16037 11308
rect 16071 11305 16083 11339
rect 19061 11339 19119 11345
rect 16025 11299 16083 11305
rect 16132 11308 18828 11336
rect 13722 11228 13728 11280
rect 13780 11268 13786 11280
rect 16132 11268 16160 11308
rect 13780 11240 16160 11268
rect 13780 11228 13786 11240
rect 4525 11203 4583 11209
rect 4525 11200 4537 11203
rect 4212 11172 4537 11200
rect 4212 11160 4218 11172
rect 4525 11169 4537 11172
rect 4571 11169 4583 11203
rect 4525 11163 4583 11169
rect 4709 11203 4767 11209
rect 4709 11169 4721 11203
rect 4755 11169 4767 11203
rect 15010 11200 15016 11212
rect 4709 11163 4767 11169
rect 14108 11172 15016 11200
rect 3605 11135 3663 11141
rect 3605 11101 3617 11135
rect 3651 11101 3663 11135
rect 3605 11095 3663 11101
rect 3973 11135 4031 11141
rect 3973 11101 3985 11135
rect 4019 11101 4031 11135
rect 3973 11095 4031 11101
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 4080 11064 4108 11095
rect 4246 11092 4252 11144
rect 4304 11092 4310 11144
rect 4338 11092 4344 11144
rect 4396 11092 4402 11144
rect 4430 11092 4436 11144
rect 4488 11092 4494 11144
rect 4798 11092 4804 11144
rect 4856 11092 4862 11144
rect 8665 11135 8723 11141
rect 8665 11101 8677 11135
rect 8711 11132 8723 11135
rect 9398 11132 9404 11144
rect 8711 11104 9404 11132
rect 8711 11101 8723 11104
rect 8665 11095 8723 11101
rect 9398 11092 9404 11104
rect 9456 11092 9462 11144
rect 4448 11064 4476 11092
rect 4080 11036 4476 11064
rect 10689 11067 10747 11073
rect 10689 11033 10701 11067
rect 10735 11064 10747 11067
rect 10873 11067 10931 11073
rect 10873 11064 10885 11067
rect 10735 11036 10885 11064
rect 10735 11033 10747 11036
rect 10689 11027 10747 11033
rect 10873 11033 10885 11036
rect 10919 11064 10931 11067
rect 11422 11064 11428 11076
rect 10919 11036 11428 11064
rect 10919 11033 10931 11036
rect 10873 11027 10931 11033
rect 11422 11024 11428 11036
rect 11480 11024 11486 11076
rect 13998 11024 14004 11076
rect 14056 11064 14062 11076
rect 14108 11073 14136 11172
rect 15010 11160 15016 11172
rect 15068 11160 15074 11212
rect 15381 11203 15439 11209
rect 15381 11169 15393 11203
rect 15427 11169 15439 11203
rect 15381 11163 15439 11169
rect 15194 11132 15200 11144
rect 14292 11104 15200 11132
rect 14292 11076 14320 11104
rect 15194 11092 15200 11104
rect 15252 11132 15258 11144
rect 15396 11132 15424 11163
rect 17586 11160 17592 11212
rect 17644 11160 17650 11212
rect 15252 11104 15424 11132
rect 15252 11092 15258 11104
rect 15562 11092 15568 11144
rect 15620 11132 15626 11144
rect 16022 11132 16028 11144
rect 15620 11104 16028 11132
rect 15620 11092 15626 11104
rect 16022 11092 16028 11104
rect 16080 11132 16086 11144
rect 16482 11132 16488 11144
rect 16080 11104 16488 11132
rect 16080 11092 16086 11104
rect 16482 11092 16488 11104
rect 16540 11132 16546 11144
rect 16577 11135 16635 11141
rect 16577 11132 16589 11135
rect 16540 11104 16589 11132
rect 16540 11092 16546 11104
rect 16577 11101 16589 11104
rect 16623 11101 16635 11135
rect 16577 11095 16635 11101
rect 17310 11092 17316 11144
rect 17368 11092 17374 11144
rect 18800 11132 18828 11308
rect 19061 11305 19073 11339
rect 19107 11336 19119 11339
rect 19426 11336 19432 11348
rect 19107 11308 19432 11336
rect 19107 11305 19119 11308
rect 19061 11299 19119 11305
rect 19426 11296 19432 11308
rect 19484 11336 19490 11348
rect 19484 11308 20024 11336
rect 19484 11296 19490 11308
rect 19996 11268 20024 11308
rect 20622 11268 20628 11280
rect 19996 11240 20628 11268
rect 19996 11209 20024 11240
rect 20622 11228 20628 11240
rect 20680 11228 20686 11280
rect 23474 11228 23480 11280
rect 23532 11268 23538 11280
rect 24578 11268 24584 11280
rect 23532 11240 24584 11268
rect 23532 11228 23538 11240
rect 24578 11228 24584 11240
rect 24636 11268 24642 11280
rect 24636 11240 24992 11268
rect 24636 11228 24642 11240
rect 19981 11203 20039 11209
rect 19981 11169 19993 11203
rect 20027 11169 20039 11203
rect 19981 11163 20039 11169
rect 20073 11203 20131 11209
rect 20073 11169 20085 11203
rect 20119 11169 20131 11203
rect 20073 11163 20131 11169
rect 20088 11132 20116 11163
rect 22002 11160 22008 11212
rect 22060 11200 22066 11212
rect 22373 11203 22431 11209
rect 22373 11200 22385 11203
rect 22060 11172 22385 11200
rect 22060 11160 22066 11172
rect 22373 11169 22385 11172
rect 22419 11169 22431 11203
rect 22373 11163 22431 11169
rect 24762 11160 24768 11212
rect 24820 11200 24826 11212
rect 24964 11209 24992 11240
rect 24857 11203 24915 11209
rect 24857 11200 24869 11203
rect 24820 11172 24869 11200
rect 24820 11160 24826 11172
rect 24857 11169 24869 11172
rect 24903 11169 24915 11203
rect 24857 11163 24915 11169
rect 24949 11203 25007 11209
rect 24949 11169 24961 11203
rect 24995 11169 25007 11203
rect 24949 11163 25007 11169
rect 18800 11104 20116 11132
rect 14093 11067 14151 11073
rect 14093 11064 14105 11067
rect 14056 11036 14105 11064
rect 14056 11024 14062 11036
rect 14093 11033 14105 11036
rect 14139 11033 14151 11067
rect 14093 11027 14151 11033
rect 14274 11024 14280 11076
rect 14332 11024 14338 11076
rect 14829 11067 14887 11073
rect 14829 11033 14841 11067
rect 14875 11064 14887 11067
rect 15378 11064 15384 11076
rect 14875 11036 15384 11064
rect 14875 11033 14887 11036
rect 14829 11027 14887 11033
rect 15378 11024 15384 11036
rect 15436 11064 15442 11076
rect 15657 11067 15715 11073
rect 15657 11064 15669 11067
rect 15436 11036 15669 11064
rect 15436 11024 15442 11036
rect 15657 11033 15669 11036
rect 15703 11033 15715 11067
rect 15657 11027 15715 11033
rect 18046 11024 18052 11076
rect 18104 11024 18110 11076
rect 19889 11067 19947 11073
rect 19889 11033 19901 11067
rect 19935 11064 19947 11067
rect 19935 11036 20668 11064
rect 19935 11033 19947 11036
rect 19889 11027 19947 11033
rect 3510 10956 3516 11008
rect 3568 10996 3574 11008
rect 3878 10996 3884 11008
rect 3568 10968 3884 10996
rect 3568 10956 3574 10968
rect 3878 10956 3884 10968
rect 3936 10956 3942 11008
rect 9398 10956 9404 11008
rect 9456 10956 9462 11008
rect 14921 10999 14979 11005
rect 14921 10965 14933 10999
rect 14967 10996 14979 10999
rect 15286 10996 15292 11008
rect 14967 10968 15292 10996
rect 14967 10965 14979 10968
rect 14921 10959 14979 10965
rect 15286 10956 15292 10968
rect 15344 10996 15350 11008
rect 15565 10999 15623 11005
rect 15565 10996 15577 10999
rect 15344 10968 15577 10996
rect 15344 10956 15350 10968
rect 15565 10965 15577 10968
rect 15611 10965 15623 10999
rect 15565 10959 15623 10965
rect 19518 10956 19524 11008
rect 19576 10956 19582 11008
rect 20640 11005 20668 11036
rect 21634 11024 21640 11076
rect 21692 11024 21698 11076
rect 22094 11024 22100 11076
rect 22152 11024 22158 11076
rect 24670 11024 24676 11076
rect 24728 11064 24734 11076
rect 24765 11067 24823 11073
rect 24765 11064 24777 11067
rect 24728 11036 24777 11064
rect 24728 11024 24734 11036
rect 24765 11033 24777 11036
rect 24811 11033 24823 11067
rect 24765 11027 24823 11033
rect 20625 10999 20683 11005
rect 20625 10965 20637 10999
rect 20671 10996 20683 10999
rect 20714 10996 20720 11008
rect 20671 10968 20720 10996
rect 20671 10965 20683 10968
rect 20625 10959 20683 10965
rect 20714 10956 20720 10968
rect 20772 10956 20778 11008
rect 24394 10956 24400 11008
rect 24452 10956 24458 11008
rect 1104 10906 28888 10928
rect 1104 10854 3658 10906
rect 3710 10854 3722 10906
rect 3774 10854 3786 10906
rect 3838 10854 3850 10906
rect 3902 10854 3914 10906
rect 3966 10854 3978 10906
rect 4030 10854 11658 10906
rect 11710 10854 11722 10906
rect 11774 10854 11786 10906
rect 11838 10854 11850 10906
rect 11902 10854 11914 10906
rect 11966 10854 11978 10906
rect 12030 10854 19658 10906
rect 19710 10854 19722 10906
rect 19774 10854 19786 10906
rect 19838 10854 19850 10906
rect 19902 10854 19914 10906
rect 19966 10854 19978 10906
rect 20030 10854 27658 10906
rect 27710 10854 27722 10906
rect 27774 10854 27786 10906
rect 27838 10854 27850 10906
rect 27902 10854 27914 10906
rect 27966 10854 27978 10906
rect 28030 10854 28888 10906
rect 1104 10832 28888 10854
rect 1394 10752 1400 10804
rect 1452 10792 1458 10804
rect 1673 10795 1731 10801
rect 1673 10792 1685 10795
rect 1452 10764 1685 10792
rect 1452 10752 1458 10764
rect 1673 10761 1685 10764
rect 1719 10761 1731 10795
rect 1673 10755 1731 10761
rect 3510 10752 3516 10804
rect 3568 10792 3574 10804
rect 3605 10795 3663 10801
rect 3605 10792 3617 10795
rect 3568 10764 3617 10792
rect 3568 10752 3574 10764
rect 3605 10761 3617 10764
rect 3651 10761 3663 10795
rect 3605 10755 3663 10761
rect 4065 10795 4123 10801
rect 4065 10761 4077 10795
rect 4111 10792 4123 10795
rect 4798 10792 4804 10804
rect 4111 10764 4804 10792
rect 4111 10761 4123 10764
rect 4065 10755 4123 10761
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 9674 10752 9680 10804
rect 9732 10752 9738 10804
rect 10045 10795 10103 10801
rect 10045 10761 10057 10795
rect 10091 10792 10103 10795
rect 10778 10792 10784 10804
rect 10091 10764 10784 10792
rect 10091 10761 10103 10764
rect 10045 10755 10103 10761
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 11532 10764 13860 10792
rect 6914 10724 6920 10736
rect 3252 10696 6920 10724
rect 1302 10616 1308 10668
rect 1360 10656 1366 10668
rect 3252 10665 3280 10696
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 1360 10628 1409 10656
rect 1360 10616 1366 10628
rect 1397 10625 1409 10628
rect 1443 10656 1455 10659
rect 1857 10659 1915 10665
rect 1857 10656 1869 10659
rect 1443 10628 1869 10656
rect 1443 10625 1455 10628
rect 1397 10619 1455 10625
rect 1857 10625 1869 10628
rect 1903 10625 1915 10659
rect 1857 10619 1915 10625
rect 3237 10659 3295 10665
rect 3237 10625 3249 10659
rect 3283 10625 3295 10659
rect 3237 10619 3295 10625
rect 3326 10616 3332 10668
rect 3384 10656 3390 10668
rect 3866 10665 3894 10696
rect 6914 10684 6920 10696
rect 6972 10684 6978 10736
rect 7282 10684 7288 10736
rect 7340 10684 7346 10736
rect 9582 10724 9588 10736
rect 8956 10696 9588 10724
rect 3697 10659 3755 10665
rect 3697 10656 3709 10659
rect 3384 10628 3709 10656
rect 3384 10616 3390 10628
rect 3697 10625 3709 10628
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 3851 10659 3909 10665
rect 3851 10625 3863 10659
rect 3897 10656 3909 10659
rect 8956 10656 8984 10696
rect 9582 10684 9588 10696
rect 9640 10724 9646 10736
rect 10686 10724 10692 10736
rect 9640 10696 10692 10724
rect 9640 10684 9646 10696
rect 10686 10684 10692 10696
rect 10744 10684 10750 10736
rect 3897 10628 3931 10656
rect 8864 10628 8984 10656
rect 9033 10659 9091 10665
rect 3897 10625 3909 10628
rect 3851 10619 3909 10625
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 3344 10588 3372 10616
rect 2832 10560 3372 10588
rect 2832 10548 2838 10560
rect 6362 10548 6368 10600
rect 6420 10548 6426 10600
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10588 6699 10591
rect 7098 10588 7104 10600
rect 6687 10560 7104 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 7098 10548 7104 10560
rect 7156 10548 7162 10600
rect 8864 10597 8892 10628
rect 9033 10625 9045 10659
rect 9079 10625 9091 10659
rect 9033 10619 9091 10625
rect 8849 10591 8907 10597
rect 8849 10557 8861 10591
rect 8895 10557 8907 10591
rect 8849 10551 8907 10557
rect 8938 10548 8944 10600
rect 8996 10548 9002 10600
rect 1581 10523 1639 10529
rect 1581 10489 1593 10523
rect 1627 10520 1639 10523
rect 2222 10520 2228 10532
rect 1627 10492 2228 10520
rect 1627 10489 1639 10492
rect 1581 10483 1639 10489
rect 2222 10480 2228 10492
rect 2280 10480 2286 10532
rect 8110 10412 8116 10464
rect 8168 10452 8174 10464
rect 9048 10452 9076 10619
rect 11330 10616 11336 10668
rect 11388 10656 11394 10668
rect 11532 10665 11560 10764
rect 12434 10684 12440 10736
rect 12492 10684 12498 10736
rect 13832 10665 13860 10764
rect 20622 10752 20628 10804
rect 20680 10792 20686 10804
rect 20809 10795 20867 10801
rect 20809 10792 20821 10795
rect 20680 10764 20821 10792
rect 20680 10752 20686 10764
rect 20809 10761 20821 10764
rect 20855 10761 20867 10795
rect 20809 10755 20867 10761
rect 21269 10795 21327 10801
rect 21269 10761 21281 10795
rect 21315 10792 21327 10795
rect 24673 10795 24731 10801
rect 24673 10792 24685 10795
rect 21315 10764 24685 10792
rect 21315 10761 21327 10764
rect 21269 10755 21327 10761
rect 24673 10761 24685 10764
rect 24719 10761 24731 10795
rect 24673 10755 24731 10761
rect 18046 10724 18052 10736
rect 15318 10696 18052 10724
rect 18046 10684 18052 10696
rect 18104 10684 18110 10736
rect 20714 10684 20720 10736
rect 20772 10724 20778 10736
rect 20901 10727 20959 10733
rect 20901 10724 20913 10727
rect 20772 10696 20913 10724
rect 20772 10684 20778 10696
rect 20901 10693 20913 10696
rect 20947 10693 20959 10727
rect 20901 10687 20959 10693
rect 23845 10727 23903 10733
rect 23845 10693 23857 10727
rect 23891 10724 23903 10727
rect 24762 10724 24768 10736
rect 23891 10696 24768 10724
rect 23891 10693 23903 10696
rect 23845 10687 23903 10693
rect 24762 10684 24768 10696
rect 24820 10684 24826 10736
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 11388 10628 11529 10656
rect 11388 10616 11394 10628
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 11517 10619 11575 10625
rect 13817 10659 13875 10665
rect 13817 10625 13829 10659
rect 13863 10625 13875 10659
rect 13817 10619 13875 10625
rect 17954 10616 17960 10668
rect 18012 10656 18018 10668
rect 19245 10659 19303 10665
rect 19245 10656 19257 10659
rect 18012 10628 19257 10656
rect 18012 10616 18018 10628
rect 19245 10625 19257 10628
rect 19291 10625 19303 10659
rect 19245 10619 19303 10625
rect 23753 10659 23811 10665
rect 23753 10625 23765 10659
rect 23799 10656 23811 10659
rect 24581 10659 24639 10665
rect 23799 10628 24532 10656
rect 23799 10625 23811 10628
rect 23753 10619 23811 10625
rect 10137 10591 10195 10597
rect 10137 10588 10149 10591
rect 9416 10560 10149 10588
rect 9416 10529 9444 10560
rect 10137 10557 10149 10560
rect 10183 10557 10195 10591
rect 10137 10551 10195 10557
rect 10321 10591 10379 10597
rect 10321 10557 10333 10591
rect 10367 10588 10379 10591
rect 10367 10560 10456 10588
rect 10367 10557 10379 10560
rect 10321 10551 10379 10557
rect 9401 10523 9459 10529
rect 9401 10489 9413 10523
rect 9447 10489 9459 10523
rect 9401 10483 9459 10489
rect 8168 10424 9076 10452
rect 9585 10455 9643 10461
rect 8168 10412 8174 10424
rect 9585 10421 9597 10455
rect 9631 10452 9643 10455
rect 10428 10452 10456 10560
rect 11790 10548 11796 10600
rect 11848 10548 11854 10600
rect 14090 10548 14096 10600
rect 14148 10548 14154 10600
rect 15286 10548 15292 10600
rect 15344 10588 15350 10600
rect 15565 10591 15623 10597
rect 15565 10588 15577 10591
rect 15344 10560 15577 10588
rect 15344 10548 15350 10560
rect 15565 10557 15577 10560
rect 15611 10557 15623 10591
rect 15565 10551 15623 10557
rect 20717 10591 20775 10597
rect 20717 10557 20729 10591
rect 20763 10588 20775 10591
rect 20806 10588 20812 10600
rect 20763 10560 20812 10588
rect 20763 10557 20775 10560
rect 20717 10551 20775 10557
rect 20806 10548 20812 10560
rect 20864 10548 20870 10600
rect 23658 10548 23664 10600
rect 23716 10588 23722 10600
rect 23937 10591 23995 10597
rect 23937 10588 23949 10591
rect 23716 10560 23949 10588
rect 23716 10548 23722 10560
rect 23937 10557 23949 10560
rect 23983 10588 23995 10591
rect 24210 10588 24216 10600
rect 23983 10560 24216 10588
rect 23983 10557 23995 10560
rect 23937 10551 23995 10557
rect 24210 10548 24216 10560
rect 24268 10548 24274 10600
rect 24504 10588 24532 10628
rect 24581 10625 24593 10659
rect 24627 10656 24639 10659
rect 25038 10656 25044 10668
rect 24627 10628 25044 10656
rect 24627 10625 24639 10628
rect 24581 10619 24639 10625
rect 25038 10616 25044 10628
rect 25096 10616 25102 10668
rect 24670 10588 24676 10600
rect 24504 10560 24676 10588
rect 24670 10548 24676 10560
rect 24728 10548 24734 10600
rect 24765 10591 24823 10597
rect 24765 10557 24777 10591
rect 24811 10557 24823 10591
rect 24765 10551 24823 10557
rect 24486 10480 24492 10532
rect 24544 10520 24550 10532
rect 24780 10520 24808 10551
rect 24544 10492 24808 10520
rect 24544 10480 24550 10492
rect 12158 10452 12164 10464
rect 9631 10424 12164 10452
rect 9631 10421 9643 10424
rect 9585 10415 9643 10421
rect 12158 10412 12164 10424
rect 12216 10412 12222 10464
rect 13262 10412 13268 10464
rect 13320 10412 13326 10464
rect 19429 10455 19487 10461
rect 19429 10421 19441 10455
rect 19475 10452 19487 10455
rect 19886 10452 19892 10464
rect 19475 10424 19892 10452
rect 19475 10421 19487 10424
rect 19429 10415 19487 10421
rect 19886 10412 19892 10424
rect 19944 10412 19950 10464
rect 23382 10412 23388 10464
rect 23440 10412 23446 10464
rect 23658 10412 23664 10464
rect 23716 10452 23722 10464
rect 24213 10455 24271 10461
rect 24213 10452 24225 10455
rect 23716 10424 24225 10452
rect 23716 10412 23722 10424
rect 24213 10421 24225 10424
rect 24259 10421 24271 10455
rect 24213 10415 24271 10421
rect 1104 10362 28888 10384
rect 1104 10310 2918 10362
rect 2970 10310 2982 10362
rect 3034 10310 3046 10362
rect 3098 10310 3110 10362
rect 3162 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 10918 10362
rect 10970 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 11238 10362
rect 11290 10310 18918 10362
rect 18970 10310 18982 10362
rect 19034 10310 19046 10362
rect 19098 10310 19110 10362
rect 19162 10310 19174 10362
rect 19226 10310 19238 10362
rect 19290 10310 26918 10362
rect 26970 10310 26982 10362
rect 27034 10310 27046 10362
rect 27098 10310 27110 10362
rect 27162 10310 27174 10362
rect 27226 10310 27238 10362
rect 27290 10310 28888 10362
rect 1104 10288 28888 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 2590 10248 2596 10260
rect 1627 10220 2596 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 2590 10208 2596 10220
rect 2648 10208 2654 10260
rect 6751 10251 6809 10257
rect 6751 10217 6763 10251
rect 6797 10248 6809 10251
rect 7006 10248 7012 10260
rect 6797 10220 7012 10248
rect 6797 10217 6809 10220
rect 6751 10211 6809 10217
rect 7006 10208 7012 10220
rect 7064 10208 7070 10260
rect 7098 10208 7104 10260
rect 7156 10208 7162 10260
rect 11609 10251 11667 10257
rect 11609 10217 11621 10251
rect 11655 10248 11667 10251
rect 11790 10248 11796 10260
rect 11655 10220 11796 10248
rect 11655 10217 11667 10220
rect 11609 10211 11667 10217
rect 11790 10208 11796 10220
rect 11848 10208 11854 10260
rect 14090 10208 14096 10260
rect 14148 10208 14154 10260
rect 10778 10180 10784 10192
rect 9140 10152 10784 10180
rect 6362 10072 6368 10124
rect 6420 10112 6426 10124
rect 6420 10084 7052 10112
rect 6420 10072 6426 10084
rect 1302 10004 1308 10056
rect 1360 10044 1366 10056
rect 7024 10053 7052 10084
rect 7558 10072 7564 10124
rect 7616 10072 7622 10124
rect 7650 10072 7656 10124
rect 7708 10072 7714 10124
rect 9140 10121 9168 10152
rect 10778 10140 10784 10152
rect 10836 10180 10842 10192
rect 13446 10180 13452 10192
rect 10836 10152 13452 10180
rect 10836 10140 10842 10152
rect 13446 10140 13452 10152
rect 13504 10140 13510 10192
rect 8757 10115 8815 10121
rect 8757 10081 8769 10115
rect 8803 10112 8815 10115
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 8803 10084 9137 10112
rect 8803 10081 8815 10084
rect 8757 10075 8815 10081
rect 9125 10081 9137 10084
rect 9171 10081 9183 10115
rect 9125 10075 9183 10081
rect 12158 10072 12164 10124
rect 12216 10072 12222 10124
rect 14737 10115 14795 10121
rect 14737 10081 14749 10115
rect 14783 10112 14795 10115
rect 17862 10112 17868 10124
rect 14783 10084 17868 10112
rect 14783 10081 14795 10084
rect 14737 10075 14795 10081
rect 17862 10072 17868 10084
rect 17920 10072 17926 10124
rect 19518 10072 19524 10124
rect 19576 10112 19582 10124
rect 19705 10115 19763 10121
rect 19705 10112 19717 10115
rect 19576 10084 19717 10112
rect 19576 10072 19582 10084
rect 19705 10081 19717 10084
rect 19751 10081 19763 10115
rect 19705 10075 19763 10081
rect 19886 10072 19892 10124
rect 19944 10112 19950 10124
rect 24486 10112 24492 10124
rect 19944 10084 24492 10112
rect 19944 10072 19950 10084
rect 24486 10072 24492 10084
rect 24544 10072 24550 10124
rect 1397 10047 1455 10053
rect 1397 10044 1409 10047
rect 1360 10016 1409 10044
rect 1360 10004 1366 10016
rect 1397 10013 1409 10016
rect 1443 10044 1455 10047
rect 1673 10047 1731 10053
rect 1673 10044 1685 10047
rect 1443 10016 1685 10044
rect 1443 10013 1455 10016
rect 1397 10007 1455 10013
rect 1673 10013 1685 10016
rect 1719 10013 1731 10047
rect 1673 10007 1731 10013
rect 7009 10047 7067 10053
rect 7009 10013 7021 10047
rect 7055 10044 7067 10047
rect 9398 10044 9404 10056
rect 7055 10016 9404 10044
rect 7055 10013 7067 10016
rect 7009 10007 7067 10013
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 11977 10047 12035 10053
rect 11977 10013 11989 10047
rect 12023 10044 12035 10047
rect 13262 10044 13268 10056
rect 12023 10016 13268 10044
rect 12023 10013 12035 10016
rect 11977 10007 12035 10013
rect 13262 10004 13268 10016
rect 13320 10004 13326 10056
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10044 14519 10047
rect 15286 10044 15292 10056
rect 14507 10016 15292 10044
rect 14507 10013 14519 10016
rect 14461 10007 14519 10013
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 6270 9936 6276 9988
rect 6328 9976 6334 9988
rect 7282 9976 7288 9988
rect 6328 9948 7288 9976
rect 6328 9936 6334 9948
rect 7282 9936 7288 9948
rect 7340 9936 7346 9988
rect 7469 9979 7527 9985
rect 7469 9945 7481 9979
rect 7515 9976 7527 9979
rect 8110 9976 8116 9988
rect 7515 9948 8116 9976
rect 7515 9945 7527 9948
rect 7469 9939 7527 9945
rect 8110 9936 8116 9948
rect 8168 9976 8174 9988
rect 9309 9979 9367 9985
rect 9309 9976 9321 9979
rect 8168 9948 9321 9976
rect 8168 9936 8174 9948
rect 9309 9945 9321 9948
rect 9355 9945 9367 9979
rect 14553 9979 14611 9985
rect 14553 9976 14565 9979
rect 9309 9939 9367 9945
rect 9692 9948 14565 9976
rect 5261 9911 5319 9917
rect 5261 9877 5273 9911
rect 5307 9908 5319 9911
rect 6730 9908 6736 9920
rect 5307 9880 6736 9908
rect 5307 9877 5319 9880
rect 5261 9871 5319 9877
rect 6730 9868 6736 9880
rect 6788 9908 6794 9920
rect 8938 9908 8944 9920
rect 6788 9880 8944 9908
rect 6788 9868 6794 9880
rect 8938 9868 8944 9880
rect 8996 9908 9002 9920
rect 9692 9917 9720 9948
rect 14553 9945 14565 9948
rect 14599 9945 14611 9979
rect 14553 9939 14611 9945
rect 9217 9911 9275 9917
rect 9217 9908 9229 9911
rect 8996 9880 9229 9908
rect 8996 9868 9002 9880
rect 9217 9877 9229 9880
rect 9263 9877 9275 9911
rect 9217 9871 9275 9877
rect 9677 9911 9735 9917
rect 9677 9877 9689 9911
rect 9723 9877 9735 9911
rect 9677 9871 9735 9877
rect 12066 9868 12072 9920
rect 12124 9868 12130 9920
rect 18138 9868 18144 9920
rect 18196 9908 18202 9920
rect 19245 9911 19303 9917
rect 19245 9908 19257 9911
rect 18196 9880 19257 9908
rect 18196 9868 18202 9880
rect 19245 9877 19257 9880
rect 19291 9877 19303 9911
rect 19245 9871 19303 9877
rect 19518 9868 19524 9920
rect 19576 9908 19582 9920
rect 19613 9911 19671 9917
rect 19613 9908 19625 9911
rect 19576 9880 19625 9908
rect 19576 9868 19582 9880
rect 19613 9877 19625 9880
rect 19659 9877 19671 9911
rect 19613 9871 19671 9877
rect 1104 9818 28888 9840
rect 1104 9766 3658 9818
rect 3710 9766 3722 9818
rect 3774 9766 3786 9818
rect 3838 9766 3850 9818
rect 3902 9766 3914 9818
rect 3966 9766 3978 9818
rect 4030 9766 11658 9818
rect 11710 9766 11722 9818
rect 11774 9766 11786 9818
rect 11838 9766 11850 9818
rect 11902 9766 11914 9818
rect 11966 9766 11978 9818
rect 12030 9766 19658 9818
rect 19710 9766 19722 9818
rect 19774 9766 19786 9818
rect 19838 9766 19850 9818
rect 19902 9766 19914 9818
rect 19966 9766 19978 9818
rect 20030 9766 27658 9818
rect 27710 9766 27722 9818
rect 27774 9766 27786 9818
rect 27838 9766 27850 9818
rect 27902 9766 27914 9818
rect 27966 9766 27978 9818
rect 28030 9766 28888 9818
rect 1104 9744 28888 9766
rect 1578 9664 1584 9716
rect 1636 9664 1642 9716
rect 7006 9664 7012 9716
rect 7064 9704 7070 9716
rect 7101 9707 7159 9713
rect 7101 9704 7113 9707
rect 7064 9676 7113 9704
rect 7064 9664 7070 9676
rect 7101 9673 7113 9676
rect 7147 9673 7159 9707
rect 7101 9667 7159 9673
rect 12066 9664 12072 9716
rect 12124 9704 12130 9716
rect 12253 9707 12311 9713
rect 12253 9704 12265 9707
rect 12124 9676 12265 9704
rect 12124 9664 12130 9676
rect 12253 9673 12265 9676
rect 12299 9673 12311 9707
rect 12253 9667 12311 9673
rect 18046 9664 18052 9716
rect 18104 9704 18110 9716
rect 18104 9676 18276 9704
rect 18104 9664 18110 9676
rect 6730 9596 6736 9648
rect 6788 9596 6794 9648
rect 18138 9596 18144 9648
rect 18196 9596 18202 9648
rect 18248 9636 18276 9676
rect 19518 9664 19524 9716
rect 19576 9704 19582 9716
rect 19613 9707 19671 9713
rect 19613 9704 19625 9707
rect 19576 9676 19625 9704
rect 19576 9664 19582 9676
rect 19613 9673 19625 9676
rect 19659 9673 19671 9707
rect 19613 9667 19671 9673
rect 22465 9707 22523 9713
rect 22465 9673 22477 9707
rect 22511 9704 22523 9707
rect 23382 9704 23388 9716
rect 22511 9676 23388 9704
rect 22511 9673 22523 9676
rect 22465 9667 22523 9673
rect 23382 9664 23388 9676
rect 23440 9664 23446 9716
rect 18248 9608 18630 9636
rect 23658 9596 23664 9648
rect 23716 9596 23722 9648
rect 25130 9636 25136 9648
rect 24886 9608 25136 9636
rect 25130 9596 25136 9608
rect 25188 9596 25194 9648
rect 1302 9528 1308 9580
rect 1360 9568 1366 9580
rect 1397 9571 1455 9577
rect 1397 9568 1409 9571
rect 1360 9540 1409 9568
rect 1360 9528 1366 9540
rect 1397 9537 1409 9540
rect 1443 9568 1455 9571
rect 1673 9571 1731 9577
rect 1673 9568 1685 9571
rect 1443 9540 1685 9568
rect 1443 9537 1455 9540
rect 1397 9531 1455 9537
rect 1673 9537 1685 9540
rect 1719 9537 1731 9571
rect 7650 9568 7656 9580
rect 1673 9531 1731 9537
rect 6564 9540 7656 9568
rect 5442 9460 5448 9512
rect 5500 9500 5506 9512
rect 6564 9509 6592 9540
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 11514 9528 11520 9580
rect 11572 9568 11578 9580
rect 11885 9571 11943 9577
rect 11885 9568 11897 9571
rect 11572 9540 11897 9568
rect 11572 9528 11578 9540
rect 11885 9537 11897 9540
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 14369 9571 14427 9577
rect 14369 9537 14381 9571
rect 14415 9568 14427 9571
rect 15378 9568 15384 9580
rect 14415 9540 15384 9568
rect 14415 9537 14427 9540
rect 14369 9531 14427 9537
rect 15378 9528 15384 9540
rect 15436 9568 15442 9580
rect 15838 9568 15844 9580
rect 15436 9540 15844 9568
rect 15436 9528 15442 9540
rect 15838 9528 15844 9540
rect 15896 9528 15902 9580
rect 17310 9528 17316 9580
rect 17368 9568 17374 9580
rect 17865 9571 17923 9577
rect 17865 9568 17877 9571
rect 17368 9540 17877 9568
rect 17368 9528 17374 9540
rect 17865 9537 17877 9540
rect 17911 9537 17923 9571
rect 17865 9531 17923 9537
rect 22370 9528 22376 9580
rect 22428 9528 22434 9580
rect 6549 9503 6607 9509
rect 6549 9500 6561 9503
rect 5500 9472 6561 9500
rect 5500 9460 5506 9472
rect 6549 9469 6561 9472
rect 6595 9469 6607 9503
rect 6549 9463 6607 9469
rect 6638 9460 6644 9512
rect 6696 9460 6702 9512
rect 11609 9503 11667 9509
rect 11609 9500 11621 9503
rect 11256 9472 11621 9500
rect 7834 9324 7840 9376
rect 7892 9364 7898 9376
rect 11256 9373 11284 9472
rect 11609 9469 11621 9472
rect 11655 9469 11667 9503
rect 11609 9463 11667 9469
rect 11793 9503 11851 9509
rect 11793 9469 11805 9503
rect 11839 9500 11851 9503
rect 11974 9500 11980 9512
rect 11839 9472 11980 9500
rect 11839 9469 11851 9472
rect 11793 9463 11851 9469
rect 11624 9432 11652 9463
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 14093 9503 14151 9509
rect 14093 9469 14105 9503
rect 14139 9469 14151 9503
rect 14093 9463 14151 9469
rect 12526 9432 12532 9444
rect 11624 9404 12532 9432
rect 12526 9392 12532 9404
rect 12584 9392 12590 9444
rect 14108 9432 14136 9463
rect 14182 9460 14188 9512
rect 14240 9500 14246 9512
rect 14277 9503 14335 9509
rect 14277 9500 14289 9503
rect 14240 9472 14289 9500
rect 14240 9460 14246 9472
rect 14277 9469 14289 9472
rect 14323 9469 14335 9503
rect 14277 9463 14335 9469
rect 22002 9460 22008 9512
rect 22060 9460 22066 9512
rect 22649 9503 22707 9509
rect 22649 9469 22661 9503
rect 22695 9500 22707 9503
rect 22738 9500 22744 9512
rect 22695 9472 22744 9500
rect 22695 9469 22707 9472
rect 22649 9463 22707 9469
rect 22738 9460 22744 9472
rect 22796 9460 22802 9512
rect 23385 9503 23443 9509
rect 23385 9469 23397 9503
rect 23431 9469 23443 9503
rect 23385 9463 23443 9469
rect 14826 9432 14832 9444
rect 14108 9404 14832 9432
rect 14826 9392 14832 9404
rect 14884 9392 14890 9444
rect 21818 9392 21824 9444
rect 21876 9432 21882 9444
rect 22020 9432 22048 9460
rect 23400 9432 23428 9463
rect 25038 9460 25044 9512
rect 25096 9500 25102 9512
rect 25133 9503 25191 9509
rect 25133 9500 25145 9503
rect 25096 9472 25145 9500
rect 25096 9460 25102 9472
rect 25133 9469 25145 9472
rect 25179 9469 25191 9503
rect 25133 9463 25191 9469
rect 21876 9404 23428 9432
rect 21876 9392 21882 9404
rect 11241 9367 11299 9373
rect 11241 9364 11253 9367
rect 7892 9336 11253 9364
rect 7892 9324 7898 9336
rect 11241 9333 11253 9336
rect 11287 9333 11299 9367
rect 11241 9327 11299 9333
rect 14366 9324 14372 9376
rect 14424 9364 14430 9376
rect 14737 9367 14795 9373
rect 14737 9364 14749 9367
rect 14424 9336 14749 9364
rect 14424 9324 14430 9336
rect 14737 9333 14749 9336
rect 14783 9333 14795 9367
rect 14737 9327 14795 9333
rect 22005 9367 22063 9373
rect 22005 9333 22017 9367
rect 22051 9364 22063 9367
rect 22094 9364 22100 9376
rect 22051 9336 22100 9364
rect 22051 9333 22063 9336
rect 22005 9327 22063 9333
rect 22094 9324 22100 9336
rect 22152 9324 22158 9376
rect 1104 9274 28888 9296
rect 1104 9222 2918 9274
rect 2970 9222 2982 9274
rect 3034 9222 3046 9274
rect 3098 9222 3110 9274
rect 3162 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 10918 9274
rect 10970 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 11238 9274
rect 11290 9222 18918 9274
rect 18970 9222 18982 9274
rect 19034 9222 19046 9274
rect 19098 9222 19110 9274
rect 19162 9222 19174 9274
rect 19226 9222 19238 9274
rect 19290 9222 26918 9274
rect 26970 9222 26982 9274
rect 27034 9222 27046 9274
rect 27098 9222 27110 9274
rect 27162 9222 27174 9274
rect 27226 9222 27238 9274
rect 27290 9222 28888 9274
rect 1104 9200 28888 9222
rect 3973 9163 4031 9169
rect 3973 9129 3985 9163
rect 4019 9160 4031 9163
rect 4246 9160 4252 9172
rect 4019 9132 4252 9160
rect 4019 9129 4031 9132
rect 3973 9123 4031 9129
rect 4246 9120 4252 9132
rect 4304 9160 4310 9172
rect 5442 9160 5448 9172
rect 4304 9132 5448 9160
rect 4304 9120 4310 9132
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 7285 9163 7343 9169
rect 7285 9129 7297 9163
rect 7331 9160 7343 9163
rect 7558 9160 7564 9172
rect 7331 9132 7564 9160
rect 7331 9129 7343 9132
rect 7285 9123 7343 9129
rect 7558 9120 7564 9132
rect 7616 9120 7622 9172
rect 11974 9160 11980 9172
rect 7668 9132 11980 9160
rect 3510 9052 3516 9104
rect 3568 9092 3574 9104
rect 7668 9092 7696 9132
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 12437 9163 12495 9169
rect 12437 9129 12449 9163
rect 12483 9160 12495 9163
rect 14182 9160 14188 9172
rect 12483 9132 14188 9160
rect 12483 9129 12495 9132
rect 12437 9123 12495 9129
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 15838 9120 15844 9172
rect 15896 9120 15902 9172
rect 19334 9120 19340 9172
rect 19392 9160 19398 9172
rect 20441 9163 20499 9169
rect 20441 9160 20453 9163
rect 19392 9132 20453 9160
rect 19392 9120 19398 9132
rect 20441 9129 20453 9132
rect 20487 9129 20499 9163
rect 20441 9123 20499 9129
rect 3568 9064 7696 9092
rect 3568 9052 3574 9064
rect 6270 9024 6276 9036
rect 3160 8996 6276 9024
rect 3160 8968 3188 8996
rect 6270 8984 6276 8996
rect 6328 8984 6334 9036
rect 7193 9027 7251 9033
rect 7193 8993 7205 9027
rect 7239 9024 7251 9027
rect 7834 9024 7840 9036
rect 7239 8996 7840 9024
rect 7239 8993 7251 8996
rect 7193 8987 7251 8993
rect 7834 8984 7840 8996
rect 7892 8984 7898 9036
rect 9398 8984 9404 9036
rect 9456 9024 9462 9036
rect 9861 9027 9919 9033
rect 9861 9024 9873 9027
rect 9456 8996 9873 9024
rect 9456 8984 9462 8996
rect 9861 8993 9873 8996
rect 9907 8993 9919 9027
rect 9861 8987 9919 8993
rect 11330 8984 11336 9036
rect 11388 9024 11394 9036
rect 11793 9027 11851 9033
rect 11793 9024 11805 9027
rect 11388 8996 11805 9024
rect 11388 8984 11394 8996
rect 11793 8993 11805 8996
rect 11839 8993 11851 9027
rect 11793 8987 11851 8993
rect 11974 8984 11980 9036
rect 12032 8984 12038 9036
rect 14366 8984 14372 9036
rect 14424 8984 14430 9036
rect 1578 8916 1584 8968
rect 1636 8956 1642 8968
rect 1765 8959 1823 8965
rect 1765 8956 1777 8959
rect 1636 8928 1777 8956
rect 1636 8916 1642 8928
rect 1765 8925 1777 8928
rect 1811 8925 1823 8959
rect 1765 8919 1823 8925
rect 3142 8916 3148 8968
rect 3200 8916 3206 8968
rect 3418 8916 3424 8968
rect 3476 8956 3482 8968
rect 4157 8959 4215 8965
rect 4157 8956 4169 8959
rect 3476 8928 4169 8956
rect 3476 8916 3482 8928
rect 4157 8925 4169 8928
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 12434 8956 12440 8968
rect 11296 8928 12440 8956
rect 11296 8916 11302 8928
rect 12434 8916 12440 8928
rect 12492 8916 12498 8968
rect 14090 8916 14096 8968
rect 14148 8916 14154 8968
rect 20456 8956 20484 9123
rect 20625 8959 20683 8965
rect 20625 8956 20637 8959
rect 20456 8928 20637 8956
rect 20625 8925 20637 8928
rect 20671 8925 20683 8959
rect 20625 8919 20683 8925
rect 21266 8916 21272 8968
rect 21324 8956 21330 8968
rect 22925 8959 22983 8965
rect 22925 8956 22937 8959
rect 21324 8928 22937 8956
rect 21324 8916 21330 8928
rect 22925 8925 22937 8928
rect 22971 8925 22983 8959
rect 22925 8919 22983 8925
rect 2038 8848 2044 8900
rect 2096 8848 2102 8900
rect 3881 8891 3939 8897
rect 3881 8857 3893 8891
rect 3927 8888 3939 8891
rect 4706 8888 4712 8900
rect 3927 8860 4712 8888
rect 3927 8857 3939 8860
rect 3881 8851 3939 8857
rect 4706 8848 4712 8860
rect 4764 8888 4770 8900
rect 10137 8891 10195 8897
rect 4764 8860 9674 8888
rect 4764 8848 4770 8860
rect 1302 8780 1308 8832
rect 1360 8820 1366 8832
rect 1397 8823 1455 8829
rect 1397 8820 1409 8823
rect 1360 8792 1409 8820
rect 1360 8780 1366 8792
rect 1397 8789 1409 8792
rect 1443 8789 1455 8823
rect 1397 8783 1455 8789
rect 4338 8780 4344 8832
rect 4396 8820 4402 8832
rect 4525 8823 4583 8829
rect 4525 8820 4537 8823
rect 4396 8792 4537 8820
rect 4396 8780 4402 8792
rect 4525 8789 4537 8792
rect 4571 8789 4583 8823
rect 4525 8783 4583 8789
rect 6086 8780 6092 8832
rect 6144 8820 6150 8832
rect 7650 8820 7656 8832
rect 6144 8792 7656 8820
rect 6144 8780 6150 8792
rect 7650 8780 7656 8792
rect 7708 8780 7714 8832
rect 7742 8780 7748 8832
rect 7800 8780 7806 8832
rect 9646 8820 9674 8860
rect 10137 8857 10149 8891
rect 10183 8888 10195 8891
rect 10226 8888 10232 8900
rect 10183 8860 10232 8888
rect 10183 8857 10195 8860
rect 10137 8851 10195 8857
rect 10226 8848 10232 8860
rect 10284 8848 10290 8900
rect 12069 8891 12127 8897
rect 12069 8888 12081 8891
rect 11624 8860 12081 8888
rect 11054 8820 11060 8832
rect 9646 8792 11060 8820
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 11514 8780 11520 8832
rect 11572 8820 11578 8832
rect 11624 8829 11652 8860
rect 12069 8857 12081 8860
rect 12115 8857 12127 8891
rect 12069 8851 12127 8857
rect 15378 8848 15384 8900
rect 15436 8848 15442 8900
rect 11609 8823 11667 8829
rect 11609 8820 11621 8823
rect 11572 8792 11621 8820
rect 11572 8780 11578 8792
rect 11609 8789 11621 8792
rect 11655 8789 11667 8823
rect 11609 8783 11667 8789
rect 21818 8780 21824 8832
rect 21876 8820 21882 8832
rect 21913 8823 21971 8829
rect 21913 8820 21925 8823
rect 21876 8792 21925 8820
rect 21876 8780 21882 8792
rect 21913 8789 21925 8792
rect 21959 8789 21971 8823
rect 21913 8783 21971 8789
rect 23109 8823 23167 8829
rect 23109 8789 23121 8823
rect 23155 8820 23167 8823
rect 23382 8820 23388 8832
rect 23155 8792 23388 8820
rect 23155 8789 23167 8792
rect 23109 8783 23167 8789
rect 23382 8780 23388 8792
rect 23440 8780 23446 8832
rect 1104 8730 28888 8752
rect 1104 8678 3658 8730
rect 3710 8678 3722 8730
rect 3774 8678 3786 8730
rect 3838 8678 3850 8730
rect 3902 8678 3914 8730
rect 3966 8678 3978 8730
rect 4030 8678 11658 8730
rect 11710 8678 11722 8730
rect 11774 8678 11786 8730
rect 11838 8678 11850 8730
rect 11902 8678 11914 8730
rect 11966 8678 11978 8730
rect 12030 8678 19658 8730
rect 19710 8678 19722 8730
rect 19774 8678 19786 8730
rect 19838 8678 19850 8730
rect 19902 8678 19914 8730
rect 19966 8678 19978 8730
rect 20030 8678 27658 8730
rect 27710 8678 27722 8730
rect 27774 8678 27786 8730
rect 27838 8678 27850 8730
rect 27902 8678 27914 8730
rect 27966 8678 27978 8730
rect 28030 8678 28888 8730
rect 1104 8656 28888 8678
rect 2038 8576 2044 8628
rect 2096 8616 2102 8628
rect 2593 8619 2651 8625
rect 2593 8616 2605 8619
rect 2096 8588 2605 8616
rect 2096 8576 2102 8588
rect 2593 8585 2605 8588
rect 2639 8585 2651 8619
rect 2593 8579 2651 8585
rect 2961 8619 3019 8625
rect 2961 8585 2973 8619
rect 3007 8616 3019 8619
rect 3510 8616 3516 8628
rect 3007 8588 3516 8616
rect 3007 8585 3019 8588
rect 2961 8579 3019 8585
rect 3510 8576 3516 8588
rect 3568 8576 3574 8628
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8616 4307 8619
rect 6638 8616 6644 8628
rect 4295 8588 6644 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 7929 8619 7987 8625
rect 7929 8616 7941 8619
rect 7800 8588 7941 8616
rect 7800 8576 7806 8588
rect 7929 8585 7941 8588
rect 7975 8585 7987 8619
rect 7929 8579 7987 8585
rect 10226 8576 10232 8628
rect 10284 8576 10290 8628
rect 10597 8619 10655 8625
rect 10597 8585 10609 8619
rect 10643 8616 10655 8619
rect 11514 8616 11520 8628
rect 10643 8588 11520 8616
rect 10643 8585 10655 8588
rect 10597 8579 10655 8585
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 17310 8576 17316 8628
rect 17368 8616 17374 8628
rect 20809 8619 20867 8625
rect 20809 8616 20821 8619
rect 17368 8588 20821 8616
rect 17368 8576 17374 8588
rect 20809 8585 20821 8588
rect 20855 8585 20867 8619
rect 20809 8579 20867 8585
rect 24305 8619 24363 8625
rect 24305 8585 24317 8619
rect 24351 8616 24363 8619
rect 24394 8616 24400 8628
rect 24351 8588 24400 8616
rect 24351 8585 24363 8588
rect 24305 8579 24363 8585
rect 24394 8576 24400 8588
rect 24452 8576 24458 8628
rect 7650 8508 7656 8560
rect 7708 8548 7714 8560
rect 8021 8551 8079 8557
rect 8021 8548 8033 8551
rect 7708 8520 8033 8548
rect 7708 8508 7714 8520
rect 8021 8517 8033 8520
rect 8067 8517 8079 8551
rect 8021 8511 8079 8517
rect 19426 8508 19432 8560
rect 19484 8548 19490 8560
rect 19521 8551 19579 8557
rect 19521 8548 19533 8551
rect 19484 8520 19533 8548
rect 19484 8508 19490 8520
rect 19521 8517 19533 8520
rect 19567 8517 19579 8551
rect 19521 8511 19579 8517
rect 22094 8508 22100 8560
rect 22152 8508 22158 8560
rect 23382 8548 23388 8560
rect 23322 8520 23388 8548
rect 23382 8508 23388 8520
rect 23440 8548 23446 8560
rect 25130 8548 25136 8560
rect 23440 8520 25136 8548
rect 23440 8508 23446 8520
rect 25130 8508 25136 8520
rect 25188 8508 25194 8560
rect 1302 8440 1308 8492
rect 1360 8480 1366 8492
rect 1397 8483 1455 8489
rect 1397 8480 1409 8483
rect 1360 8452 1409 8480
rect 1360 8440 1366 8452
rect 1397 8449 1409 8452
rect 1443 8449 1455 8483
rect 1397 8443 1455 8449
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3694 8480 3700 8492
rect 3099 8452 3700 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 3786 8440 3792 8492
rect 3844 8440 3850 8492
rect 3878 8440 3884 8492
rect 3936 8440 3942 8492
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 4341 8483 4399 8489
rect 4341 8480 4353 8483
rect 4212 8452 4353 8480
rect 4212 8440 4218 8452
rect 4341 8449 4353 8452
rect 4387 8449 4399 8483
rect 11330 8480 11336 8492
rect 4341 8443 4399 8449
rect 7852 8452 11336 8480
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8412 1731 8415
rect 2774 8412 2780 8424
rect 1719 8384 2780 8412
rect 1719 8381 1731 8384
rect 1673 8375 1731 8381
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8381 3295 8415
rect 3237 8375 3295 8381
rect 3605 8415 3663 8421
rect 3605 8381 3617 8415
rect 3651 8412 3663 8415
rect 7190 8412 7196 8424
rect 3651 8384 7196 8412
rect 3651 8381 3663 8384
rect 3605 8375 3663 8381
rect 3142 8344 3148 8356
rect 2792 8316 3148 8344
rect 2792 8288 2820 8316
rect 3142 8304 3148 8316
rect 3200 8304 3206 8356
rect 3252 8344 3280 8375
rect 4246 8344 4252 8356
rect 3252 8316 4252 8344
rect 4246 8304 4252 8316
rect 4304 8304 4310 8356
rect 4540 8353 4568 8384
rect 7190 8372 7196 8384
rect 7248 8372 7254 8424
rect 7852 8421 7880 8452
rect 11330 8440 11336 8452
rect 11388 8480 11394 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 11388 8452 11529 8480
rect 11388 8440 11394 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 18046 8440 18052 8492
rect 18104 8440 18110 8492
rect 24397 8483 24455 8489
rect 24397 8449 24409 8483
rect 24443 8480 24455 8483
rect 24762 8480 24768 8492
rect 24443 8452 24768 8480
rect 24443 8449 24455 8452
rect 24397 8443 24455 8449
rect 24762 8440 24768 8452
rect 24820 8440 24826 8492
rect 7837 8415 7895 8421
rect 7837 8412 7849 8415
rect 7484 8384 7849 8412
rect 4525 8347 4583 8353
rect 4525 8313 4537 8347
rect 4571 8313 4583 8347
rect 4525 8307 4583 8313
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7484 8353 7512 8384
rect 7837 8381 7849 8384
rect 7883 8381 7895 8415
rect 10689 8415 10747 8421
rect 10689 8412 10701 8415
rect 7837 8375 7895 8381
rect 8404 8384 10701 8412
rect 8404 8353 8432 8384
rect 10689 8381 10701 8384
rect 10735 8381 10747 8415
rect 10689 8375 10747 8381
rect 10873 8415 10931 8421
rect 10873 8381 10885 8415
rect 10919 8412 10931 8415
rect 11054 8412 11060 8424
rect 10919 8384 11060 8412
rect 10919 8381 10931 8384
rect 10873 8375 10931 8381
rect 11054 8372 11060 8384
rect 11112 8412 11118 8424
rect 12158 8412 12164 8424
rect 11112 8384 12164 8412
rect 11112 8372 11118 8384
rect 12158 8372 12164 8384
rect 12216 8372 12222 8424
rect 17681 8415 17739 8421
rect 17681 8381 17693 8415
rect 17727 8412 17739 8415
rect 18782 8412 18788 8424
rect 17727 8384 18788 8412
rect 17727 8381 17739 8384
rect 17681 8375 17739 8381
rect 18782 8372 18788 8384
rect 18840 8372 18846 8424
rect 19153 8415 19211 8421
rect 19153 8381 19165 8415
rect 19199 8412 19211 8415
rect 19429 8415 19487 8421
rect 19199 8384 19380 8412
rect 19199 8381 19211 8384
rect 19153 8375 19211 8381
rect 7469 8347 7527 8353
rect 7469 8344 7481 8347
rect 6972 8316 7481 8344
rect 6972 8304 6978 8316
rect 7469 8313 7481 8316
rect 7515 8313 7527 8347
rect 7469 8307 7527 8313
rect 8389 8347 8447 8353
rect 8389 8313 8401 8347
rect 8435 8313 8447 8347
rect 19352 8344 19380 8384
rect 19429 8381 19441 8415
rect 19475 8412 19487 8415
rect 21818 8412 21824 8424
rect 19475 8384 21824 8412
rect 19475 8381 19487 8384
rect 19429 8375 19487 8381
rect 21818 8372 21824 8384
rect 21876 8372 21882 8424
rect 24213 8415 24271 8421
rect 24213 8381 24225 8415
rect 24259 8412 24271 8415
rect 24486 8412 24492 8424
rect 24259 8384 24492 8412
rect 24259 8381 24271 8384
rect 24213 8375 24271 8381
rect 24486 8372 24492 8384
rect 24544 8372 24550 8424
rect 19518 8344 19524 8356
rect 19352 8316 19524 8344
rect 8389 8307 8447 8313
rect 19518 8304 19524 8316
rect 19576 8304 19582 8356
rect 23382 8304 23388 8356
rect 23440 8344 23446 8356
rect 23569 8347 23627 8353
rect 23569 8344 23581 8347
rect 23440 8316 23581 8344
rect 23440 8304 23446 8316
rect 23569 8313 23581 8316
rect 23615 8313 23627 8347
rect 23569 8307 23627 8313
rect 2774 8236 2780 8288
rect 2832 8236 2838 8288
rect 14550 8236 14556 8288
rect 14608 8276 14614 8288
rect 16758 8276 16764 8288
rect 14608 8248 16764 8276
rect 14608 8236 14614 8248
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 24670 8236 24676 8288
rect 24728 8276 24734 8288
rect 24765 8279 24823 8285
rect 24765 8276 24777 8279
rect 24728 8248 24777 8276
rect 24728 8236 24734 8248
rect 24765 8245 24777 8248
rect 24811 8245 24823 8279
rect 24765 8239 24823 8245
rect 1104 8186 28888 8208
rect 1104 8134 2918 8186
rect 2970 8134 2982 8186
rect 3034 8134 3046 8186
rect 3098 8134 3110 8186
rect 3162 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 10918 8186
rect 10970 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 11238 8186
rect 11290 8134 18918 8186
rect 18970 8134 18982 8186
rect 19034 8134 19046 8186
rect 19098 8134 19110 8186
rect 19162 8134 19174 8186
rect 19226 8134 19238 8186
rect 19290 8134 26918 8186
rect 26970 8134 26982 8186
rect 27034 8134 27046 8186
rect 27098 8134 27110 8186
rect 27162 8134 27174 8186
rect 27226 8134 27238 8186
rect 27290 8134 28888 8186
rect 1104 8112 28888 8134
rect 3694 8032 3700 8084
rect 3752 8072 3758 8084
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 3752 8044 3801 8072
rect 3752 8032 3758 8044
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 3789 8035 3847 8041
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 8205 8075 8263 8081
rect 8205 8072 8217 8075
rect 7800 8044 8217 8072
rect 7800 8032 7806 8044
rect 8205 8041 8217 8044
rect 8251 8041 8263 8075
rect 17589 8075 17647 8081
rect 17589 8072 17601 8075
rect 8205 8035 8263 8041
rect 15948 8044 17601 8072
rect 2501 8007 2559 8013
rect 2501 7973 2513 8007
rect 2547 8004 2559 8007
rect 4154 8004 4160 8016
rect 2547 7976 4160 8004
rect 2547 7973 2559 7976
rect 2501 7967 2559 7973
rect 4154 7964 4160 7976
rect 4212 7964 4218 8016
rect 4430 8004 4436 8016
rect 4264 7976 4436 8004
rect 1302 7896 1308 7948
rect 1360 7936 1366 7948
rect 1397 7939 1455 7945
rect 1397 7936 1409 7939
rect 1360 7908 1409 7936
rect 1360 7896 1366 7908
rect 1397 7905 1409 7908
rect 1443 7905 1455 7939
rect 1397 7899 1455 7905
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 4264 7936 4292 7976
rect 4430 7964 4436 7976
rect 4488 7964 4494 8016
rect 1719 7908 4292 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 4338 7896 4344 7948
rect 4396 7936 4402 7948
rect 4709 7939 4767 7945
rect 4709 7936 4721 7939
rect 4396 7908 4721 7936
rect 4396 7896 4402 7908
rect 4709 7905 4721 7908
rect 4755 7936 4767 7939
rect 7098 7936 7104 7948
rect 4755 7908 7104 7936
rect 4755 7905 4767 7908
rect 4709 7899 4767 7905
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 1210 7828 1216 7880
rect 1268 7868 1274 7880
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 1268 7840 2329 7868
rect 1268 7828 1274 7840
rect 2317 7837 2329 7840
rect 2363 7868 2375 7871
rect 2593 7871 2651 7877
rect 2593 7868 2605 7871
rect 2363 7840 2605 7868
rect 2363 7837 2375 7840
rect 2317 7831 2375 7837
rect 2593 7837 2605 7840
rect 2639 7837 2651 7871
rect 2593 7831 2651 7837
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 6457 7871 6515 7877
rect 6457 7868 6469 7871
rect 4120 7840 6469 7868
rect 4120 7828 4126 7840
rect 6457 7837 6469 7840
rect 6503 7837 6515 7871
rect 15948 7854 15976 8044
rect 17589 8041 17601 8044
rect 17635 8072 17647 8075
rect 18046 8072 18052 8084
rect 17635 8044 18052 8072
rect 17635 8041 17647 8044
rect 17589 8035 17647 8041
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 19334 8032 19340 8084
rect 19392 8032 19398 8084
rect 19518 8032 19524 8084
rect 19576 8032 19582 8084
rect 20438 8032 20444 8084
rect 20496 8072 20502 8084
rect 27893 8075 27951 8081
rect 27893 8072 27905 8075
rect 20496 8044 27905 8072
rect 20496 8032 20502 8044
rect 27893 8041 27905 8044
rect 27939 8041 27951 8075
rect 27893 8035 27951 8041
rect 17862 7964 17868 8016
rect 17920 8004 17926 8016
rect 17957 8007 18015 8013
rect 17957 8004 17969 8007
rect 17920 7976 17969 8004
rect 17920 7964 17926 7976
rect 17957 7973 17969 7976
rect 18003 8004 18015 8007
rect 19886 8004 19892 8016
rect 18003 7976 19892 8004
rect 18003 7973 18015 7976
rect 17957 7967 18015 7973
rect 19886 7964 19892 7976
rect 19944 7964 19950 8016
rect 19996 7976 20300 8004
rect 17310 7896 17316 7948
rect 17368 7936 17374 7948
rect 17368 7908 18184 7936
rect 17368 7896 17374 7908
rect 17773 7871 17831 7877
rect 6457 7831 6515 7837
rect 17773 7837 17785 7871
rect 17819 7868 17831 7871
rect 17954 7868 17960 7880
rect 17819 7840 17960 7868
rect 17819 7837 17831 7840
rect 17773 7831 17831 7837
rect 3510 7760 3516 7812
rect 3568 7800 3574 7812
rect 3786 7800 3792 7812
rect 3568 7772 3792 7800
rect 3568 7760 3574 7772
rect 3786 7760 3792 7772
rect 3844 7800 3850 7812
rect 4249 7803 4307 7809
rect 4249 7800 4261 7803
rect 3844 7772 4261 7800
rect 3844 7760 3850 7772
rect 4249 7769 4261 7772
rect 4295 7769 4307 7803
rect 4249 7763 4307 7769
rect 3878 7692 3884 7744
rect 3936 7732 3942 7744
rect 4154 7732 4160 7744
rect 3936 7704 4160 7732
rect 3936 7692 3942 7704
rect 4154 7692 4160 7704
rect 4212 7692 4218 7744
rect 6472 7732 6500 7831
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 18156 7877 18184 7908
rect 18690 7896 18696 7948
rect 18748 7936 18754 7948
rect 19996 7936 20024 7976
rect 18748 7908 20024 7936
rect 18748 7896 18754 7908
rect 20070 7896 20076 7948
rect 20128 7896 20134 7948
rect 20272 7936 20300 7976
rect 20530 7964 20536 8016
rect 20588 8004 20594 8016
rect 20588 7976 21312 8004
rect 20588 7964 20594 7976
rect 21284 7945 21312 7976
rect 20901 7939 20959 7945
rect 20901 7936 20913 7939
rect 20272 7908 20913 7936
rect 20901 7905 20913 7908
rect 20947 7905 20959 7939
rect 20901 7899 20959 7905
rect 21269 7939 21327 7945
rect 21269 7905 21281 7939
rect 21315 7905 21327 7939
rect 21269 7899 21327 7905
rect 24670 7896 24676 7948
rect 24728 7896 24734 7948
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7837 18199 7871
rect 18141 7831 18199 7837
rect 19610 7828 19616 7880
rect 19668 7868 19674 7880
rect 20809 7871 20867 7877
rect 20809 7868 20821 7871
rect 19668 7840 20821 7868
rect 19668 7828 19674 7840
rect 20809 7837 20821 7840
rect 20855 7868 20867 7871
rect 21453 7871 21511 7877
rect 21453 7868 21465 7871
rect 20855 7840 21465 7868
rect 20855 7837 20867 7840
rect 20809 7831 20867 7837
rect 21453 7837 21465 7840
rect 21499 7837 21511 7871
rect 21453 7831 21511 7837
rect 21818 7828 21824 7880
rect 21876 7868 21882 7880
rect 24394 7868 24400 7880
rect 21876 7840 24400 7868
rect 21876 7828 21882 7840
rect 24394 7828 24400 7840
rect 24452 7828 24458 7880
rect 27908 7868 27936 8035
rect 28077 7871 28135 7877
rect 28077 7868 28089 7871
rect 27908 7840 28089 7868
rect 28077 7837 28089 7840
rect 28123 7837 28135 7871
rect 28077 7831 28135 7837
rect 6730 7760 6736 7812
rect 6788 7760 6794 7812
rect 7282 7760 7288 7812
rect 7340 7760 7346 7812
rect 17034 7760 17040 7812
rect 17092 7760 17098 7812
rect 17494 7760 17500 7812
rect 17552 7800 17558 7812
rect 20717 7803 20775 7809
rect 17552 7772 20484 7800
rect 17552 7760 17558 7772
rect 6914 7732 6920 7744
rect 6472 7704 6920 7732
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 15565 7735 15623 7741
rect 15565 7701 15577 7735
rect 15611 7732 15623 7735
rect 16942 7732 16948 7744
rect 15611 7704 16948 7732
rect 15611 7701 15623 7704
rect 15565 7695 15623 7701
rect 16942 7692 16948 7704
rect 17000 7692 17006 7744
rect 18782 7692 18788 7744
rect 18840 7732 18846 7744
rect 19518 7732 19524 7744
rect 18840 7704 19524 7732
rect 18840 7692 18846 7704
rect 19518 7692 19524 7704
rect 19576 7732 19582 7744
rect 19889 7735 19947 7741
rect 19889 7732 19901 7735
rect 19576 7704 19901 7732
rect 19576 7692 19582 7704
rect 19889 7701 19901 7704
rect 19935 7701 19947 7735
rect 19889 7695 19947 7701
rect 19981 7735 20039 7741
rect 19981 7701 19993 7735
rect 20027 7732 20039 7735
rect 20349 7735 20407 7741
rect 20349 7732 20361 7735
rect 20027 7704 20361 7732
rect 20027 7701 20039 7704
rect 19981 7695 20039 7701
rect 20349 7701 20361 7704
rect 20395 7701 20407 7735
rect 20456 7732 20484 7772
rect 20717 7769 20729 7803
rect 20763 7800 20775 7803
rect 21545 7803 21603 7809
rect 21545 7800 21557 7803
rect 20763 7772 21557 7800
rect 20763 7769 20775 7772
rect 20717 7763 20775 7769
rect 21545 7769 21557 7772
rect 21591 7800 21603 7803
rect 22370 7800 22376 7812
rect 21591 7772 22376 7800
rect 21591 7769 21603 7772
rect 21545 7763 21603 7769
rect 22370 7760 22376 7772
rect 22428 7800 22434 7812
rect 23382 7800 23388 7812
rect 22428 7772 23388 7800
rect 22428 7760 22434 7772
rect 23382 7760 23388 7772
rect 23440 7760 23446 7812
rect 25130 7760 25136 7812
rect 25188 7760 25194 7812
rect 28350 7760 28356 7812
rect 28408 7760 28414 7812
rect 21266 7732 21272 7744
rect 20456 7704 21272 7732
rect 20349 7695 20407 7701
rect 21266 7692 21272 7704
rect 21324 7692 21330 7744
rect 21913 7735 21971 7741
rect 21913 7701 21925 7735
rect 21959 7732 21971 7735
rect 22278 7732 22284 7744
rect 21959 7704 22284 7732
rect 21959 7701 21971 7704
rect 21913 7695 21971 7701
rect 22278 7692 22284 7704
rect 22336 7692 22342 7744
rect 24762 7692 24768 7744
rect 24820 7732 24826 7744
rect 26145 7735 26203 7741
rect 26145 7732 26157 7735
rect 24820 7704 26157 7732
rect 24820 7692 24826 7704
rect 26145 7701 26157 7704
rect 26191 7701 26203 7735
rect 26145 7695 26203 7701
rect 1104 7642 28888 7664
rect 1104 7590 3658 7642
rect 3710 7590 3722 7642
rect 3774 7590 3786 7642
rect 3838 7590 3850 7642
rect 3902 7590 3914 7642
rect 3966 7590 3978 7642
rect 4030 7590 11658 7642
rect 11710 7590 11722 7642
rect 11774 7590 11786 7642
rect 11838 7590 11850 7642
rect 11902 7590 11914 7642
rect 11966 7590 11978 7642
rect 12030 7590 19658 7642
rect 19710 7590 19722 7642
rect 19774 7590 19786 7642
rect 19838 7590 19850 7642
rect 19902 7590 19914 7642
rect 19966 7590 19978 7642
rect 20030 7590 27658 7642
rect 27710 7590 27722 7642
rect 27774 7590 27786 7642
rect 27838 7590 27850 7642
rect 27902 7590 27914 7642
rect 27966 7590 27978 7642
rect 28030 7590 28888 7642
rect 1104 7568 28888 7590
rect 1302 7488 1308 7540
rect 1360 7528 1366 7540
rect 1397 7531 1455 7537
rect 1397 7528 1409 7531
rect 1360 7500 1409 7528
rect 1360 7488 1366 7500
rect 1397 7497 1409 7500
rect 1443 7497 1455 7531
rect 1397 7491 1455 7497
rect 1578 7488 1584 7540
rect 1636 7528 1642 7540
rect 3326 7528 3332 7540
rect 1636 7500 3332 7528
rect 1636 7488 1642 7500
rect 3326 7488 3332 7500
rect 3384 7528 3390 7540
rect 4062 7528 4068 7540
rect 3384 7500 4068 7528
rect 3384 7488 3390 7500
rect 4062 7488 4068 7500
rect 4120 7528 4126 7540
rect 4120 7500 4384 7528
rect 4120 7488 4126 7500
rect 2590 7420 2596 7472
rect 2648 7420 2654 7472
rect 3602 7420 3608 7472
rect 3660 7460 3666 7472
rect 3660 7432 4016 7460
rect 3660 7420 3666 7432
rect 1578 7352 1584 7404
rect 1636 7352 1642 7404
rect 3510 7352 3516 7404
rect 3568 7392 3574 7404
rect 3789 7395 3847 7401
rect 3789 7392 3801 7395
rect 3568 7364 3801 7392
rect 3568 7352 3574 7364
rect 1857 7327 1915 7333
rect 1857 7293 1869 7327
rect 1903 7324 1915 7327
rect 1903 7296 3464 7324
rect 1903 7293 1915 7296
rect 1857 7287 1915 7293
rect 3436 7265 3464 7296
rect 3421 7259 3479 7265
rect 3421 7225 3433 7259
rect 3467 7225 3479 7259
rect 3421 7219 3479 7225
rect 3329 7191 3387 7197
rect 3329 7157 3341 7191
rect 3375 7188 3387 7191
rect 3712 7188 3740 7364
rect 3789 7361 3801 7364
rect 3835 7361 3847 7395
rect 3789 7355 3847 7361
rect 3988 7333 4016 7432
rect 4356 7401 4384 7500
rect 6730 7488 6736 7540
rect 6788 7528 6794 7540
rect 7193 7531 7251 7537
rect 7193 7528 7205 7531
rect 6788 7500 7205 7528
rect 6788 7488 6794 7500
rect 7193 7497 7205 7500
rect 7239 7497 7251 7531
rect 7193 7491 7251 7497
rect 7561 7531 7619 7537
rect 7561 7497 7573 7531
rect 7607 7528 7619 7531
rect 7742 7528 7748 7540
rect 7607 7500 7748 7528
rect 7607 7497 7619 7500
rect 7561 7491 7619 7497
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 8846 7488 8852 7540
rect 8904 7488 8910 7540
rect 14737 7531 14795 7537
rect 14737 7497 14749 7531
rect 14783 7528 14795 7531
rect 14783 7500 15332 7528
rect 14783 7497 14795 7500
rect 14737 7491 14795 7497
rect 5626 7420 5632 7472
rect 5684 7420 5690 7472
rect 14826 7420 14832 7472
rect 14884 7420 14890 7472
rect 15304 7469 15332 7500
rect 15378 7488 15384 7540
rect 15436 7488 15442 7540
rect 16669 7531 16727 7537
rect 16669 7497 16681 7531
rect 16715 7528 16727 7531
rect 17034 7528 17040 7540
rect 16715 7500 17040 7528
rect 16715 7497 16727 7500
rect 16669 7491 16727 7497
rect 17034 7488 17040 7500
rect 17092 7488 17098 7540
rect 17129 7531 17187 7537
rect 17129 7497 17141 7531
rect 17175 7528 17187 7531
rect 18417 7531 18475 7537
rect 18417 7528 18429 7531
rect 17175 7500 18429 7528
rect 17175 7497 17187 7500
rect 17129 7491 17187 7497
rect 18417 7497 18429 7500
rect 18463 7497 18475 7531
rect 18417 7491 18475 7497
rect 18782 7488 18788 7540
rect 18840 7528 18846 7540
rect 18877 7531 18935 7537
rect 18877 7528 18889 7531
rect 18840 7500 18889 7528
rect 18840 7488 18846 7500
rect 18877 7497 18889 7500
rect 18923 7497 18935 7531
rect 18877 7491 18935 7497
rect 24762 7488 24768 7540
rect 24820 7528 24826 7540
rect 24857 7531 24915 7537
rect 24857 7528 24869 7531
rect 24820 7500 24869 7528
rect 24820 7488 24826 7500
rect 24857 7497 24869 7500
rect 24903 7497 24915 7531
rect 24857 7491 24915 7497
rect 24949 7531 25007 7537
rect 24949 7497 24961 7531
rect 24995 7528 25007 7531
rect 25038 7528 25044 7540
rect 24995 7500 25044 7528
rect 24995 7497 25007 7500
rect 24949 7491 25007 7497
rect 15289 7463 15347 7469
rect 15289 7429 15301 7463
rect 15335 7460 15347 7463
rect 17494 7460 17500 7472
rect 15335 7432 17500 7460
rect 15335 7429 15347 7432
rect 15289 7423 15347 7429
rect 17494 7420 17500 7432
rect 17552 7420 17558 7472
rect 21634 7420 21640 7472
rect 21692 7460 21698 7472
rect 24029 7463 24087 7469
rect 21692 7432 22586 7460
rect 21692 7420 21698 7432
rect 24029 7429 24041 7463
rect 24075 7460 24087 7463
rect 24780 7460 24808 7488
rect 24075 7432 24808 7460
rect 24075 7429 24087 7432
rect 24029 7423 24087 7429
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7361 4399 7395
rect 14550 7392 14556 7404
rect 4341 7355 4399 7361
rect 14384 7364 14556 7392
rect 3881 7327 3939 7333
rect 3881 7293 3893 7327
rect 3927 7293 3939 7327
rect 3881 7287 3939 7293
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7293 4031 7327
rect 3973 7287 4031 7293
rect 3375 7160 3740 7188
rect 3896 7188 3924 7287
rect 4614 7284 4620 7336
rect 4672 7284 4678 7336
rect 7650 7284 7656 7336
rect 7708 7284 7714 7336
rect 7834 7284 7840 7336
rect 7892 7284 7898 7336
rect 5994 7188 6000 7200
rect 3896 7160 6000 7188
rect 3375 7157 3387 7160
rect 3329 7151 3387 7157
rect 5994 7148 6000 7160
rect 6052 7148 6058 7200
rect 6086 7148 6092 7200
rect 6144 7148 6150 7200
rect 14182 7148 14188 7200
rect 14240 7188 14246 7200
rect 14384 7197 14412 7364
rect 14550 7352 14556 7364
rect 14608 7352 14614 7404
rect 15013 7395 15071 7401
rect 15013 7361 15025 7395
rect 15059 7361 15071 7395
rect 15013 7355 15071 7361
rect 15028 7324 15056 7355
rect 15562 7352 15568 7404
rect 15620 7392 15626 7404
rect 15841 7395 15899 7401
rect 15841 7392 15853 7395
rect 15620 7364 15853 7392
rect 15620 7352 15626 7364
rect 15841 7361 15853 7364
rect 15887 7361 15899 7395
rect 15841 7355 15899 7361
rect 16942 7352 16948 7404
rect 17000 7392 17006 7404
rect 17037 7395 17095 7401
rect 17037 7392 17049 7395
rect 17000 7364 17049 7392
rect 17000 7352 17006 7364
rect 17037 7361 17049 7364
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 18785 7395 18843 7401
rect 18785 7361 18797 7395
rect 18831 7392 18843 7395
rect 19610 7392 19616 7404
rect 18831 7364 19616 7392
rect 18831 7361 18843 7364
rect 18785 7355 18843 7361
rect 19610 7352 19616 7364
rect 19668 7352 19674 7404
rect 24121 7395 24179 7401
rect 24121 7361 24133 7395
rect 24167 7392 24179 7395
rect 24964 7392 24992 7491
rect 25038 7488 25044 7500
rect 25096 7488 25102 7540
rect 24167 7364 24992 7392
rect 24167 7361 24179 7364
rect 24121 7355 24179 7361
rect 17313 7327 17371 7333
rect 15028 7296 15792 7324
rect 15764 7265 15792 7296
rect 17313 7293 17325 7327
rect 17359 7324 17371 7327
rect 17862 7324 17868 7336
rect 17359 7296 17868 7324
rect 17359 7293 17371 7296
rect 17313 7287 17371 7293
rect 17862 7284 17868 7296
rect 17920 7284 17926 7336
rect 18690 7284 18696 7336
rect 18748 7324 18754 7336
rect 18969 7327 19027 7333
rect 18969 7324 18981 7327
rect 18748 7296 18981 7324
rect 18748 7284 18754 7296
rect 18969 7293 18981 7296
rect 19015 7293 19027 7327
rect 18969 7287 19027 7293
rect 21358 7284 21364 7336
rect 21416 7324 21422 7336
rect 21818 7324 21824 7336
rect 21416 7296 21824 7324
rect 21416 7284 21422 7296
rect 21818 7284 21824 7296
rect 21876 7284 21882 7336
rect 22094 7284 22100 7336
rect 22152 7284 22158 7336
rect 24210 7284 24216 7336
rect 24268 7284 24274 7336
rect 24578 7284 24584 7336
rect 24636 7324 24642 7336
rect 24762 7324 24768 7336
rect 24636 7296 24768 7324
rect 24636 7284 24642 7296
rect 24762 7284 24768 7296
rect 24820 7324 24826 7336
rect 25041 7327 25099 7333
rect 25041 7324 25053 7327
rect 24820 7296 25053 7324
rect 24820 7284 24826 7296
rect 25041 7293 25053 7296
rect 25087 7293 25099 7327
rect 25041 7287 25099 7293
rect 15749 7259 15807 7265
rect 15749 7225 15761 7259
rect 15795 7256 15807 7259
rect 17954 7256 17960 7268
rect 15795 7228 17960 7256
rect 15795 7225 15807 7228
rect 15749 7219 15807 7225
rect 17954 7216 17960 7228
rect 18012 7216 18018 7268
rect 14369 7191 14427 7197
rect 14369 7188 14381 7191
rect 14240 7160 14381 7188
rect 14240 7148 14246 7160
rect 14369 7157 14381 7160
rect 14415 7157 14427 7191
rect 14369 7151 14427 7157
rect 22554 7148 22560 7200
rect 22612 7188 22618 7200
rect 23569 7191 23627 7197
rect 23569 7188 23581 7191
rect 22612 7160 23581 7188
rect 22612 7148 22618 7160
rect 23569 7157 23581 7160
rect 23615 7157 23627 7191
rect 23569 7151 23627 7157
rect 23658 7148 23664 7200
rect 23716 7148 23722 7200
rect 24489 7191 24547 7197
rect 24489 7157 24501 7191
rect 24535 7188 24547 7191
rect 24670 7188 24676 7200
rect 24535 7160 24676 7188
rect 24535 7157 24547 7160
rect 24489 7151 24547 7157
rect 24670 7148 24676 7160
rect 24728 7148 24734 7200
rect 1104 7098 28888 7120
rect 1104 7046 2918 7098
rect 2970 7046 2982 7098
rect 3034 7046 3046 7098
rect 3098 7046 3110 7098
rect 3162 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 10918 7098
rect 10970 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 11238 7098
rect 11290 7046 18918 7098
rect 18970 7046 18982 7098
rect 19034 7046 19046 7098
rect 19098 7046 19110 7098
rect 19162 7046 19174 7098
rect 19226 7046 19238 7098
rect 19290 7046 26918 7098
rect 26970 7046 26982 7098
rect 27034 7046 27046 7098
rect 27098 7046 27110 7098
rect 27162 7046 27174 7098
rect 27226 7046 27238 7098
rect 27290 7046 28888 7098
rect 1104 7024 28888 7046
rect 4614 6944 4620 6996
rect 4672 6984 4678 6996
rect 4801 6987 4859 6993
rect 4801 6984 4813 6987
rect 4672 6956 4813 6984
rect 4672 6944 4678 6956
rect 4801 6953 4813 6956
rect 4847 6953 4859 6987
rect 4801 6947 4859 6953
rect 22094 6944 22100 6996
rect 22152 6984 22158 6996
rect 22189 6987 22247 6993
rect 22189 6984 22201 6987
rect 22152 6956 22201 6984
rect 22152 6944 22158 6956
rect 22189 6953 22201 6956
rect 22235 6953 22247 6987
rect 22189 6947 22247 6953
rect 1949 6919 2007 6925
rect 1949 6885 1961 6919
rect 1995 6885 2007 6919
rect 1949 6879 2007 6885
rect 1964 6848 1992 6879
rect 2682 6876 2688 6928
rect 2740 6916 2746 6928
rect 2774 6916 2780 6928
rect 2740 6888 2780 6916
rect 2740 6876 2746 6888
rect 2774 6876 2780 6888
rect 2832 6876 2838 6928
rect 3418 6848 3424 6860
rect 1964 6820 3424 6848
rect 3418 6808 3424 6820
rect 3476 6808 3482 6860
rect 5442 6808 5448 6860
rect 5500 6808 5506 6860
rect 6914 6808 6920 6860
rect 6972 6848 6978 6860
rect 7009 6851 7067 6857
rect 7009 6848 7021 6851
rect 6972 6820 7021 6848
rect 6972 6808 6978 6820
rect 7009 6817 7021 6820
rect 7055 6817 7067 6851
rect 13081 6851 13139 6857
rect 13081 6848 13093 6851
rect 7009 6811 7067 6817
rect 10980 6820 13093 6848
rect 1302 6740 1308 6792
rect 1360 6780 1366 6792
rect 1765 6783 1823 6789
rect 1765 6780 1777 6783
rect 1360 6752 1777 6780
rect 1360 6740 1366 6752
rect 1765 6749 1777 6752
rect 1811 6780 1823 6783
rect 2225 6783 2283 6789
rect 2225 6780 2237 6783
rect 1811 6752 2237 6780
rect 1811 6749 1823 6752
rect 1765 6743 1823 6749
rect 2225 6749 2237 6752
rect 2271 6749 2283 6783
rect 2225 6743 2283 6749
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6780 5227 6783
rect 6086 6780 6092 6792
rect 5215 6752 6092 6780
rect 5215 6749 5227 6752
rect 5169 6743 5227 6749
rect 6086 6740 6092 6752
rect 6144 6740 6150 6792
rect 10980 6789 11008 6820
rect 13081 6817 13093 6820
rect 13127 6848 13139 6851
rect 13814 6848 13820 6860
rect 13127 6820 13820 6848
rect 13127 6817 13139 6820
rect 13081 6811 13139 6817
rect 13814 6808 13820 6820
rect 13872 6848 13878 6860
rect 14090 6848 14096 6860
rect 13872 6820 14096 6848
rect 13872 6808 13878 6820
rect 14090 6808 14096 6820
rect 14148 6808 14154 6860
rect 19518 6808 19524 6860
rect 19576 6848 19582 6860
rect 19705 6851 19763 6857
rect 19705 6848 19717 6851
rect 19576 6820 19717 6848
rect 19576 6808 19582 6820
rect 19705 6817 19717 6820
rect 19751 6817 19763 6851
rect 19705 6811 19763 6817
rect 19889 6851 19947 6857
rect 19889 6817 19901 6851
rect 19935 6848 19947 6851
rect 20530 6848 20536 6860
rect 19935 6820 20536 6848
rect 19935 6817 19947 6820
rect 19889 6811 19947 6817
rect 10689 6783 10747 6789
rect 10689 6749 10701 6783
rect 10735 6780 10747 6783
rect 10965 6783 11023 6789
rect 10965 6780 10977 6783
rect 10735 6752 10977 6780
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 10965 6749 10977 6752
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 11330 6740 11336 6792
rect 11388 6780 11394 6792
rect 11388 6752 11560 6780
rect 11388 6740 11394 6752
rect 11532 6724 11560 6752
rect 19334 6740 19340 6792
rect 19392 6780 19398 6792
rect 19904 6780 19932 6811
rect 20530 6808 20536 6820
rect 20588 6808 20594 6860
rect 22002 6808 22008 6860
rect 22060 6848 22066 6860
rect 22738 6848 22744 6860
rect 22060 6820 22744 6848
rect 22060 6808 22066 6820
rect 22738 6808 22744 6820
rect 22796 6808 22802 6860
rect 19392 6752 19932 6780
rect 19392 6740 19398 6752
rect 22554 6740 22560 6792
rect 22612 6740 22618 6792
rect 22649 6783 22707 6789
rect 22649 6749 22661 6783
rect 22695 6780 22707 6783
rect 23658 6780 23664 6792
rect 22695 6752 23664 6780
rect 22695 6749 22707 6752
rect 22649 6743 22707 6749
rect 23658 6740 23664 6752
rect 23716 6740 23722 6792
rect 1210 6672 1216 6724
rect 1268 6712 1274 6724
rect 1489 6715 1547 6721
rect 1489 6712 1501 6715
rect 1268 6684 1501 6712
rect 1268 6672 1274 6684
rect 1489 6681 1501 6684
rect 1535 6681 1547 6715
rect 1489 6675 1547 6681
rect 1673 6715 1731 6721
rect 1673 6681 1685 6715
rect 1719 6712 1731 6715
rect 2041 6715 2099 6721
rect 2041 6712 2053 6715
rect 1719 6684 2053 6712
rect 1719 6681 1731 6684
rect 1673 6675 1731 6681
rect 2041 6681 2053 6684
rect 2087 6712 2099 6715
rect 3418 6712 3424 6724
rect 2087 6684 3424 6712
rect 2087 6681 2099 6684
rect 2041 6675 2099 6681
rect 1504 6644 1532 6675
rect 3418 6672 3424 6684
rect 3476 6672 3482 6724
rect 8754 6672 8760 6724
rect 8812 6672 8818 6724
rect 8846 6672 8852 6724
rect 8904 6712 8910 6724
rect 8904 6684 9246 6712
rect 8904 6672 8910 6684
rect 10318 6672 10324 6724
rect 10376 6712 10382 6724
rect 10413 6715 10471 6721
rect 10413 6712 10425 6715
rect 10376 6684 10425 6712
rect 10376 6672 10382 6684
rect 10413 6681 10425 6684
rect 10459 6681 10471 6715
rect 10413 6675 10471 6681
rect 11514 6672 11520 6724
rect 11572 6712 11578 6724
rect 11572 6684 11638 6712
rect 11572 6672 11578 6684
rect 12802 6672 12808 6724
rect 12860 6672 12866 6724
rect 13722 6672 13728 6724
rect 13780 6672 13786 6724
rect 14366 6672 14372 6724
rect 14424 6672 14430 6724
rect 15378 6672 15384 6724
rect 15436 6672 15442 6724
rect 19610 6672 19616 6724
rect 19668 6712 19674 6724
rect 22572 6712 22600 6740
rect 19668 6684 22600 6712
rect 19668 6672 19674 6684
rect 2409 6647 2467 6653
rect 2409 6644 2421 6647
rect 1504 6616 2421 6644
rect 2409 6613 2421 6616
rect 2455 6613 2467 6647
rect 2409 6607 2467 6613
rect 5261 6647 5319 6653
rect 5261 6613 5273 6647
rect 5307 6644 5319 6647
rect 5534 6644 5540 6656
rect 5307 6616 5540 6644
rect 5307 6613 5319 6616
rect 5261 6607 5319 6613
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 8018 6604 8024 6656
rect 8076 6644 8082 6656
rect 8941 6647 8999 6653
rect 8941 6644 8953 6647
rect 8076 6616 8953 6644
rect 8076 6604 8082 6616
rect 8941 6613 8953 6616
rect 8987 6613 8999 6647
rect 8941 6607 8999 6613
rect 11330 6604 11336 6656
rect 11388 6604 11394 6656
rect 13817 6647 13875 6653
rect 13817 6613 13829 6647
rect 13863 6644 13875 6647
rect 14090 6644 14096 6656
rect 13863 6616 14096 6644
rect 13863 6613 13875 6616
rect 13817 6607 13875 6613
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 14734 6604 14740 6656
rect 14792 6644 14798 6656
rect 15841 6647 15899 6653
rect 15841 6644 15853 6647
rect 14792 6616 15853 6644
rect 14792 6604 14798 6616
rect 15841 6613 15853 6616
rect 15887 6613 15899 6647
rect 15841 6607 15899 6613
rect 18506 6604 18512 6656
rect 18564 6644 18570 6656
rect 19245 6647 19303 6653
rect 19245 6644 19257 6647
rect 18564 6616 19257 6644
rect 18564 6604 18570 6616
rect 19245 6613 19257 6616
rect 19291 6613 19303 6647
rect 19245 6607 19303 6613
rect 1104 6554 28888 6576
rect 1104 6502 3658 6554
rect 3710 6502 3722 6554
rect 3774 6502 3786 6554
rect 3838 6502 3850 6554
rect 3902 6502 3914 6554
rect 3966 6502 3978 6554
rect 4030 6502 11658 6554
rect 11710 6502 11722 6554
rect 11774 6502 11786 6554
rect 11838 6502 11850 6554
rect 11902 6502 11914 6554
rect 11966 6502 11978 6554
rect 12030 6502 19658 6554
rect 19710 6502 19722 6554
rect 19774 6502 19786 6554
rect 19838 6502 19850 6554
rect 19902 6502 19914 6554
rect 19966 6502 19978 6554
rect 20030 6502 27658 6554
rect 27710 6502 27722 6554
rect 27774 6502 27786 6554
rect 27838 6502 27850 6554
rect 27902 6502 27914 6554
rect 27966 6502 27978 6554
rect 28030 6502 28888 6554
rect 1104 6480 28888 6502
rect 7650 6400 7656 6452
rect 7708 6440 7714 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 7708 6412 7849 6440
rect 7708 6400 7714 6412
rect 7837 6409 7849 6412
rect 7883 6409 7895 6443
rect 7837 6403 7895 6409
rect 8754 6400 8760 6452
rect 8812 6440 8818 6452
rect 8849 6443 8907 6449
rect 8849 6440 8861 6443
rect 8812 6412 8861 6440
rect 8812 6400 8818 6412
rect 8849 6409 8861 6412
rect 8895 6440 8907 6443
rect 11422 6440 11428 6452
rect 8895 6412 11428 6440
rect 8895 6409 8907 6412
rect 8849 6403 8907 6409
rect 11422 6400 11428 6412
rect 11480 6440 11486 6452
rect 11480 6412 11560 6440
rect 11480 6400 11486 6412
rect 6914 6332 6920 6384
rect 6972 6372 6978 6384
rect 7101 6375 7159 6381
rect 7101 6372 7113 6375
rect 6972 6344 7113 6372
rect 6972 6332 6978 6344
rect 7101 6341 7113 6344
rect 7147 6341 7159 6375
rect 7101 6335 7159 6341
rect 7190 6332 7196 6384
rect 7248 6372 7254 6384
rect 8110 6372 8116 6384
rect 7248 6344 8116 6372
rect 7248 6332 7254 6344
rect 8110 6332 8116 6344
rect 8168 6372 8174 6384
rect 9582 6372 9588 6384
rect 8168 6344 9588 6372
rect 8168 6332 8174 6344
rect 9582 6332 9588 6344
rect 9640 6372 9646 6384
rect 11532 6381 11560 6412
rect 14366 6400 14372 6452
rect 14424 6400 14430 6452
rect 14734 6400 14740 6452
rect 14792 6400 14798 6452
rect 14829 6443 14887 6449
rect 14829 6409 14841 6443
rect 14875 6440 14887 6443
rect 16669 6443 16727 6449
rect 16669 6440 16681 6443
rect 14875 6412 16681 6440
rect 14875 6409 14887 6412
rect 14829 6403 14887 6409
rect 16669 6409 16681 6412
rect 16715 6409 16727 6443
rect 16669 6403 16727 6409
rect 16942 6400 16948 6452
rect 17000 6440 17006 6452
rect 17129 6443 17187 6449
rect 17129 6440 17141 6443
rect 17000 6412 17141 6440
rect 17000 6400 17006 6412
rect 17129 6409 17141 6412
rect 17175 6409 17187 6443
rect 17129 6403 17187 6409
rect 20898 6400 20904 6452
rect 20956 6440 20962 6452
rect 21177 6443 21235 6449
rect 21177 6440 21189 6443
rect 20956 6412 21189 6440
rect 20956 6400 20962 6412
rect 21177 6409 21189 6412
rect 21223 6440 21235 6443
rect 21634 6440 21640 6452
rect 21223 6412 21640 6440
rect 21223 6409 21235 6412
rect 21177 6403 21235 6409
rect 21634 6400 21640 6412
rect 21692 6400 21698 6452
rect 11517 6375 11575 6381
rect 9640 6344 11376 6372
rect 9640 6332 9646 6344
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 1489 6307 1547 6313
rect 1489 6304 1501 6307
rect 1360 6276 1501 6304
rect 1360 6264 1366 6276
rect 1489 6273 1501 6276
rect 1535 6304 1547 6307
rect 1949 6307 2007 6313
rect 1949 6304 1961 6307
rect 1535 6276 1961 6304
rect 1535 6273 1547 6276
rect 1489 6267 1547 6273
rect 1949 6273 1961 6276
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 8202 6264 8208 6316
rect 8260 6264 8266 6316
rect 9953 6307 10011 6313
rect 9953 6304 9965 6307
rect 8312 6276 9965 6304
rect 3237 6239 3295 6245
rect 3237 6205 3249 6239
rect 3283 6236 3295 6239
rect 3602 6236 3608 6248
rect 3283 6208 3608 6236
rect 3283 6205 3295 6208
rect 3237 6199 3295 6205
rect 3602 6196 3608 6208
rect 3660 6236 3666 6248
rect 3660 6208 6868 6236
rect 3660 6196 3666 6208
rect 1673 6171 1731 6177
rect 1673 6137 1685 6171
rect 1719 6168 1731 6171
rect 1857 6171 1915 6177
rect 1857 6168 1869 6171
rect 1719 6140 1869 6168
rect 1719 6137 1731 6140
rect 1673 6131 1731 6137
rect 1857 6137 1869 6140
rect 1903 6168 1915 6171
rect 6178 6168 6184 6180
rect 1903 6140 6184 6168
rect 1903 6137 1915 6140
rect 1857 6131 1915 6137
rect 6178 6128 6184 6140
rect 6236 6128 6242 6180
rect 3694 6060 3700 6112
rect 3752 6060 3758 6112
rect 6840 6100 6868 6208
rect 8018 6196 8024 6248
rect 8076 6236 8082 6248
rect 8312 6245 8340 6276
rect 9953 6273 9965 6276
rect 9999 6273 10011 6307
rect 9953 6267 10011 6273
rect 10686 6264 10692 6316
rect 10744 6304 10750 6316
rect 10965 6307 11023 6313
rect 10965 6304 10977 6307
rect 10744 6276 10977 6304
rect 10744 6264 10750 6276
rect 10965 6273 10977 6276
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 8297 6239 8355 6245
rect 8297 6236 8309 6239
rect 8076 6208 8309 6236
rect 8076 6196 8082 6208
rect 8297 6205 8309 6208
rect 8343 6205 8355 6239
rect 8297 6199 8355 6205
rect 8481 6239 8539 6245
rect 8481 6205 8493 6239
rect 8527 6236 8539 6239
rect 9493 6239 9551 6245
rect 8527 6208 8984 6236
rect 8527 6205 8539 6208
rect 8481 6199 8539 6205
rect 7098 6128 7104 6180
rect 7156 6168 7162 6180
rect 7745 6171 7803 6177
rect 7745 6168 7757 6171
rect 7156 6140 7757 6168
rect 7156 6128 7162 6140
rect 7745 6137 7757 6140
rect 7791 6168 7803 6171
rect 8496 6168 8524 6199
rect 7791 6140 8524 6168
rect 7791 6137 7803 6140
rect 7745 6131 7803 6137
rect 8846 6100 8852 6112
rect 6840 6072 8852 6100
rect 8846 6060 8852 6072
rect 8904 6060 8910 6112
rect 8956 6100 8984 6208
rect 9493 6205 9505 6239
rect 9539 6236 9551 6239
rect 9766 6236 9772 6248
rect 9539 6208 9772 6236
rect 9539 6205 9551 6208
rect 9493 6199 9551 6205
rect 9766 6196 9772 6208
rect 9824 6196 9830 6248
rect 9861 6239 9919 6245
rect 9861 6205 9873 6239
rect 9907 6236 9919 6239
rect 11057 6239 11115 6245
rect 9907 6208 10640 6236
rect 9907 6205 9919 6208
rect 9861 6199 9919 6205
rect 10318 6128 10324 6180
rect 10376 6128 10382 6180
rect 10612 6177 10640 6208
rect 11057 6205 11069 6239
rect 11103 6205 11115 6239
rect 11057 6199 11115 6205
rect 11241 6239 11299 6245
rect 11241 6205 11253 6239
rect 11287 6236 11299 6239
rect 11348 6236 11376 6344
rect 11517 6341 11529 6375
rect 11563 6372 11575 6375
rect 13357 6375 13415 6381
rect 13357 6372 13369 6375
rect 11563 6344 13369 6372
rect 11563 6341 11575 6344
rect 11517 6335 11575 6341
rect 13357 6341 13369 6344
rect 13403 6341 13415 6375
rect 13357 6335 13415 6341
rect 14001 6375 14059 6381
rect 14001 6341 14013 6375
rect 14047 6372 14059 6375
rect 14752 6372 14780 6400
rect 14047 6344 14780 6372
rect 14844 6344 17356 6372
rect 14047 6341 14059 6344
rect 14001 6335 14059 6341
rect 13265 6307 13323 6313
rect 13265 6273 13277 6307
rect 13311 6304 13323 6307
rect 13814 6304 13820 6316
rect 13311 6276 13820 6304
rect 13311 6273 13323 6276
rect 13265 6267 13323 6273
rect 13814 6264 13820 6276
rect 13872 6264 13878 6316
rect 13906 6264 13912 6316
rect 13964 6264 13970 6316
rect 14090 6264 14096 6316
rect 14148 6304 14154 6316
rect 14844 6304 14872 6344
rect 14148 6276 14872 6304
rect 15197 6307 15255 6313
rect 14148 6264 14154 6276
rect 13722 6236 13728 6248
rect 11287 6208 13728 6236
rect 11287 6205 11299 6208
rect 11241 6199 11299 6205
rect 10597 6171 10655 6177
rect 10597 6137 10609 6171
rect 10643 6137 10655 6171
rect 11072 6168 11100 6199
rect 13722 6196 13728 6208
rect 13780 6196 13786 6248
rect 14200 6245 14228 6276
rect 15197 6273 15209 6307
rect 15243 6273 15255 6307
rect 15197 6267 15255 6273
rect 14185 6239 14243 6245
rect 14185 6205 14197 6239
rect 14231 6205 14243 6239
rect 14185 6199 14243 6205
rect 14826 6196 14832 6248
rect 14884 6236 14890 6248
rect 14921 6239 14979 6245
rect 14921 6236 14933 6239
rect 14884 6208 14933 6236
rect 14884 6196 14890 6208
rect 14921 6205 14933 6208
rect 14967 6205 14979 6239
rect 14921 6199 14979 6205
rect 11330 6168 11336 6180
rect 11072 6140 11336 6168
rect 10597 6131 10655 6137
rect 11330 6128 11336 6140
rect 11388 6128 11394 6180
rect 15212 6168 15240 6267
rect 17034 6264 17040 6316
rect 17092 6264 17098 6316
rect 17328 6245 17356 6344
rect 21266 6332 21272 6384
rect 21324 6332 21330 6384
rect 17313 6239 17371 6245
rect 17313 6205 17325 6239
rect 17359 6236 17371 6239
rect 18690 6236 18696 6248
rect 17359 6208 18696 6236
rect 17359 6205 17371 6208
rect 17313 6199 17371 6205
rect 18690 6196 18696 6208
rect 18748 6196 18754 6248
rect 15565 6171 15623 6177
rect 15565 6168 15577 6171
rect 12406 6140 15577 6168
rect 10778 6100 10784 6112
rect 8956 6072 10784 6100
rect 10778 6060 10784 6072
rect 10836 6100 10842 6112
rect 12406 6100 12434 6140
rect 15565 6137 15577 6140
rect 15611 6137 15623 6171
rect 15565 6131 15623 6137
rect 10836 6072 12434 6100
rect 10836 6060 10842 6072
rect 12710 6060 12716 6112
rect 12768 6100 12774 6112
rect 13541 6103 13599 6109
rect 13541 6100 13553 6103
rect 12768 6072 13553 6100
rect 12768 6060 12774 6072
rect 13541 6069 13553 6072
rect 13587 6069 13599 6103
rect 13541 6063 13599 6069
rect 15381 6103 15439 6109
rect 15381 6069 15393 6103
rect 15427 6100 15439 6103
rect 16666 6100 16672 6112
rect 15427 6072 16672 6100
rect 15427 6069 15439 6072
rect 15381 6063 15439 6069
rect 16666 6060 16672 6072
rect 16724 6060 16730 6112
rect 1104 6010 28888 6032
rect 1104 5958 2918 6010
rect 2970 5958 2982 6010
rect 3034 5958 3046 6010
rect 3098 5958 3110 6010
rect 3162 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 10918 6010
rect 10970 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 11238 6010
rect 11290 5958 18918 6010
rect 18970 5958 18982 6010
rect 19034 5958 19046 6010
rect 19098 5958 19110 6010
rect 19162 5958 19174 6010
rect 19226 5958 19238 6010
rect 19290 5958 26918 6010
rect 26970 5958 26982 6010
rect 27034 5958 27046 6010
rect 27098 5958 27110 6010
rect 27162 5958 27174 6010
rect 27226 5958 27238 6010
rect 27290 5958 28888 6010
rect 1104 5936 28888 5958
rect 2961 5899 3019 5905
rect 2961 5865 2973 5899
rect 3007 5896 3019 5899
rect 3050 5896 3056 5908
rect 3007 5868 3056 5896
rect 3007 5865 3019 5868
rect 2961 5859 3019 5865
rect 3050 5856 3056 5868
rect 3108 5896 3114 5908
rect 3602 5896 3608 5908
rect 3108 5868 3608 5896
rect 3108 5856 3114 5868
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 5534 5856 5540 5908
rect 5592 5856 5598 5908
rect 5994 5856 6000 5908
rect 6052 5896 6058 5908
rect 7561 5899 7619 5905
rect 7561 5896 7573 5899
rect 6052 5868 7573 5896
rect 6052 5856 6058 5868
rect 7561 5865 7573 5868
rect 7607 5865 7619 5899
rect 7561 5859 7619 5865
rect 9766 5856 9772 5908
rect 9824 5896 9830 5908
rect 12158 5896 12164 5908
rect 9824 5868 12164 5896
rect 9824 5856 9830 5868
rect 12158 5856 12164 5868
rect 12216 5856 12222 5908
rect 12253 5899 12311 5905
rect 12253 5865 12265 5899
rect 12299 5896 12311 5899
rect 12802 5896 12808 5908
rect 12299 5868 12808 5896
rect 12299 5865 12311 5868
rect 12253 5859 12311 5865
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 17954 5856 17960 5908
rect 18012 5896 18018 5908
rect 18012 5868 21864 5896
rect 18012 5856 18018 5868
rect 2225 5831 2283 5837
rect 2225 5797 2237 5831
rect 2271 5828 2283 5831
rect 2409 5831 2467 5837
rect 2409 5828 2421 5831
rect 2271 5800 2421 5828
rect 2271 5797 2283 5800
rect 2225 5791 2283 5797
rect 2409 5797 2421 5800
rect 2455 5828 2467 5831
rect 2685 5831 2743 5837
rect 2685 5828 2697 5831
rect 2455 5800 2697 5828
rect 2455 5797 2467 5800
rect 2409 5791 2467 5797
rect 2685 5797 2697 5800
rect 2731 5828 2743 5831
rect 6086 5828 6092 5840
rect 2731 5800 6092 5828
rect 2731 5797 2743 5800
rect 2685 5791 2743 5797
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 1397 5695 1455 5701
rect 1397 5692 1409 5695
rect 1360 5664 1409 5692
rect 1360 5652 1366 5664
rect 1397 5661 1409 5664
rect 1443 5692 1455 5695
rect 1673 5695 1731 5701
rect 1673 5692 1685 5695
rect 1443 5664 1685 5692
rect 1443 5661 1455 5664
rect 1397 5655 1455 5661
rect 1673 5661 1685 5664
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 2498 5652 2504 5704
rect 2556 5652 2562 5704
rect 2792 5701 2820 5800
rect 6086 5788 6092 5800
rect 6144 5788 6150 5840
rect 11606 5828 11612 5840
rect 6196 5800 11612 5828
rect 4985 5763 5043 5769
rect 4985 5729 4997 5763
rect 5031 5760 5043 5763
rect 5718 5760 5724 5772
rect 5031 5732 5724 5760
rect 5031 5729 5043 5732
rect 4985 5723 5043 5729
rect 5718 5720 5724 5732
rect 5776 5720 5782 5772
rect 6196 5760 6224 5800
rect 11606 5788 11612 5800
rect 11664 5788 11670 5840
rect 5828 5732 6224 5760
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 3513 5695 3571 5701
rect 3513 5661 3525 5695
rect 3559 5692 3571 5695
rect 3694 5692 3700 5704
rect 3559 5664 3700 5692
rect 3559 5661 3571 5664
rect 3513 5655 3571 5661
rect 3694 5652 3700 5664
rect 3752 5692 3758 5704
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 3752 5664 4077 5692
rect 3752 5652 3758 5664
rect 4065 5661 4077 5664
rect 4111 5692 4123 5695
rect 4433 5695 4491 5701
rect 4433 5692 4445 5695
rect 4111 5664 4445 5692
rect 4111 5661 4123 5664
rect 4065 5655 4123 5661
rect 4433 5661 4445 5664
rect 4479 5692 4491 5695
rect 5828 5692 5856 5732
rect 8018 5720 8024 5772
rect 8076 5720 8082 5772
rect 8110 5720 8116 5772
rect 8168 5720 8174 5772
rect 10778 5720 10784 5772
rect 10836 5760 10842 5772
rect 11425 5763 11483 5769
rect 11425 5760 11437 5763
rect 10836 5732 11437 5760
rect 10836 5720 10842 5732
rect 11425 5729 11437 5732
rect 11471 5729 11483 5763
rect 12176 5760 12204 5856
rect 14090 5788 14096 5840
rect 14148 5788 14154 5840
rect 14734 5828 14740 5840
rect 14568 5800 14740 5828
rect 14568 5769 14596 5800
rect 14734 5788 14740 5800
rect 14792 5788 14798 5840
rect 14826 5788 14832 5840
rect 14884 5828 14890 5840
rect 17218 5828 17224 5840
rect 14884 5800 17224 5828
rect 14884 5788 14890 5800
rect 17218 5788 17224 5800
rect 17276 5828 17282 5840
rect 17276 5800 18644 5828
rect 17276 5788 17282 5800
rect 12805 5763 12863 5769
rect 12805 5760 12817 5763
rect 12176 5732 12817 5760
rect 11425 5723 11483 5729
rect 12805 5729 12817 5732
rect 12851 5729 12863 5763
rect 12805 5723 12863 5729
rect 14553 5763 14611 5769
rect 14553 5729 14565 5763
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 14645 5763 14703 5769
rect 14645 5729 14657 5763
rect 14691 5760 14703 5763
rect 16666 5760 16672 5772
rect 14691 5732 16672 5760
rect 14691 5729 14703 5732
rect 14645 5723 14703 5729
rect 16666 5720 16672 5732
rect 16724 5760 16730 5772
rect 16724 5732 18092 5760
rect 16724 5720 16730 5732
rect 4479 5664 5856 5692
rect 7929 5695 7987 5701
rect 4479 5661 4491 5664
rect 4433 5655 4491 5661
rect 7929 5661 7941 5695
rect 7975 5692 7987 5695
rect 8202 5692 8208 5704
rect 7975 5664 8208 5692
rect 7975 5661 7987 5664
rect 7929 5655 7987 5661
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 11330 5652 11336 5704
rect 11388 5692 11394 5704
rect 12621 5695 12679 5701
rect 12621 5692 12633 5695
rect 11388 5664 12633 5692
rect 11388 5652 11394 5664
rect 12621 5661 12633 5664
rect 12667 5661 12679 5695
rect 12621 5655 12679 5661
rect 12710 5652 12716 5704
rect 12768 5652 12774 5704
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 14461 5695 14519 5701
rect 14461 5692 14473 5695
rect 13964 5664 14473 5692
rect 13964 5652 13970 5664
rect 14461 5661 14473 5664
rect 14507 5661 14519 5695
rect 14461 5655 14519 5661
rect 16485 5695 16543 5701
rect 16485 5661 16497 5695
rect 16531 5692 16543 5695
rect 16942 5692 16948 5704
rect 16531 5664 16948 5692
rect 16531 5661 16543 5664
rect 16485 5655 16543 5661
rect 16942 5652 16948 5664
rect 17000 5652 17006 5704
rect 18064 5692 18092 5732
rect 18506 5720 18512 5772
rect 18564 5720 18570 5772
rect 18616 5769 18644 5800
rect 18601 5763 18659 5769
rect 18601 5729 18613 5763
rect 18647 5729 18659 5763
rect 18601 5723 18659 5729
rect 21358 5720 21364 5772
rect 21416 5760 21422 5772
rect 21637 5763 21695 5769
rect 21637 5760 21649 5763
rect 21416 5732 21649 5760
rect 21416 5720 21422 5732
rect 21637 5729 21649 5732
rect 21683 5729 21695 5763
rect 21637 5723 21695 5729
rect 19334 5692 19340 5704
rect 18064 5664 19340 5692
rect 19334 5652 19340 5664
rect 19392 5652 19398 5704
rect 21836 5701 21864 5868
rect 21821 5695 21879 5701
rect 21821 5661 21833 5695
rect 21867 5661 21879 5695
rect 21821 5655 21879 5661
rect 3329 5627 3387 5633
rect 3329 5624 3341 5627
rect 1596 5596 3341 5624
rect 1596 5565 1624 5596
rect 3329 5593 3341 5596
rect 3375 5593 3387 5627
rect 4249 5627 4307 5633
rect 4249 5624 4261 5627
rect 3329 5587 3387 5593
rect 3896 5596 4261 5624
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5525 1639 5559
rect 1581 5519 1639 5525
rect 3234 5516 3240 5568
rect 3292 5556 3298 5568
rect 3896 5565 3924 5596
rect 4249 5593 4261 5596
rect 4295 5624 4307 5627
rect 4295 5596 6040 5624
rect 4295 5593 4307 5596
rect 4249 5587 4307 5593
rect 3881 5559 3939 5565
rect 3881 5556 3893 5559
rect 3292 5528 3893 5556
rect 3292 5516 3298 5528
rect 3881 5525 3893 5528
rect 3927 5525 3939 5559
rect 3881 5519 3939 5525
rect 4982 5516 4988 5568
rect 5040 5556 5046 5568
rect 5077 5559 5135 5565
rect 5077 5556 5089 5559
rect 5040 5528 5089 5556
rect 5040 5516 5046 5528
rect 5077 5525 5089 5528
rect 5123 5525 5135 5559
rect 5077 5519 5135 5525
rect 5166 5516 5172 5568
rect 5224 5516 5230 5568
rect 5718 5516 5724 5568
rect 5776 5516 5782 5568
rect 6012 5556 6040 5596
rect 6086 5584 6092 5636
rect 6144 5624 6150 5636
rect 14182 5624 14188 5636
rect 6144 5596 14188 5624
rect 6144 5584 6150 5596
rect 14182 5584 14188 5596
rect 14240 5584 14246 5636
rect 16393 5627 16451 5633
rect 16393 5593 16405 5627
rect 16439 5624 16451 5627
rect 17034 5624 17040 5636
rect 16439 5596 17040 5624
rect 16439 5593 16451 5596
rect 16393 5587 16451 5593
rect 17034 5584 17040 5596
rect 17092 5624 17098 5636
rect 17092 5596 19932 5624
rect 17092 5584 17098 5596
rect 9766 5556 9772 5568
rect 6012 5528 9772 5556
rect 9766 5516 9772 5528
rect 9824 5516 9830 5568
rect 10870 5516 10876 5568
rect 10928 5516 10934 5568
rect 10962 5516 10968 5568
rect 11020 5556 11026 5568
rect 11241 5559 11299 5565
rect 11241 5556 11253 5559
rect 11020 5528 11253 5556
rect 11020 5516 11026 5528
rect 11241 5525 11253 5528
rect 11287 5556 11299 5559
rect 11330 5556 11336 5568
rect 11287 5528 11336 5556
rect 11287 5525 11299 5528
rect 11241 5519 11299 5525
rect 11330 5516 11336 5528
rect 11388 5516 11394 5568
rect 11606 5516 11612 5568
rect 11664 5556 11670 5568
rect 15562 5556 15568 5568
rect 11664 5528 15568 5556
rect 11664 5516 11670 5528
rect 15562 5516 15568 5528
rect 15620 5516 15626 5568
rect 16022 5516 16028 5568
rect 16080 5516 16086 5568
rect 17954 5516 17960 5568
rect 18012 5556 18018 5568
rect 18049 5559 18107 5565
rect 18049 5556 18061 5559
rect 18012 5528 18061 5556
rect 18012 5516 18018 5528
rect 18049 5525 18061 5528
rect 18095 5525 18107 5559
rect 18049 5519 18107 5525
rect 18414 5516 18420 5568
rect 18472 5516 18478 5568
rect 19904 5565 19932 5596
rect 20898 5584 20904 5636
rect 20956 5584 20962 5636
rect 21361 5627 21419 5633
rect 21361 5593 21373 5627
rect 21407 5624 21419 5627
rect 21450 5624 21456 5636
rect 21407 5596 21456 5624
rect 21407 5593 21419 5596
rect 21361 5587 21419 5593
rect 21450 5584 21456 5596
rect 21508 5584 21514 5636
rect 22002 5584 22008 5636
rect 22060 5584 22066 5636
rect 19889 5559 19947 5565
rect 19889 5525 19901 5559
rect 19935 5556 19947 5559
rect 21174 5556 21180 5568
rect 19935 5528 21180 5556
rect 19935 5525 19947 5528
rect 19889 5519 19947 5525
rect 21174 5516 21180 5528
rect 21232 5516 21238 5568
rect 1104 5466 28888 5488
rect 1104 5414 3658 5466
rect 3710 5414 3722 5466
rect 3774 5414 3786 5466
rect 3838 5414 3850 5466
rect 3902 5414 3914 5466
rect 3966 5414 3978 5466
rect 4030 5414 11658 5466
rect 11710 5414 11722 5466
rect 11774 5414 11786 5466
rect 11838 5414 11850 5466
rect 11902 5414 11914 5466
rect 11966 5414 11978 5466
rect 12030 5414 19658 5466
rect 19710 5414 19722 5466
rect 19774 5414 19786 5466
rect 19838 5414 19850 5466
rect 19902 5414 19914 5466
rect 19966 5414 19978 5466
rect 20030 5414 27658 5466
rect 27710 5414 27722 5466
rect 27774 5414 27786 5466
rect 27838 5414 27850 5466
rect 27902 5414 27914 5466
rect 27966 5414 27978 5466
rect 28030 5414 28888 5466
rect 1104 5392 28888 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 2498 5352 2504 5364
rect 1627 5324 2504 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 2498 5312 2504 5324
rect 2556 5312 2562 5364
rect 2682 5312 2688 5364
rect 2740 5312 2746 5364
rect 3237 5355 3295 5361
rect 3237 5321 3249 5355
rect 3283 5352 3295 5355
rect 3283 5324 3648 5352
rect 3283 5321 3295 5324
rect 3237 5315 3295 5321
rect 2133 5287 2191 5293
rect 2133 5253 2145 5287
rect 2179 5284 2191 5287
rect 2700 5284 2728 5312
rect 3620 5293 3648 5324
rect 3694 5312 3700 5364
rect 3752 5352 3758 5364
rect 5169 5355 5227 5361
rect 3752 5324 4936 5352
rect 3752 5312 3758 5324
rect 3605 5287 3663 5293
rect 2179 5256 2728 5284
rect 2884 5256 3556 5284
rect 2179 5253 2191 5256
rect 2133 5247 2191 5253
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 1360 5188 1409 5216
rect 1360 5176 1366 5188
rect 1397 5185 1409 5188
rect 1443 5216 1455 5219
rect 1673 5219 1731 5225
rect 1673 5216 1685 5219
rect 1443 5188 1685 5216
rect 1443 5185 1455 5188
rect 1397 5179 1455 5185
rect 1673 5185 1685 5188
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 2240 5012 2268 5256
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5216 2743 5219
rect 2884 5216 2912 5256
rect 2731 5188 2912 5216
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 2317 5083 2375 5089
rect 2317 5049 2329 5083
rect 2363 5080 2375 5083
rect 2590 5080 2596 5092
rect 2363 5052 2596 5080
rect 2363 5049 2375 5052
rect 2317 5043 2375 5049
rect 2590 5040 2596 5052
rect 2648 5080 2654 5092
rect 2774 5080 2780 5092
rect 2648 5052 2780 5080
rect 2648 5040 2654 5052
rect 2774 5040 2780 5052
rect 2832 5040 2838 5092
rect 2884 5089 2912 5188
rect 3050 5176 3056 5228
rect 3108 5176 3114 5228
rect 3234 5176 3240 5228
rect 3292 5216 3298 5228
rect 3421 5219 3479 5225
rect 3421 5216 3433 5219
rect 3292 5188 3433 5216
rect 3292 5176 3298 5188
rect 3421 5185 3433 5188
rect 3467 5185 3479 5219
rect 3528 5216 3556 5256
rect 3605 5253 3617 5287
rect 3651 5284 3663 5287
rect 4706 5284 4712 5296
rect 3651 5256 4712 5284
rect 3651 5253 3663 5256
rect 3605 5247 3663 5253
rect 4706 5244 4712 5256
rect 4764 5244 4770 5296
rect 4246 5216 4252 5228
rect 3528 5188 4252 5216
rect 3421 5179 3479 5185
rect 3436 5148 3464 5179
rect 4246 5176 4252 5188
rect 4304 5176 4310 5228
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 4341 5179 4399 5185
rect 3510 5148 3516 5160
rect 3436 5120 3516 5148
rect 3510 5108 3516 5120
rect 3568 5108 3574 5160
rect 4065 5151 4123 5157
rect 4065 5117 4077 5151
rect 4111 5148 4123 5151
rect 4356 5148 4384 5179
rect 4111 5120 4384 5148
rect 4908 5148 4936 5324
rect 5169 5321 5181 5355
rect 5215 5352 5227 5355
rect 10870 5352 10876 5364
rect 5215 5324 10876 5352
rect 5215 5321 5227 5324
rect 5169 5315 5227 5321
rect 10870 5312 10876 5324
rect 10928 5312 10934 5364
rect 15378 5312 15384 5364
rect 15436 5352 15442 5364
rect 15436 5324 18092 5352
rect 15436 5312 15442 5324
rect 6178 5284 6184 5296
rect 5552 5256 6184 5284
rect 4982 5176 4988 5228
rect 5040 5216 5046 5228
rect 5552 5225 5580 5256
rect 6178 5244 6184 5256
rect 6236 5244 6242 5296
rect 13998 5284 14004 5296
rect 12406 5256 14004 5284
rect 5077 5219 5135 5225
rect 5077 5216 5089 5219
rect 5040 5188 5089 5216
rect 5040 5176 5046 5188
rect 5077 5185 5089 5188
rect 5123 5185 5135 5219
rect 5077 5179 5135 5185
rect 5537 5219 5595 5225
rect 5537 5185 5549 5219
rect 5583 5185 5595 5219
rect 5537 5179 5595 5185
rect 5350 5148 5356 5160
rect 4908 5120 5356 5148
rect 4111 5117 4123 5120
rect 4065 5111 4123 5117
rect 2869 5083 2927 5089
rect 2869 5049 2881 5083
rect 2915 5049 2927 5083
rect 2869 5043 2927 5049
rect 3418 5040 3424 5092
rect 3476 5080 3482 5092
rect 4080 5080 4108 5111
rect 3476 5052 4108 5080
rect 4356 5080 4384 5120
rect 5350 5108 5356 5120
rect 5408 5108 5414 5160
rect 12406 5080 12434 5256
rect 13998 5244 14004 5256
rect 14056 5244 14062 5296
rect 17681 5287 17739 5293
rect 17681 5253 17693 5287
rect 17727 5284 17739 5287
rect 17954 5284 17960 5296
rect 17727 5256 17960 5284
rect 17727 5253 17739 5256
rect 17681 5247 17739 5253
rect 17954 5244 17960 5256
rect 18012 5244 18018 5296
rect 18064 5284 18092 5324
rect 18414 5312 18420 5364
rect 18472 5352 18478 5364
rect 19153 5355 19211 5361
rect 19153 5352 19165 5355
rect 18472 5324 19165 5352
rect 18472 5312 18478 5324
rect 19153 5321 19165 5324
rect 19199 5321 19211 5355
rect 19153 5315 19211 5321
rect 21174 5312 21180 5364
rect 21232 5312 21238 5364
rect 21450 5312 21456 5364
rect 21508 5352 21514 5364
rect 21545 5355 21603 5361
rect 21545 5352 21557 5355
rect 21508 5324 21557 5352
rect 21508 5312 21514 5324
rect 21545 5321 21557 5324
rect 21591 5321 21603 5355
rect 21545 5315 21603 5321
rect 24394 5312 24400 5364
rect 24452 5352 24458 5364
rect 24452 5324 25084 5352
rect 24452 5312 24458 5324
rect 18064 5256 18170 5284
rect 20898 5244 20904 5296
rect 20956 5284 20962 5296
rect 21818 5284 21824 5296
rect 20956 5256 21824 5284
rect 20956 5244 20962 5256
rect 21818 5244 21824 5256
rect 21876 5284 21882 5296
rect 21876 5256 23598 5284
rect 21876 5244 21882 5256
rect 17310 5176 17316 5228
rect 17368 5216 17374 5228
rect 25056 5225 25084 5324
rect 17405 5219 17463 5225
rect 17405 5216 17417 5219
rect 17368 5188 17417 5216
rect 17368 5176 17374 5188
rect 17405 5185 17417 5188
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 25041 5219 25099 5225
rect 25041 5185 25053 5219
rect 25087 5185 25099 5219
rect 25041 5179 25099 5185
rect 20714 5108 20720 5160
rect 20772 5148 20778 5160
rect 20901 5151 20959 5157
rect 20901 5148 20913 5151
rect 20772 5120 20913 5148
rect 20772 5108 20778 5120
rect 20901 5117 20913 5120
rect 20947 5117 20959 5151
rect 20901 5111 20959 5117
rect 21085 5151 21143 5157
rect 21085 5117 21097 5151
rect 21131 5148 21143 5151
rect 21910 5148 21916 5160
rect 21131 5120 21916 5148
rect 21131 5117 21143 5120
rect 21085 5111 21143 5117
rect 21910 5108 21916 5120
rect 21968 5108 21974 5160
rect 24765 5151 24823 5157
rect 24765 5117 24777 5151
rect 24811 5148 24823 5151
rect 25130 5148 25136 5160
rect 24811 5120 25136 5148
rect 24811 5117 24823 5120
rect 24765 5111 24823 5117
rect 25130 5108 25136 5120
rect 25188 5108 25194 5160
rect 4356 5052 12434 5080
rect 3476 5040 3482 5052
rect 2501 5015 2559 5021
rect 2501 5012 2513 5015
rect 2240 4984 2513 5012
rect 2501 4981 2513 4984
rect 2547 4981 2559 5015
rect 2501 4975 2559 4981
rect 3050 4972 3056 5024
rect 3108 5012 3114 5024
rect 3602 5012 3608 5024
rect 3108 4984 3608 5012
rect 3108 4972 3114 4984
rect 3602 4972 3608 4984
rect 3660 4972 3666 5024
rect 4249 5015 4307 5021
rect 4249 4981 4261 5015
rect 4295 5012 4307 5015
rect 4525 5015 4583 5021
rect 4525 5012 4537 5015
rect 4295 4984 4537 5012
rect 4295 4981 4307 4984
rect 4249 4975 4307 4981
rect 4525 4981 4537 4984
rect 4571 5012 4583 5015
rect 4614 5012 4620 5024
rect 4571 4984 4620 5012
rect 4571 4981 4583 4984
rect 4525 4975 4583 4981
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 4706 4972 4712 5024
rect 4764 4972 4770 5024
rect 5718 4972 5724 5024
rect 5776 5012 5782 5024
rect 5997 5015 6055 5021
rect 5997 5012 6009 5015
rect 5776 4984 6009 5012
rect 5776 4972 5782 4984
rect 5997 4981 6009 4984
rect 6043 5012 6055 5015
rect 6822 5012 6828 5024
rect 6043 4984 6828 5012
rect 6043 4981 6055 4984
rect 5997 4975 6055 4981
rect 6822 4972 6828 4984
rect 6880 5012 6886 5024
rect 8294 5012 8300 5024
rect 6880 4984 8300 5012
rect 6880 4972 6886 4984
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 23290 4972 23296 5024
rect 23348 4972 23354 5024
rect 1104 4922 28888 4944
rect 1104 4870 2918 4922
rect 2970 4870 2982 4922
rect 3034 4870 3046 4922
rect 3098 4870 3110 4922
rect 3162 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 10918 4922
rect 10970 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 11238 4922
rect 11290 4870 18918 4922
rect 18970 4870 18982 4922
rect 19034 4870 19046 4922
rect 19098 4870 19110 4922
rect 19162 4870 19174 4922
rect 19226 4870 19238 4922
rect 19290 4870 26918 4922
rect 26970 4870 26982 4922
rect 27034 4870 27046 4922
rect 27098 4870 27110 4922
rect 27162 4870 27174 4922
rect 27226 4870 27238 4922
rect 27290 4870 28888 4922
rect 1104 4848 28888 4870
rect 2958 4768 2964 4820
rect 3016 4808 3022 4820
rect 3145 4811 3203 4817
rect 3145 4808 3157 4811
rect 3016 4780 3157 4808
rect 3016 4768 3022 4780
rect 3145 4777 3157 4780
rect 3191 4808 3203 4811
rect 4062 4808 4068 4820
rect 3191 4780 4068 4808
rect 3191 4777 3203 4780
rect 3145 4771 3203 4777
rect 4062 4768 4068 4780
rect 4120 4768 4126 4820
rect 4246 4768 4252 4820
rect 4304 4808 4310 4820
rect 4304 4780 7052 4808
rect 4304 4768 4310 4780
rect 3510 4700 3516 4752
rect 3568 4700 3574 4752
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 3326 4672 3332 4684
rect 1443 4644 3332 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 3326 4632 3332 4644
rect 3384 4672 3390 4684
rect 3789 4675 3847 4681
rect 3789 4672 3801 4675
rect 3384 4644 3801 4672
rect 3384 4632 3390 4644
rect 3789 4641 3801 4644
rect 3835 4641 3847 4675
rect 3789 4635 3847 4641
rect 4065 4675 4123 4681
rect 4065 4641 4077 4675
rect 4111 4672 4123 4675
rect 4706 4672 4712 4684
rect 4111 4644 4712 4672
rect 4111 4641 4123 4644
rect 4065 4635 4123 4641
rect 4706 4632 4712 4644
rect 4764 4632 4770 4684
rect 6914 4632 6920 4684
rect 6972 4632 6978 4684
rect 7024 4672 7052 4780
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 8665 4811 8723 4817
rect 8665 4808 8677 4811
rect 8260 4780 8677 4808
rect 8260 4768 8266 4780
rect 8665 4777 8677 4780
rect 8711 4777 8723 4811
rect 8665 4771 8723 4777
rect 12526 4768 12532 4820
rect 12584 4808 12590 4820
rect 18141 4811 18199 4817
rect 18141 4808 18153 4811
rect 12584 4780 18153 4808
rect 12584 4768 12590 4780
rect 18141 4777 18153 4780
rect 18187 4777 18199 4811
rect 18141 4771 18199 4777
rect 9674 4672 9680 4684
rect 7024 4644 9680 4672
rect 9674 4632 9680 4644
rect 9732 4672 9738 4684
rect 11514 4672 11520 4684
rect 9732 4644 11520 4672
rect 9732 4632 9738 4644
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 14826 4632 14832 4684
rect 14884 4672 14890 4684
rect 15197 4675 15255 4681
rect 15197 4672 15209 4675
rect 14884 4644 15209 4672
rect 14884 4632 14890 4644
rect 15197 4641 15209 4644
rect 15243 4641 15255 4675
rect 15197 4635 15255 4641
rect 2774 4564 2780 4616
rect 2832 4564 2838 4616
rect 3237 4607 3295 4613
rect 3237 4573 3249 4607
rect 3283 4604 3295 4607
rect 3602 4604 3608 4616
rect 3283 4576 3608 4604
rect 3283 4573 3295 4576
rect 3237 4567 3295 4573
rect 3602 4564 3608 4576
rect 3660 4564 3666 4616
rect 14737 4607 14795 4613
rect 14737 4573 14749 4607
rect 14783 4604 14795 4607
rect 16022 4604 16028 4616
rect 14783 4576 16028 4604
rect 14783 4573 14795 4576
rect 14737 4567 14795 4573
rect 16022 4564 16028 4576
rect 16080 4564 16086 4616
rect 18156 4604 18184 4771
rect 18506 4768 18512 4820
rect 18564 4768 18570 4820
rect 21910 4768 21916 4820
rect 21968 4768 21974 4820
rect 25130 4768 25136 4820
rect 25188 4768 25194 4820
rect 22002 4700 22008 4752
rect 22060 4740 22066 4752
rect 22060 4712 24532 4740
rect 22060 4700 22066 4712
rect 18506 4632 18512 4684
rect 18564 4672 18570 4684
rect 22557 4675 22615 4681
rect 22557 4672 22569 4675
rect 18564 4644 22569 4672
rect 18564 4632 18570 4644
rect 22557 4641 22569 4644
rect 22603 4672 22615 4675
rect 24210 4672 24216 4684
rect 22603 4644 24216 4672
rect 22603 4641 22615 4644
rect 22557 4635 22615 4641
rect 24210 4632 24216 4644
rect 24268 4632 24274 4684
rect 24504 4681 24532 4712
rect 24489 4675 24547 4681
rect 24489 4641 24501 4675
rect 24535 4641 24547 4675
rect 24489 4635 24547 4641
rect 24670 4632 24676 4684
rect 24728 4632 24734 4684
rect 18325 4607 18383 4613
rect 18325 4604 18337 4607
rect 18156 4576 18337 4604
rect 18325 4573 18337 4576
rect 18371 4573 18383 4607
rect 18325 4567 18383 4573
rect 22281 4607 22339 4613
rect 22281 4573 22293 4607
rect 22327 4604 22339 4607
rect 23290 4604 23296 4616
rect 22327 4576 23296 4604
rect 22327 4573 22339 4576
rect 22281 4567 22339 4573
rect 23290 4564 23296 4576
rect 23348 4604 23354 4616
rect 24765 4607 24823 4613
rect 24765 4604 24777 4607
rect 23348 4576 24777 4604
rect 23348 4564 23354 4576
rect 24765 4573 24777 4576
rect 24811 4573 24823 4607
rect 24765 4567 24823 4573
rect 1670 4496 1676 4548
rect 1728 4496 1734 4548
rect 2792 4468 2820 4564
rect 5290 4508 5672 4536
rect 5368 4468 5396 4508
rect 5644 4480 5672 4508
rect 7190 4496 7196 4548
rect 7248 4496 7254 4548
rect 7300 4508 7682 4536
rect 2792 4440 5396 4468
rect 5442 4428 5448 4480
rect 5500 4468 5506 4480
rect 5537 4471 5595 4477
rect 5537 4468 5549 4471
rect 5500 4440 5549 4468
rect 5500 4428 5506 4440
rect 5537 4437 5549 4440
rect 5583 4437 5595 4471
rect 5537 4431 5595 4437
rect 5626 4428 5632 4480
rect 5684 4468 5690 4480
rect 7300 4468 7328 4508
rect 13906 4496 13912 4548
rect 13964 4536 13970 4548
rect 15381 4539 15439 4545
rect 13964 4508 14872 4536
rect 13964 4496 13970 4508
rect 5684 4440 7328 4468
rect 14277 4471 14335 4477
rect 5684 4428 5690 4440
rect 14277 4437 14289 4471
rect 14323 4468 14335 4471
rect 14366 4468 14372 4480
rect 14323 4440 14372 4468
rect 14323 4437 14335 4440
rect 14277 4431 14335 4437
rect 14366 4428 14372 4440
rect 14424 4428 14430 4480
rect 14645 4471 14703 4477
rect 14645 4437 14657 4471
rect 14691 4468 14703 4471
rect 14734 4468 14740 4480
rect 14691 4440 14740 4468
rect 14691 4437 14703 4440
rect 14645 4431 14703 4437
rect 14734 4428 14740 4440
rect 14792 4428 14798 4480
rect 14844 4468 14872 4508
rect 15381 4505 15393 4539
rect 15427 4536 15439 4539
rect 17862 4536 17868 4548
rect 15427 4508 17868 4536
rect 15427 4505 15439 4508
rect 15381 4499 15439 4505
rect 17862 4496 17868 4508
rect 17920 4496 17926 4548
rect 15473 4471 15531 4477
rect 15473 4468 15485 4471
rect 14844 4440 15485 4468
rect 15473 4437 15485 4440
rect 15519 4437 15531 4471
rect 15473 4431 15531 4437
rect 15654 4428 15660 4480
rect 15712 4468 15718 4480
rect 15841 4471 15899 4477
rect 15841 4468 15853 4471
rect 15712 4440 15853 4468
rect 15712 4428 15718 4440
rect 15841 4437 15853 4440
rect 15887 4437 15899 4471
rect 15841 4431 15899 4437
rect 22370 4428 22376 4480
rect 22428 4428 22434 4480
rect 1104 4378 28888 4400
rect 1104 4326 3658 4378
rect 3710 4326 3722 4378
rect 3774 4326 3786 4378
rect 3838 4326 3850 4378
rect 3902 4326 3914 4378
rect 3966 4326 3978 4378
rect 4030 4326 11658 4378
rect 11710 4326 11722 4378
rect 11774 4326 11786 4378
rect 11838 4326 11850 4378
rect 11902 4326 11914 4378
rect 11966 4326 11978 4378
rect 12030 4326 19658 4378
rect 19710 4326 19722 4378
rect 19774 4326 19786 4378
rect 19838 4326 19850 4378
rect 19902 4326 19914 4378
rect 19966 4326 19978 4378
rect 20030 4326 27658 4378
rect 27710 4326 27722 4378
rect 27774 4326 27786 4378
rect 27838 4326 27850 4378
rect 27902 4326 27914 4378
rect 27966 4326 27978 4378
rect 28030 4326 28888 4378
rect 1104 4304 28888 4326
rect 1670 4224 1676 4276
rect 1728 4264 1734 4276
rect 2593 4267 2651 4273
rect 2593 4264 2605 4267
rect 1728 4236 2605 4264
rect 1728 4224 1734 4236
rect 2593 4233 2605 4236
rect 2639 4233 2651 4267
rect 2593 4227 2651 4233
rect 2958 4224 2964 4276
rect 3016 4224 3022 4276
rect 4617 4267 4675 4273
rect 4617 4233 4629 4267
rect 4663 4264 4675 4267
rect 4982 4264 4988 4276
rect 4663 4236 4988 4264
rect 4663 4233 4675 4236
rect 4617 4227 4675 4233
rect 4982 4224 4988 4236
rect 5040 4264 5046 4276
rect 5442 4264 5448 4276
rect 5040 4236 5448 4264
rect 5040 4224 5046 4236
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 7190 4224 7196 4276
rect 7248 4264 7254 4276
rect 7469 4267 7527 4273
rect 7469 4264 7481 4267
rect 7248 4236 7481 4264
rect 7248 4224 7254 4236
rect 7469 4233 7481 4236
rect 7515 4233 7527 4267
rect 7469 4227 7527 4233
rect 7837 4267 7895 4273
rect 7837 4233 7849 4267
rect 7883 4264 7895 4267
rect 8202 4264 8208 4276
rect 7883 4236 8208 4264
rect 7883 4233 7895 4236
rect 7837 4227 7895 4233
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 17862 4224 17868 4276
rect 17920 4224 17926 4276
rect 18325 4267 18383 4273
rect 18325 4233 18337 4267
rect 18371 4264 18383 4267
rect 18414 4264 18420 4276
rect 18371 4236 18420 4264
rect 18371 4233 18383 4236
rect 18325 4227 18383 4233
rect 18414 4224 18420 4236
rect 18472 4264 18478 4276
rect 19153 4267 19211 4273
rect 19153 4264 19165 4267
rect 18472 4236 19165 4264
rect 18472 4224 18478 4236
rect 19153 4233 19165 4236
rect 19199 4233 19211 4267
rect 19153 4227 19211 4233
rect 22189 4267 22247 4273
rect 22189 4233 22201 4267
rect 22235 4264 22247 4267
rect 22370 4264 22376 4276
rect 22235 4236 22376 4264
rect 22235 4233 22247 4236
rect 22189 4227 22247 4233
rect 22370 4224 22376 4236
rect 22428 4224 22434 4276
rect 23017 4267 23075 4273
rect 23017 4233 23029 4267
rect 23063 4264 23075 4267
rect 23290 4264 23296 4276
rect 23063 4236 23296 4264
rect 23063 4233 23075 4236
rect 23017 4227 23075 4233
rect 23290 4224 23296 4236
rect 23348 4224 23354 4276
rect 4525 4199 4583 4205
rect 4525 4165 4537 4199
rect 4571 4196 4583 4199
rect 5166 4196 5172 4208
rect 4571 4168 5172 4196
rect 4571 4165 4583 4168
rect 4525 4159 4583 4165
rect 5166 4156 5172 4168
rect 5224 4156 5230 4208
rect 8665 4199 8723 4205
rect 8665 4165 8677 4199
rect 8711 4196 8723 4199
rect 9306 4196 9312 4208
rect 8711 4168 9312 4196
rect 8711 4165 8723 4168
rect 8665 4159 8723 4165
rect 9306 4156 9312 4168
rect 9364 4196 9370 4208
rect 10873 4199 10931 4205
rect 10873 4196 10885 4199
rect 9364 4168 10885 4196
rect 9364 4156 9370 4168
rect 10873 4165 10885 4168
rect 10919 4165 10931 4199
rect 10873 4159 10931 4165
rect 11330 4156 11336 4208
rect 11388 4196 11394 4208
rect 11790 4196 11796 4208
rect 11388 4168 11796 4196
rect 11388 4156 11394 4168
rect 11790 4156 11796 4168
rect 11848 4196 11854 4208
rect 11885 4199 11943 4205
rect 11885 4196 11897 4199
rect 11848 4168 11897 4196
rect 11848 4156 11854 4168
rect 11885 4165 11897 4168
rect 11931 4165 11943 4199
rect 11885 4159 11943 4165
rect 11977 4199 12035 4205
rect 11977 4165 11989 4199
rect 12023 4196 12035 4199
rect 12158 4196 12164 4208
rect 12023 4168 12164 4196
rect 12023 4165 12035 4168
rect 11977 4159 12035 4165
rect 12158 4156 12164 4168
rect 12216 4156 12222 4208
rect 15378 4196 15384 4208
rect 15226 4168 15384 4196
rect 15378 4156 15384 4168
rect 15436 4156 15442 4208
rect 15654 4156 15660 4208
rect 15712 4156 15718 4208
rect 18233 4199 18291 4205
rect 18233 4165 18245 4199
rect 18279 4196 18291 4199
rect 19061 4199 19119 4205
rect 19061 4196 19073 4199
rect 18279 4168 19073 4196
rect 18279 4165 18291 4168
rect 18233 4159 18291 4165
rect 19061 4165 19073 4168
rect 19107 4196 19119 4199
rect 20438 4196 20444 4208
rect 19107 4168 20444 4196
rect 19107 4165 19119 4168
rect 19061 4159 19119 4165
rect 20438 4156 20444 4168
rect 20496 4156 20502 4208
rect 22388 4196 22416 4224
rect 22830 4196 22836 4208
rect 22388 4168 22836 4196
rect 22830 4156 22836 4168
rect 22888 4196 22894 4208
rect 23109 4199 23167 4205
rect 23109 4196 23121 4199
rect 22888 4168 23121 4196
rect 22888 4156 22894 4168
rect 23109 4165 23121 4168
rect 23155 4165 23167 4199
rect 23109 4159 23167 4165
rect 4614 4088 4620 4140
rect 4672 4128 4678 4140
rect 5077 4131 5135 4137
rect 5077 4128 5089 4131
rect 4672 4100 5089 4128
rect 4672 4088 4678 4100
rect 4816 4069 4844 4100
rect 5077 4097 5089 4100
rect 5123 4128 5135 4131
rect 12437 4131 12495 4137
rect 5123 4100 12388 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 8956 4072 8984 4100
rect 3053 4063 3111 4069
rect 3053 4029 3065 4063
rect 3099 4029 3111 4063
rect 3053 4023 3111 4029
rect 3237 4063 3295 4069
rect 3237 4029 3249 4063
rect 3283 4060 3295 4063
rect 4801 4063 4859 4069
rect 3283 4032 4752 4060
rect 3283 4029 3295 4032
rect 3237 4023 3295 4029
rect 3068 3992 3096 4023
rect 4157 3995 4215 4001
rect 4157 3992 4169 3995
rect 3068 3964 4169 3992
rect 4157 3961 4169 3964
rect 4203 3961 4215 3995
rect 4724 3992 4752 4032
rect 4801 4029 4813 4063
rect 4847 4029 4859 4063
rect 4801 4023 4859 4029
rect 7929 4063 7987 4069
rect 7929 4029 7941 4063
rect 7975 4029 7987 4063
rect 7929 4023 7987 4029
rect 5350 3992 5356 4004
rect 4724 3964 5356 3992
rect 4157 3955 4215 3961
rect 5350 3952 5356 3964
rect 5408 3952 5414 4004
rect 7944 3992 7972 4023
rect 8110 4020 8116 4072
rect 8168 4020 8174 4072
rect 8754 4020 8760 4072
rect 8812 4020 8818 4072
rect 8938 4020 8944 4072
rect 8996 4020 9002 4072
rect 10689 4063 10747 4069
rect 10689 4029 10701 4063
rect 10735 4029 10747 4063
rect 10689 4023 10747 4029
rect 8297 3995 8355 4001
rect 8297 3992 8309 3995
rect 7944 3964 8309 3992
rect 8297 3961 8309 3964
rect 8343 3961 8355 3995
rect 10704 3992 10732 4023
rect 10778 4020 10784 4072
rect 10836 4020 10842 4072
rect 12066 4020 12072 4072
rect 12124 4020 12130 4072
rect 12084 3992 12112 4020
rect 10704 3964 12112 3992
rect 8297 3955 8355 3961
rect 11241 3927 11299 3933
rect 11241 3893 11253 3927
rect 11287 3924 11299 3927
rect 11422 3924 11428 3936
rect 11287 3896 11428 3924
rect 11287 3893 11299 3896
rect 11241 3887 11299 3893
rect 11422 3884 11428 3896
rect 11480 3884 11486 3936
rect 11517 3927 11575 3933
rect 11517 3893 11529 3927
rect 11563 3924 11575 3927
rect 11882 3924 11888 3936
rect 11563 3896 11888 3924
rect 11563 3893 11575 3896
rect 11517 3887 11575 3893
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 12360 3924 12388 4100
rect 12437 4097 12449 4131
rect 12483 4128 12495 4131
rect 12526 4128 12532 4140
rect 12483 4100 12532 4128
rect 12483 4097 12495 4100
rect 12437 4091 12495 4097
rect 12452 3924 12480 4091
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 15933 4131 15991 4137
rect 15933 4097 15945 4131
rect 15979 4128 15991 4131
rect 17310 4128 17316 4140
rect 15979 4100 17316 4128
rect 15979 4097 15991 4100
rect 15933 4091 15991 4097
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 22278 4088 22284 4140
rect 22336 4088 22342 4140
rect 13906 4020 13912 4072
rect 13964 4060 13970 4072
rect 14185 4063 14243 4069
rect 14185 4060 14197 4063
rect 13964 4032 14197 4060
rect 13964 4020 13970 4032
rect 14185 4029 14197 4032
rect 14231 4029 14243 4063
rect 14185 4023 14243 4029
rect 18506 4020 18512 4072
rect 18564 4020 18570 4072
rect 19245 4063 19303 4069
rect 19245 4029 19257 4063
rect 19291 4029 19303 4063
rect 19245 4023 19303 4029
rect 18598 3952 18604 4004
rect 18656 3992 18662 4004
rect 19260 3992 19288 4023
rect 20714 4020 20720 4072
rect 20772 4060 20778 4072
rect 22002 4060 22008 4072
rect 20772 4032 22008 4060
rect 20772 4020 20778 4032
rect 22002 4020 22008 4032
rect 22060 4060 22066 4072
rect 22373 4063 22431 4069
rect 22373 4060 22385 4063
rect 22060 4032 22385 4060
rect 22060 4020 22066 4032
rect 22373 4029 22385 4032
rect 22419 4029 22431 4063
rect 22373 4023 22431 4029
rect 23293 4063 23351 4069
rect 23293 4029 23305 4063
rect 23339 4060 23351 4063
rect 24762 4060 24768 4072
rect 23339 4032 24768 4060
rect 23339 4029 23351 4032
rect 23293 4023 23351 4029
rect 23308 3992 23336 4023
rect 24762 4020 24768 4032
rect 24820 4020 24826 4072
rect 18656 3964 23336 3992
rect 18656 3952 18662 3964
rect 12802 3924 12808 3936
rect 12360 3896 12808 3924
rect 12802 3884 12808 3896
rect 12860 3884 12866 3936
rect 17402 3884 17408 3936
rect 17460 3924 17466 3936
rect 18693 3927 18751 3933
rect 18693 3924 18705 3927
rect 17460 3896 18705 3924
rect 17460 3884 17466 3896
rect 18693 3893 18705 3896
rect 18739 3893 18751 3927
rect 18693 3887 18751 3893
rect 21450 3884 21456 3936
rect 21508 3924 21514 3936
rect 21821 3927 21879 3933
rect 21821 3924 21833 3927
rect 21508 3896 21833 3924
rect 21508 3884 21514 3896
rect 21821 3893 21833 3896
rect 21867 3893 21879 3927
rect 21821 3887 21879 3893
rect 22646 3884 22652 3936
rect 22704 3884 22710 3936
rect 1104 3834 28888 3856
rect 1104 3782 2918 3834
rect 2970 3782 2982 3834
rect 3034 3782 3046 3834
rect 3098 3782 3110 3834
rect 3162 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 10918 3834
rect 10970 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 11238 3834
rect 11290 3782 18918 3834
rect 18970 3782 18982 3834
rect 19034 3782 19046 3834
rect 19098 3782 19110 3834
rect 19162 3782 19174 3834
rect 19226 3782 19238 3834
rect 19290 3782 26918 3834
rect 26970 3782 26982 3834
rect 27034 3782 27046 3834
rect 27098 3782 27110 3834
rect 27162 3782 27174 3834
rect 27226 3782 27238 3834
rect 27290 3782 28888 3834
rect 1104 3760 28888 3782
rect 5166 3680 5172 3732
rect 5224 3720 5230 3732
rect 5537 3723 5595 3729
rect 5537 3720 5549 3723
rect 5224 3692 5549 3720
rect 5224 3680 5230 3692
rect 5537 3689 5549 3692
rect 5583 3689 5595 3723
rect 5537 3683 5595 3689
rect 8481 3723 8539 3729
rect 8481 3689 8493 3723
rect 8527 3720 8539 3723
rect 8938 3720 8944 3732
rect 8527 3692 8944 3720
rect 8527 3689 8539 3692
rect 8481 3683 8539 3689
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 10413 3723 10471 3729
rect 10413 3689 10425 3723
rect 10459 3720 10471 3723
rect 11790 3720 11796 3732
rect 10459 3692 11796 3720
rect 10459 3689 10471 3692
rect 10413 3683 10471 3689
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 12158 3680 12164 3732
rect 12216 3720 12222 3732
rect 12253 3723 12311 3729
rect 12253 3720 12265 3723
rect 12216 3692 12265 3720
rect 12216 3680 12222 3692
rect 12253 3689 12265 3692
rect 12299 3689 12311 3723
rect 14734 3720 14740 3732
rect 12253 3683 12311 3689
rect 12728 3692 14740 3720
rect 12728 3596 12756 3692
rect 14734 3680 14740 3692
rect 14792 3720 14798 3732
rect 15841 3723 15899 3729
rect 15841 3720 15853 3723
rect 14792 3692 15853 3720
rect 14792 3680 14798 3692
rect 15841 3689 15853 3692
rect 15887 3689 15899 3723
rect 15841 3683 15899 3689
rect 18598 3680 18604 3732
rect 18656 3680 18662 3732
rect 22830 3680 22836 3732
rect 22888 3680 22894 3732
rect 3326 3544 3332 3596
rect 3384 3584 3390 3596
rect 3789 3587 3847 3593
rect 3789 3584 3801 3587
rect 3384 3556 3801 3584
rect 3384 3544 3390 3556
rect 3789 3553 3801 3556
rect 3835 3553 3847 3587
rect 3789 3547 3847 3553
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3584 6607 3587
rect 6822 3584 6828 3596
rect 6595 3556 6828 3584
rect 6595 3553 6607 3556
rect 6549 3547 6607 3553
rect 6822 3544 6828 3556
rect 6880 3544 6886 3596
rect 8294 3544 8300 3596
rect 8352 3584 8358 3596
rect 8757 3587 8815 3593
rect 8757 3584 8769 3587
rect 8352 3556 8769 3584
rect 8352 3544 8358 3556
rect 8757 3553 8769 3556
rect 8803 3584 8815 3587
rect 9585 3587 9643 3593
rect 9585 3584 9597 3587
rect 8803 3556 9597 3584
rect 8803 3553 8815 3556
rect 8757 3547 8815 3553
rect 9585 3553 9597 3556
rect 9631 3584 9643 3587
rect 11514 3584 11520 3596
rect 9631 3556 11520 3584
rect 9631 3553 9643 3556
rect 9585 3547 9643 3553
rect 11514 3544 11520 3556
rect 11572 3544 11578 3596
rect 11882 3544 11888 3596
rect 11940 3544 11946 3596
rect 12710 3544 12716 3596
rect 12768 3544 12774 3596
rect 12802 3544 12808 3596
rect 12860 3544 12866 3596
rect 13814 3544 13820 3596
rect 13872 3584 13878 3596
rect 14093 3587 14151 3593
rect 14093 3584 14105 3587
rect 13872 3556 14105 3584
rect 13872 3544 13878 3556
rect 14093 3553 14105 3556
rect 14139 3553 14151 3587
rect 14093 3547 14151 3553
rect 14366 3544 14372 3596
rect 14424 3544 14430 3596
rect 17310 3544 17316 3596
rect 17368 3584 17374 3596
rect 18049 3587 18107 3593
rect 18049 3584 18061 3587
rect 17368 3556 18061 3584
rect 17368 3544 17374 3556
rect 18049 3553 18061 3556
rect 18095 3584 18107 3587
rect 19245 3587 19303 3593
rect 19245 3584 19257 3587
rect 18095 3556 19257 3584
rect 18095 3553 18107 3556
rect 18049 3547 18107 3553
rect 19245 3553 19257 3556
rect 19291 3553 19303 3587
rect 19245 3547 19303 3553
rect 21085 3587 21143 3593
rect 21085 3553 21097 3587
rect 21131 3584 21143 3587
rect 21358 3584 21364 3596
rect 21131 3556 21364 3584
rect 21131 3553 21143 3556
rect 21085 3547 21143 3553
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 9306 3476 9312 3528
rect 9364 3476 9370 3528
rect 12158 3476 12164 3528
rect 12216 3516 12222 3528
rect 13832 3516 13860 3544
rect 12216 3488 13860 3516
rect 12216 3476 12222 3488
rect 15470 3476 15476 3528
rect 15528 3516 15534 3528
rect 18417 3519 18475 3525
rect 18417 3516 18429 3519
rect 15528 3488 16698 3516
rect 18248 3488 18429 3516
rect 15528 3476 15534 3488
rect 4062 3408 4068 3460
rect 4120 3408 4126 3460
rect 5626 3448 5632 3460
rect 5290 3420 5632 3448
rect 5626 3408 5632 3420
rect 5684 3408 5690 3460
rect 6822 3408 6828 3460
rect 6880 3408 6886 3460
rect 7282 3408 7288 3460
rect 7340 3408 7346 3460
rect 8754 3448 8760 3460
rect 8312 3420 8760 3448
rect 8312 3392 8340 3420
rect 8754 3408 8760 3420
rect 8812 3448 8818 3460
rect 9401 3451 9459 3457
rect 9401 3448 9413 3451
rect 8812 3420 9413 3448
rect 8812 3408 8818 3420
rect 9401 3417 9413 3420
rect 9447 3417 9459 3451
rect 9401 3411 9459 3417
rect 9674 3408 9680 3460
rect 9732 3448 9738 3460
rect 17773 3451 17831 3457
rect 9732 3420 10718 3448
rect 9732 3408 9738 3420
rect 17773 3417 17785 3451
rect 17819 3448 17831 3451
rect 17862 3448 17868 3460
rect 17819 3420 17868 3448
rect 17819 3417 17831 3420
rect 17773 3411 17831 3417
rect 17862 3408 17868 3420
rect 17920 3408 17926 3460
rect 8294 3340 8300 3392
rect 8352 3340 8358 3392
rect 8938 3340 8944 3392
rect 8996 3340 9002 3392
rect 12618 3340 12624 3392
rect 12676 3340 12682 3392
rect 16298 3340 16304 3392
rect 16356 3340 16362 3392
rect 17126 3340 17132 3392
rect 17184 3380 17190 3392
rect 18248 3389 18276 3488
rect 18417 3485 18429 3488
rect 18463 3485 18475 3519
rect 18417 3479 18475 3485
rect 19518 3408 19524 3460
rect 19576 3408 19582 3460
rect 21361 3451 21419 3457
rect 20746 3420 21220 3448
rect 18233 3383 18291 3389
rect 18233 3380 18245 3383
rect 17184 3352 18245 3380
rect 17184 3340 17190 3352
rect 18233 3349 18245 3352
rect 18279 3349 18291 3383
rect 18233 3343 18291 3349
rect 20438 3340 20444 3392
rect 20496 3380 20502 3392
rect 20993 3383 21051 3389
rect 20993 3380 21005 3383
rect 20496 3352 21005 3380
rect 20496 3340 20502 3352
rect 20993 3349 21005 3352
rect 21039 3349 21051 3383
rect 21192 3380 21220 3420
rect 21361 3417 21373 3451
rect 21407 3448 21419 3451
rect 21450 3448 21456 3460
rect 21407 3420 21456 3448
rect 21407 3417 21419 3420
rect 21361 3411 21419 3417
rect 21450 3408 21456 3420
rect 21508 3408 21514 3460
rect 21818 3448 21824 3460
rect 21560 3420 21824 3448
rect 21560 3380 21588 3420
rect 21818 3408 21824 3420
rect 21876 3408 21882 3460
rect 21192 3352 21588 3380
rect 20993 3343 21051 3349
rect 1104 3290 28888 3312
rect 1104 3238 3658 3290
rect 3710 3238 3722 3290
rect 3774 3238 3786 3290
rect 3838 3238 3850 3290
rect 3902 3238 3914 3290
rect 3966 3238 3978 3290
rect 4030 3238 11658 3290
rect 11710 3238 11722 3290
rect 11774 3238 11786 3290
rect 11838 3238 11850 3290
rect 11902 3238 11914 3290
rect 11966 3238 11978 3290
rect 12030 3238 19658 3290
rect 19710 3238 19722 3290
rect 19774 3238 19786 3290
rect 19838 3238 19850 3290
rect 19902 3238 19914 3290
rect 19966 3238 19978 3290
rect 20030 3238 27658 3290
rect 27710 3238 27722 3290
rect 27774 3238 27786 3290
rect 27838 3238 27850 3290
rect 27902 3238 27914 3290
rect 27966 3238 27978 3290
rect 28030 3238 28888 3290
rect 1104 3216 28888 3238
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 4433 3179 4491 3185
rect 4433 3176 4445 3179
rect 4120 3148 4445 3176
rect 4120 3136 4126 3148
rect 4433 3145 4445 3148
rect 4479 3145 4491 3179
rect 4433 3139 4491 3145
rect 4801 3179 4859 3185
rect 4801 3145 4813 3179
rect 4847 3176 4859 3179
rect 5166 3176 5172 3188
rect 4847 3148 5172 3176
rect 4847 3145 4859 3148
rect 4801 3139 4859 3145
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 6822 3136 6828 3188
rect 6880 3176 6886 3188
rect 7561 3179 7619 3185
rect 7561 3176 7573 3179
rect 6880 3148 7573 3176
rect 6880 3136 6886 3148
rect 7561 3145 7573 3148
rect 7607 3145 7619 3179
rect 7561 3139 7619 3145
rect 7929 3179 7987 3185
rect 7929 3145 7941 3179
rect 7975 3176 7987 3179
rect 8294 3176 8300 3188
rect 7975 3148 8300 3176
rect 7975 3145 7987 3148
rect 7929 3139 7987 3145
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 9306 3136 9312 3188
rect 9364 3176 9370 3188
rect 9493 3179 9551 3185
rect 9493 3176 9505 3179
rect 9364 3148 9505 3176
rect 9364 3136 9370 3148
rect 9493 3145 9505 3148
rect 9539 3145 9551 3179
rect 9493 3139 9551 3145
rect 10778 3136 10784 3188
rect 10836 3176 10842 3188
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 10836 3148 12173 3176
rect 10836 3136 10842 3148
rect 12161 3145 12173 3148
rect 12207 3145 12219 3179
rect 12161 3139 12219 3145
rect 12529 3179 12587 3185
rect 12529 3145 12541 3179
rect 12575 3176 12587 3179
rect 12618 3176 12624 3188
rect 12575 3148 12624 3176
rect 12575 3145 12587 3148
rect 12529 3139 12587 3145
rect 12618 3136 12624 3148
rect 12676 3176 12682 3188
rect 16298 3176 16304 3188
rect 12676 3148 16304 3176
rect 12676 3136 12682 3148
rect 16298 3136 16304 3148
rect 16356 3176 16362 3188
rect 17497 3179 17555 3185
rect 17497 3176 17509 3179
rect 16356 3148 17509 3176
rect 16356 3136 16362 3148
rect 17497 3145 17509 3148
rect 17543 3145 17555 3179
rect 17497 3139 17555 3145
rect 17862 3136 17868 3188
rect 17920 3136 17926 3188
rect 19518 3136 19524 3188
rect 19576 3176 19582 3188
rect 20073 3179 20131 3185
rect 20073 3176 20085 3179
rect 19576 3148 20085 3176
rect 19576 3136 19582 3148
rect 20073 3145 20085 3148
rect 20119 3145 20131 3179
rect 20073 3139 20131 3145
rect 20438 3136 20444 3188
rect 20496 3136 20502 3188
rect 20533 3179 20591 3185
rect 20533 3145 20545 3179
rect 20579 3176 20591 3179
rect 22646 3176 22652 3188
rect 20579 3148 22652 3176
rect 20579 3145 20591 3148
rect 20533 3139 20591 3145
rect 22646 3136 22652 3148
rect 22704 3136 22710 3188
rect 4893 3111 4951 3117
rect 4893 3077 4905 3111
rect 4939 3108 4951 3111
rect 8938 3108 8944 3120
rect 4939 3080 8944 3108
rect 4939 3077 4951 3080
rect 4893 3071 4951 3077
rect 8938 3068 8944 3080
rect 8996 3068 9002 3120
rect 9674 3068 9680 3120
rect 9732 3108 9738 3120
rect 10965 3111 11023 3117
rect 9732 3080 9798 3108
rect 9732 3068 9738 3080
rect 10965 3077 10977 3111
rect 11011 3108 11023 3111
rect 11422 3108 11428 3120
rect 11011 3080 11428 3108
rect 11011 3077 11023 3080
rect 10965 3071 11023 3077
rect 11422 3068 11428 3080
rect 11480 3068 11486 3120
rect 12710 3108 12716 3120
rect 12636 3080 12716 3108
rect 8021 3043 8079 3049
rect 8021 3009 8033 3043
rect 8067 3040 8079 3043
rect 11241 3043 11299 3049
rect 8067 3012 9812 3040
rect 8067 3009 8079 3012
rect 8021 3003 8079 3009
rect 5077 2975 5135 2981
rect 5077 2941 5089 2975
rect 5123 2972 5135 2975
rect 5350 2972 5356 2984
rect 5123 2944 5356 2972
rect 5123 2941 5135 2944
rect 5077 2935 5135 2941
rect 5350 2932 5356 2944
rect 5408 2972 5414 2984
rect 8110 2972 8116 2984
rect 5408 2944 8116 2972
rect 5408 2932 5414 2944
rect 8110 2932 8116 2944
rect 8168 2932 8174 2984
rect 9784 2972 9812 3012
rect 11241 3009 11253 3043
rect 11287 3040 11299 3043
rect 12158 3040 12164 3052
rect 11287 3012 12164 3040
rect 11287 3009 11299 3012
rect 11241 3003 11299 3009
rect 12158 3000 12164 3012
rect 12216 3000 12222 3052
rect 12636 3049 12664 3080
rect 12710 3068 12716 3080
rect 12768 3068 12774 3120
rect 17402 3068 17408 3120
rect 17460 3068 17466 3120
rect 12621 3043 12679 3049
rect 12621 3009 12633 3043
rect 12667 3009 12679 3043
rect 12621 3003 12679 3009
rect 9784 2944 11192 2972
rect 11164 2904 11192 2944
rect 11514 2932 11520 2984
rect 11572 2972 11578 2984
rect 12069 2975 12127 2981
rect 12069 2972 12081 2975
rect 11572 2944 12081 2972
rect 11572 2932 11578 2944
rect 12069 2941 12081 2944
rect 12115 2972 12127 2975
rect 12713 2975 12771 2981
rect 12713 2972 12725 2975
rect 12115 2944 12725 2972
rect 12115 2941 12127 2944
rect 12069 2935 12127 2941
rect 12713 2941 12725 2944
rect 12759 2972 12771 2975
rect 17126 2972 17132 2984
rect 12759 2944 17132 2972
rect 12759 2941 12771 2944
rect 12713 2935 12771 2941
rect 17126 2932 17132 2944
rect 17184 2932 17190 2984
rect 17218 2932 17224 2984
rect 17276 2932 17282 2984
rect 20714 2932 20720 2984
rect 20772 2932 20778 2984
rect 14090 2904 14096 2916
rect 11164 2876 14096 2904
rect 14090 2864 14096 2876
rect 14148 2864 14154 2916
rect 1104 2746 28888 2768
rect 1104 2694 2918 2746
rect 2970 2694 2982 2746
rect 3034 2694 3046 2746
rect 3098 2694 3110 2746
rect 3162 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 10918 2746
rect 10970 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 11238 2746
rect 11290 2694 18918 2746
rect 18970 2694 18982 2746
rect 19034 2694 19046 2746
rect 19098 2694 19110 2746
rect 19162 2694 19174 2746
rect 19226 2694 19238 2746
rect 19290 2694 26918 2746
rect 26970 2694 26982 2746
rect 27034 2694 27046 2746
rect 27098 2694 27110 2746
rect 27162 2694 27174 2746
rect 27226 2694 27238 2746
rect 27290 2694 28888 2746
rect 1104 2672 28888 2694
rect 1104 2202 28888 2224
rect 1104 2150 3658 2202
rect 3710 2150 3722 2202
rect 3774 2150 3786 2202
rect 3838 2150 3850 2202
rect 3902 2150 3914 2202
rect 3966 2150 3978 2202
rect 4030 2150 11658 2202
rect 11710 2150 11722 2202
rect 11774 2150 11786 2202
rect 11838 2150 11850 2202
rect 11902 2150 11914 2202
rect 11966 2150 11978 2202
rect 12030 2150 19658 2202
rect 19710 2150 19722 2202
rect 19774 2150 19786 2202
rect 19838 2150 19850 2202
rect 19902 2150 19914 2202
rect 19966 2150 19978 2202
rect 20030 2150 27658 2202
rect 27710 2150 27722 2202
rect 27774 2150 27786 2202
rect 27838 2150 27850 2202
rect 27902 2150 27914 2202
rect 27966 2150 27978 2202
rect 28030 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 2918 27718 2970 27770
rect 2982 27718 3034 27770
rect 3046 27718 3098 27770
rect 3110 27718 3162 27770
rect 3174 27718 3226 27770
rect 3238 27718 3290 27770
rect 10918 27718 10970 27770
rect 10982 27718 11034 27770
rect 11046 27718 11098 27770
rect 11110 27718 11162 27770
rect 11174 27718 11226 27770
rect 11238 27718 11290 27770
rect 18918 27718 18970 27770
rect 18982 27718 19034 27770
rect 19046 27718 19098 27770
rect 19110 27718 19162 27770
rect 19174 27718 19226 27770
rect 19238 27718 19290 27770
rect 26918 27718 26970 27770
rect 26982 27718 27034 27770
rect 27046 27718 27098 27770
rect 27110 27718 27162 27770
rect 27174 27718 27226 27770
rect 27238 27718 27290 27770
rect 3658 27174 3710 27226
rect 3722 27174 3774 27226
rect 3786 27174 3838 27226
rect 3850 27174 3902 27226
rect 3914 27174 3966 27226
rect 3978 27174 4030 27226
rect 11658 27174 11710 27226
rect 11722 27174 11774 27226
rect 11786 27174 11838 27226
rect 11850 27174 11902 27226
rect 11914 27174 11966 27226
rect 11978 27174 12030 27226
rect 19658 27174 19710 27226
rect 19722 27174 19774 27226
rect 19786 27174 19838 27226
rect 19850 27174 19902 27226
rect 19914 27174 19966 27226
rect 19978 27174 20030 27226
rect 27658 27174 27710 27226
rect 27722 27174 27774 27226
rect 27786 27174 27838 27226
rect 27850 27174 27902 27226
rect 27914 27174 27966 27226
rect 27978 27174 28030 27226
rect 2918 26630 2970 26682
rect 2982 26630 3034 26682
rect 3046 26630 3098 26682
rect 3110 26630 3162 26682
rect 3174 26630 3226 26682
rect 3238 26630 3290 26682
rect 10918 26630 10970 26682
rect 10982 26630 11034 26682
rect 11046 26630 11098 26682
rect 11110 26630 11162 26682
rect 11174 26630 11226 26682
rect 11238 26630 11290 26682
rect 18918 26630 18970 26682
rect 18982 26630 19034 26682
rect 19046 26630 19098 26682
rect 19110 26630 19162 26682
rect 19174 26630 19226 26682
rect 19238 26630 19290 26682
rect 26918 26630 26970 26682
rect 26982 26630 27034 26682
rect 27046 26630 27098 26682
rect 27110 26630 27162 26682
rect 27174 26630 27226 26682
rect 27238 26630 27290 26682
rect 3658 26086 3710 26138
rect 3722 26086 3774 26138
rect 3786 26086 3838 26138
rect 3850 26086 3902 26138
rect 3914 26086 3966 26138
rect 3978 26086 4030 26138
rect 11658 26086 11710 26138
rect 11722 26086 11774 26138
rect 11786 26086 11838 26138
rect 11850 26086 11902 26138
rect 11914 26086 11966 26138
rect 11978 26086 12030 26138
rect 19658 26086 19710 26138
rect 19722 26086 19774 26138
rect 19786 26086 19838 26138
rect 19850 26086 19902 26138
rect 19914 26086 19966 26138
rect 19978 26086 20030 26138
rect 27658 26086 27710 26138
rect 27722 26086 27774 26138
rect 27786 26086 27838 26138
rect 27850 26086 27902 26138
rect 27914 26086 27966 26138
rect 27978 26086 28030 26138
rect 2918 25542 2970 25594
rect 2982 25542 3034 25594
rect 3046 25542 3098 25594
rect 3110 25542 3162 25594
rect 3174 25542 3226 25594
rect 3238 25542 3290 25594
rect 10918 25542 10970 25594
rect 10982 25542 11034 25594
rect 11046 25542 11098 25594
rect 11110 25542 11162 25594
rect 11174 25542 11226 25594
rect 11238 25542 11290 25594
rect 18918 25542 18970 25594
rect 18982 25542 19034 25594
rect 19046 25542 19098 25594
rect 19110 25542 19162 25594
rect 19174 25542 19226 25594
rect 19238 25542 19290 25594
rect 26918 25542 26970 25594
rect 26982 25542 27034 25594
rect 27046 25542 27098 25594
rect 27110 25542 27162 25594
rect 27174 25542 27226 25594
rect 27238 25542 27290 25594
rect 1216 25168 1268 25220
rect 2504 25100 2556 25152
rect 3658 24998 3710 25050
rect 3722 24998 3774 25050
rect 3786 24998 3838 25050
rect 3850 24998 3902 25050
rect 3914 24998 3966 25050
rect 3978 24998 4030 25050
rect 11658 24998 11710 25050
rect 11722 24998 11774 25050
rect 11786 24998 11838 25050
rect 11850 24998 11902 25050
rect 11914 24998 11966 25050
rect 11978 24998 12030 25050
rect 19658 24998 19710 25050
rect 19722 24998 19774 25050
rect 19786 24998 19838 25050
rect 19850 24998 19902 25050
rect 19914 24998 19966 25050
rect 19978 24998 20030 25050
rect 27658 24998 27710 25050
rect 27722 24998 27774 25050
rect 27786 24998 27838 25050
rect 27850 24998 27902 25050
rect 27914 24998 27966 25050
rect 27978 24998 28030 25050
rect 1308 24760 1360 24812
rect 2688 24556 2740 24608
rect 2918 24454 2970 24506
rect 2982 24454 3034 24506
rect 3046 24454 3098 24506
rect 3110 24454 3162 24506
rect 3174 24454 3226 24506
rect 3238 24454 3290 24506
rect 10918 24454 10970 24506
rect 10982 24454 11034 24506
rect 11046 24454 11098 24506
rect 11110 24454 11162 24506
rect 11174 24454 11226 24506
rect 11238 24454 11290 24506
rect 18918 24454 18970 24506
rect 18982 24454 19034 24506
rect 19046 24454 19098 24506
rect 19110 24454 19162 24506
rect 19174 24454 19226 24506
rect 19238 24454 19290 24506
rect 26918 24454 26970 24506
rect 26982 24454 27034 24506
rect 27046 24454 27098 24506
rect 27110 24454 27162 24506
rect 27174 24454 27226 24506
rect 27238 24454 27290 24506
rect 5448 24216 5500 24268
rect 1308 24148 1360 24200
rect 6828 24191 6880 24200
rect 6828 24157 6837 24191
rect 6837 24157 6871 24191
rect 6871 24157 6880 24191
rect 6828 24148 6880 24157
rect 6920 24080 6972 24132
rect 7104 24123 7156 24132
rect 7104 24089 7113 24123
rect 7113 24089 7147 24123
rect 7147 24089 7156 24123
rect 7104 24080 7156 24089
rect 2044 24012 2096 24064
rect 8392 24012 8444 24064
rect 3658 23910 3710 23962
rect 3722 23910 3774 23962
rect 3786 23910 3838 23962
rect 3850 23910 3902 23962
rect 3914 23910 3966 23962
rect 3978 23910 4030 23962
rect 11658 23910 11710 23962
rect 11722 23910 11774 23962
rect 11786 23910 11838 23962
rect 11850 23910 11902 23962
rect 11914 23910 11966 23962
rect 11978 23910 12030 23962
rect 19658 23910 19710 23962
rect 19722 23910 19774 23962
rect 19786 23910 19838 23962
rect 19850 23910 19902 23962
rect 19914 23910 19966 23962
rect 19978 23910 20030 23962
rect 27658 23910 27710 23962
rect 27722 23910 27774 23962
rect 27786 23910 27838 23962
rect 27850 23910 27902 23962
rect 27914 23910 27966 23962
rect 27978 23910 28030 23962
rect 6828 23808 6880 23860
rect 1308 23672 1360 23724
rect 2688 23672 2740 23724
rect 2780 23604 2832 23656
rect 3424 23672 3476 23724
rect 3792 23672 3844 23724
rect 5448 23672 5500 23724
rect 3700 23604 3752 23656
rect 6920 23672 6972 23724
rect 7840 23715 7892 23724
rect 7840 23681 7849 23715
rect 7849 23681 7883 23715
rect 7883 23681 7892 23715
rect 7840 23672 7892 23681
rect 7932 23715 7984 23724
rect 7932 23681 7941 23715
rect 7941 23681 7975 23715
rect 7975 23681 7984 23715
rect 7932 23672 7984 23681
rect 8392 23715 8444 23724
rect 8392 23681 8401 23715
rect 8401 23681 8435 23715
rect 8435 23681 8444 23715
rect 8392 23672 8444 23681
rect 6736 23604 6788 23656
rect 7656 23647 7708 23656
rect 7656 23613 7665 23647
rect 7665 23613 7699 23647
rect 7699 23613 7708 23647
rect 7656 23604 7708 23613
rect 1400 23536 1452 23588
rect 2504 23536 2556 23588
rect 1952 23468 2004 23520
rect 2596 23468 2648 23520
rect 3424 23511 3476 23520
rect 3424 23477 3433 23511
rect 3433 23477 3467 23511
rect 3467 23477 3476 23511
rect 3424 23468 3476 23477
rect 4252 23536 4304 23588
rect 9036 23536 9088 23588
rect 5632 23468 5684 23520
rect 7104 23468 7156 23520
rect 7748 23468 7800 23520
rect 8760 23511 8812 23520
rect 8760 23477 8769 23511
rect 8769 23477 8803 23511
rect 8803 23477 8812 23511
rect 8760 23468 8812 23477
rect 2918 23366 2970 23418
rect 2982 23366 3034 23418
rect 3046 23366 3098 23418
rect 3110 23366 3162 23418
rect 3174 23366 3226 23418
rect 3238 23366 3290 23418
rect 10918 23366 10970 23418
rect 10982 23366 11034 23418
rect 11046 23366 11098 23418
rect 11110 23366 11162 23418
rect 11174 23366 11226 23418
rect 11238 23366 11290 23418
rect 18918 23366 18970 23418
rect 18982 23366 19034 23418
rect 19046 23366 19098 23418
rect 19110 23366 19162 23418
rect 19174 23366 19226 23418
rect 19238 23366 19290 23418
rect 26918 23366 26970 23418
rect 26982 23366 27034 23418
rect 27046 23366 27098 23418
rect 27110 23366 27162 23418
rect 27174 23366 27226 23418
rect 27238 23366 27290 23418
rect 1768 23264 1820 23316
rect 3332 23196 3384 23248
rect 3424 23196 3476 23248
rect 2504 23128 2556 23180
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 2320 23060 2372 23112
rect 2412 23103 2464 23112
rect 2412 23069 2421 23103
rect 2421 23069 2455 23103
rect 2455 23069 2464 23103
rect 2412 23060 2464 23069
rect 2596 23103 2648 23112
rect 2596 23069 2605 23103
rect 2605 23069 2639 23103
rect 2639 23069 2648 23103
rect 2596 23060 2648 23069
rect 2872 23060 2924 23112
rect 4712 23264 4764 23316
rect 7656 23264 7708 23316
rect 7932 23264 7984 23316
rect 5632 23196 5684 23248
rect 3792 23103 3844 23112
rect 3792 23069 3801 23103
rect 3801 23069 3835 23103
rect 3835 23069 3844 23103
rect 3792 23060 3844 23069
rect 4068 23103 4120 23112
rect 4068 23069 4077 23103
rect 4077 23069 4111 23103
rect 4111 23069 4120 23103
rect 4068 23060 4120 23069
rect 4252 23103 4304 23112
rect 4252 23069 4261 23103
rect 4261 23069 4295 23103
rect 4295 23069 4304 23103
rect 4252 23060 4304 23069
rect 4712 23103 4764 23112
rect 4712 23069 4721 23103
rect 4721 23069 4755 23103
rect 4755 23069 4764 23103
rect 4712 23060 4764 23069
rect 2504 22924 2556 22976
rect 3700 22992 3752 23044
rect 3516 22924 3568 22976
rect 4160 22967 4212 22976
rect 4160 22933 4169 22967
rect 4169 22933 4203 22967
rect 4203 22933 4212 22967
rect 4160 22924 4212 22933
rect 4252 22924 4304 22976
rect 6368 23128 6420 23180
rect 6920 23171 6972 23180
rect 6920 23137 6929 23171
rect 6929 23137 6963 23171
rect 6963 23137 6972 23171
rect 6920 23128 6972 23137
rect 8116 23239 8168 23248
rect 8116 23205 8125 23239
rect 8125 23205 8159 23239
rect 8159 23205 8168 23239
rect 8116 23196 8168 23205
rect 8484 23128 8536 23180
rect 6828 23103 6880 23112
rect 6828 23069 6837 23103
rect 6837 23069 6871 23103
rect 6871 23069 6880 23103
rect 6828 23060 6880 23069
rect 7104 23103 7156 23112
rect 7104 23069 7113 23103
rect 7113 23069 7147 23103
rect 7147 23069 7156 23103
rect 7104 23060 7156 23069
rect 7196 23103 7248 23112
rect 7196 23069 7205 23103
rect 7205 23069 7239 23103
rect 7239 23069 7248 23103
rect 7196 23060 7248 23069
rect 7748 23103 7800 23112
rect 7748 23069 7757 23103
rect 7757 23069 7791 23103
rect 7791 23069 7800 23103
rect 7748 23060 7800 23069
rect 7564 22992 7616 23044
rect 8944 22924 8996 22976
rect 3658 22822 3710 22874
rect 3722 22822 3774 22874
rect 3786 22822 3838 22874
rect 3850 22822 3902 22874
rect 3914 22822 3966 22874
rect 3978 22822 4030 22874
rect 11658 22822 11710 22874
rect 11722 22822 11774 22874
rect 11786 22822 11838 22874
rect 11850 22822 11902 22874
rect 11914 22822 11966 22874
rect 11978 22822 12030 22874
rect 19658 22822 19710 22874
rect 19722 22822 19774 22874
rect 19786 22822 19838 22874
rect 19850 22822 19902 22874
rect 19914 22822 19966 22874
rect 19978 22822 20030 22874
rect 27658 22822 27710 22874
rect 27722 22822 27774 22874
rect 27786 22822 27838 22874
rect 27850 22822 27902 22874
rect 27914 22822 27966 22874
rect 27978 22822 28030 22874
rect 2872 22720 2924 22772
rect 3424 22720 3476 22772
rect 7104 22720 7156 22772
rect 7472 22720 7524 22772
rect 1216 22584 1268 22636
rect 1952 22584 2004 22636
rect 6184 22652 6236 22704
rect 7196 22652 7248 22704
rect 2228 22627 2280 22636
rect 2228 22593 2237 22627
rect 2237 22593 2271 22627
rect 2271 22593 2280 22627
rect 2228 22584 2280 22593
rect 2688 22584 2740 22636
rect 3976 22584 4028 22636
rect 7748 22584 7800 22636
rect 7932 22627 7984 22636
rect 7932 22593 7941 22627
rect 7941 22593 7975 22627
rect 7975 22593 7984 22627
rect 7932 22584 7984 22593
rect 28080 22627 28132 22636
rect 28080 22593 28089 22627
rect 28089 22593 28123 22627
rect 28123 22593 28132 22627
rect 28080 22584 28132 22593
rect 2044 22516 2096 22568
rect 2780 22448 2832 22500
rect 2044 22380 2096 22432
rect 2596 22380 2648 22432
rect 28356 22559 28408 22568
rect 28356 22525 28365 22559
rect 28365 22525 28399 22559
rect 28399 22525 28408 22559
rect 28356 22516 28408 22525
rect 7840 22448 7892 22500
rect 6368 22380 6420 22432
rect 2918 22278 2970 22330
rect 2982 22278 3034 22330
rect 3046 22278 3098 22330
rect 3110 22278 3162 22330
rect 3174 22278 3226 22330
rect 3238 22278 3290 22330
rect 10918 22278 10970 22330
rect 10982 22278 11034 22330
rect 11046 22278 11098 22330
rect 11110 22278 11162 22330
rect 11174 22278 11226 22330
rect 11238 22278 11290 22330
rect 18918 22278 18970 22330
rect 18982 22278 19034 22330
rect 19046 22278 19098 22330
rect 19110 22278 19162 22330
rect 19174 22278 19226 22330
rect 19238 22278 19290 22330
rect 26918 22278 26970 22330
rect 26982 22278 27034 22330
rect 27046 22278 27098 22330
rect 27110 22278 27162 22330
rect 27174 22278 27226 22330
rect 27238 22278 27290 22330
rect 2412 22176 2464 22228
rect 3240 22176 3292 22228
rect 3424 22176 3476 22228
rect 5448 22176 5500 22228
rect 7932 22176 7984 22228
rect 7564 22108 7616 22160
rect 2780 22040 2832 22092
rect 2596 21972 2648 22024
rect 4160 22040 4212 22092
rect 4896 22040 4948 22092
rect 1216 21904 1268 21956
rect 2780 21947 2832 21956
rect 2780 21913 2789 21947
rect 2789 21913 2823 21947
rect 2823 21913 2832 21947
rect 2780 21904 2832 21913
rect 1860 21836 1912 21888
rect 2504 21836 2556 21888
rect 4068 21947 4120 21956
rect 4068 21913 4077 21947
rect 4077 21913 4111 21947
rect 4111 21913 4120 21947
rect 4068 21904 4120 21913
rect 3424 21836 3476 21888
rect 3976 21836 4028 21888
rect 4896 21904 4948 21956
rect 5448 22015 5500 22024
rect 5448 21981 5457 22015
rect 5457 21981 5491 22015
rect 5491 21981 5500 22015
rect 5448 21972 5500 21981
rect 5724 22040 5776 22092
rect 5632 22015 5684 22024
rect 5632 21981 5641 22015
rect 5641 21981 5675 22015
rect 5675 21981 5684 22015
rect 5632 21972 5684 21981
rect 5908 21972 5960 22024
rect 6184 22015 6236 22024
rect 6184 21981 6193 22015
rect 6193 21981 6227 22015
rect 6227 21981 6236 22015
rect 6184 21972 6236 21981
rect 6368 22015 6420 22024
rect 8760 22040 8812 22092
rect 6368 21981 6401 22015
rect 6401 21981 6420 22015
rect 6368 21972 6420 21981
rect 6920 22015 6972 22024
rect 6920 21981 6929 22015
rect 6929 21981 6963 22015
rect 6963 21981 6972 22015
rect 6920 21972 6972 21981
rect 5356 21836 5408 21888
rect 5816 21879 5868 21888
rect 5816 21845 5825 21879
rect 5825 21845 5859 21879
rect 5859 21845 5868 21879
rect 5816 21836 5868 21845
rect 6092 21904 6144 21956
rect 9036 21972 9088 22024
rect 6552 21879 6604 21888
rect 6552 21845 6561 21879
rect 6561 21845 6595 21879
rect 6595 21845 6604 21879
rect 6552 21836 6604 21845
rect 6644 21879 6696 21888
rect 6644 21845 6653 21879
rect 6653 21845 6687 21879
rect 6687 21845 6696 21879
rect 6644 21836 6696 21845
rect 8576 21836 8628 21888
rect 9496 21836 9548 21888
rect 3658 21734 3710 21786
rect 3722 21734 3774 21786
rect 3786 21734 3838 21786
rect 3850 21734 3902 21786
rect 3914 21734 3966 21786
rect 3978 21734 4030 21786
rect 11658 21734 11710 21786
rect 11722 21734 11774 21786
rect 11786 21734 11838 21786
rect 11850 21734 11902 21786
rect 11914 21734 11966 21786
rect 11978 21734 12030 21786
rect 19658 21734 19710 21786
rect 19722 21734 19774 21786
rect 19786 21734 19838 21786
rect 19850 21734 19902 21786
rect 19914 21734 19966 21786
rect 19978 21734 20030 21786
rect 27658 21734 27710 21786
rect 27722 21734 27774 21786
rect 27786 21734 27838 21786
rect 27850 21734 27902 21786
rect 27914 21734 27966 21786
rect 27978 21734 28030 21786
rect 2136 21632 2188 21684
rect 1308 21496 1360 21548
rect 3240 21564 3292 21616
rect 4896 21675 4948 21684
rect 4896 21641 4905 21675
rect 4905 21641 4939 21675
rect 4939 21641 4948 21675
rect 4896 21632 4948 21641
rect 6092 21632 6144 21684
rect 6920 21632 6972 21684
rect 5724 21564 5776 21616
rect 5816 21564 5868 21616
rect 2688 21539 2740 21548
rect 2688 21505 2697 21539
rect 2697 21505 2731 21539
rect 2731 21505 2740 21539
rect 2688 21496 2740 21505
rect 2596 21428 2648 21480
rect 3608 21496 3660 21548
rect 1216 21360 1268 21412
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 2412 21292 2464 21344
rect 2780 21292 2832 21344
rect 5908 21335 5960 21344
rect 5908 21301 5917 21335
rect 5917 21301 5951 21335
rect 5951 21301 5960 21335
rect 5908 21292 5960 21301
rect 6460 21496 6512 21548
rect 8484 21607 8536 21616
rect 8484 21573 8493 21607
rect 8493 21573 8527 21607
rect 8527 21573 8536 21607
rect 8484 21564 8536 21573
rect 7748 21539 7800 21548
rect 7748 21505 7757 21539
rect 7757 21505 7791 21539
rect 7791 21505 7800 21539
rect 7748 21496 7800 21505
rect 7932 21539 7984 21548
rect 7932 21505 7941 21539
rect 7941 21505 7975 21539
rect 7975 21505 7984 21539
rect 7932 21496 7984 21505
rect 7012 21360 7064 21412
rect 8300 21360 8352 21412
rect 6552 21292 6604 21344
rect 7196 21335 7248 21344
rect 7196 21301 7205 21335
rect 7205 21301 7239 21335
rect 7239 21301 7248 21335
rect 7196 21292 7248 21301
rect 2918 21190 2970 21242
rect 2982 21190 3034 21242
rect 3046 21190 3098 21242
rect 3110 21190 3162 21242
rect 3174 21190 3226 21242
rect 3238 21190 3290 21242
rect 10918 21190 10970 21242
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 11238 21190 11290 21242
rect 18918 21190 18970 21242
rect 18982 21190 19034 21242
rect 19046 21190 19098 21242
rect 19110 21190 19162 21242
rect 19174 21190 19226 21242
rect 19238 21190 19290 21242
rect 26918 21190 26970 21242
rect 26982 21190 27034 21242
rect 27046 21190 27098 21242
rect 27110 21190 27162 21242
rect 27174 21190 27226 21242
rect 27238 21190 27290 21242
rect 3516 21088 3568 21140
rect 5356 21131 5408 21140
rect 5356 21097 5365 21131
rect 5365 21097 5399 21131
rect 5399 21097 5408 21131
rect 5356 21088 5408 21097
rect 5908 21088 5960 21140
rect 8300 21020 8352 21072
rect 8944 21020 8996 21072
rect 2780 20952 2832 21004
rect 1308 20884 1360 20936
rect 1952 20816 2004 20868
rect 2780 20816 2832 20868
rect 2964 20927 3016 20936
rect 2964 20893 2973 20927
rect 2973 20893 3007 20927
rect 3007 20893 3016 20927
rect 2964 20884 3016 20893
rect 3516 20952 3568 21004
rect 9128 20952 9180 21004
rect 4252 20927 4304 20936
rect 4252 20893 4261 20927
rect 4261 20893 4295 20927
rect 4295 20893 4304 20927
rect 4252 20884 4304 20893
rect 5448 20927 5500 20936
rect 5448 20893 5457 20927
rect 5457 20893 5491 20927
rect 5491 20893 5500 20927
rect 5448 20884 5500 20893
rect 7012 20927 7064 20936
rect 7012 20893 7021 20927
rect 7021 20893 7055 20927
rect 7055 20893 7064 20927
rect 7012 20884 7064 20893
rect 7196 20884 7248 20936
rect 7380 20927 7432 20936
rect 7380 20893 7389 20927
rect 7389 20893 7423 20927
rect 7423 20893 7432 20927
rect 7380 20884 7432 20893
rect 3056 20816 3108 20868
rect 12900 20816 12952 20868
rect 3332 20748 3384 20800
rect 4160 20791 4212 20800
rect 4160 20757 4169 20791
rect 4169 20757 4203 20791
rect 4203 20757 4212 20791
rect 4160 20748 4212 20757
rect 4528 20791 4580 20800
rect 4528 20757 4537 20791
rect 4537 20757 4571 20791
rect 4571 20757 4580 20791
rect 4528 20748 4580 20757
rect 9864 20748 9916 20800
rect 3658 20646 3710 20698
rect 3722 20646 3774 20698
rect 3786 20646 3838 20698
rect 3850 20646 3902 20698
rect 3914 20646 3966 20698
rect 3978 20646 4030 20698
rect 11658 20646 11710 20698
rect 11722 20646 11774 20698
rect 11786 20646 11838 20698
rect 11850 20646 11902 20698
rect 11914 20646 11966 20698
rect 11978 20646 12030 20698
rect 19658 20646 19710 20698
rect 19722 20646 19774 20698
rect 19786 20646 19838 20698
rect 19850 20646 19902 20698
rect 19914 20646 19966 20698
rect 19978 20646 20030 20698
rect 27658 20646 27710 20698
rect 27722 20646 27774 20698
rect 27786 20646 27838 20698
rect 27850 20646 27902 20698
rect 27914 20646 27966 20698
rect 27978 20646 28030 20698
rect 3056 20544 3108 20596
rect 4252 20476 4304 20528
rect 5448 20476 5500 20528
rect 1308 20408 1360 20460
rect 2228 20408 2280 20460
rect 2688 20408 2740 20460
rect 8944 20408 8996 20460
rect 9128 20451 9180 20460
rect 9128 20417 9138 20451
rect 9138 20417 9172 20451
rect 9172 20417 9180 20451
rect 9128 20408 9180 20417
rect 6736 20340 6788 20392
rect 1676 20272 1728 20324
rect 2596 20272 2648 20324
rect 9588 20272 9640 20324
rect 10048 20272 10100 20324
rect 3332 20204 3384 20256
rect 5448 20204 5500 20256
rect 10232 20204 10284 20256
rect 21916 20204 21968 20256
rect 24032 20204 24084 20256
rect 2918 20102 2970 20154
rect 2982 20102 3034 20154
rect 3046 20102 3098 20154
rect 3110 20102 3162 20154
rect 3174 20102 3226 20154
rect 3238 20102 3290 20154
rect 10918 20102 10970 20154
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 11238 20102 11290 20154
rect 18918 20102 18970 20154
rect 18982 20102 19034 20154
rect 19046 20102 19098 20154
rect 19110 20102 19162 20154
rect 19174 20102 19226 20154
rect 19238 20102 19290 20154
rect 26918 20102 26970 20154
rect 26982 20102 27034 20154
rect 27046 20102 27098 20154
rect 27110 20102 27162 20154
rect 27174 20102 27226 20154
rect 27238 20102 27290 20154
rect 6828 20000 6880 20052
rect 7472 20043 7524 20052
rect 7472 20009 7481 20043
rect 7481 20009 7515 20043
rect 7515 20009 7524 20043
rect 7472 20000 7524 20009
rect 10140 20000 10192 20052
rect 23204 20000 23256 20052
rect 23572 20000 23624 20052
rect 28080 20000 28132 20052
rect 3516 19932 3568 19984
rect 4528 19932 4580 19984
rect 5816 19864 5868 19916
rect 1308 19796 1360 19848
rect 2596 19796 2648 19848
rect 6000 19796 6052 19848
rect 8024 19864 8076 19916
rect 8208 19864 8260 19916
rect 9864 19864 9916 19916
rect 12440 19864 12492 19916
rect 1952 19728 2004 19780
rect 4068 19728 4120 19780
rect 6184 19728 6236 19780
rect 9772 19839 9824 19848
rect 9772 19805 9781 19839
rect 9781 19805 9815 19839
rect 9815 19805 9824 19839
rect 9772 19796 9824 19805
rect 10048 19839 10100 19848
rect 10048 19805 10057 19839
rect 10057 19805 10091 19839
rect 10091 19805 10100 19839
rect 10048 19796 10100 19805
rect 10232 19839 10284 19848
rect 10232 19805 10241 19839
rect 10241 19805 10275 19839
rect 10275 19805 10284 19839
rect 10232 19796 10284 19805
rect 14464 19796 14516 19848
rect 9404 19771 9456 19780
rect 9404 19737 9413 19771
rect 9413 19737 9447 19771
rect 9447 19737 9456 19771
rect 9404 19728 9456 19737
rect 9588 19771 9640 19780
rect 9588 19737 9623 19771
rect 9623 19737 9640 19771
rect 9588 19728 9640 19737
rect 12624 19728 12676 19780
rect 3056 19660 3108 19712
rect 3516 19660 3568 19712
rect 12532 19703 12584 19712
rect 12532 19669 12541 19703
rect 12541 19669 12575 19703
rect 12575 19669 12584 19703
rect 12532 19660 12584 19669
rect 18144 19703 18196 19712
rect 18144 19669 18153 19703
rect 18153 19669 18187 19703
rect 18187 19669 18196 19703
rect 18144 19660 18196 19669
rect 19340 19660 19392 19712
rect 23296 19975 23348 19984
rect 23296 19941 23305 19975
rect 23305 19941 23339 19975
rect 23339 19941 23348 19975
rect 23296 19932 23348 19941
rect 22836 19907 22888 19916
rect 22836 19873 22845 19907
rect 22845 19873 22879 19907
rect 22879 19873 22888 19907
rect 22836 19864 22888 19873
rect 23020 19864 23072 19916
rect 21916 19796 21968 19848
rect 22192 19796 22244 19848
rect 23388 19728 23440 19780
rect 23572 19839 23624 19848
rect 23572 19805 23581 19839
rect 23581 19805 23615 19839
rect 23615 19805 23624 19839
rect 23572 19796 23624 19805
rect 24308 19728 24360 19780
rect 22192 19660 22244 19712
rect 23480 19703 23532 19712
rect 23480 19669 23489 19703
rect 23489 19669 23523 19703
rect 23523 19669 23532 19703
rect 23480 19660 23532 19669
rect 24216 19660 24268 19712
rect 3658 19558 3710 19610
rect 3722 19558 3774 19610
rect 3786 19558 3838 19610
rect 3850 19558 3902 19610
rect 3914 19558 3966 19610
rect 3978 19558 4030 19610
rect 11658 19558 11710 19610
rect 11722 19558 11774 19610
rect 11786 19558 11838 19610
rect 11850 19558 11902 19610
rect 11914 19558 11966 19610
rect 11978 19558 12030 19610
rect 19658 19558 19710 19610
rect 19722 19558 19774 19610
rect 19786 19558 19838 19610
rect 19850 19558 19902 19610
rect 19914 19558 19966 19610
rect 19978 19558 20030 19610
rect 27658 19558 27710 19610
rect 27722 19558 27774 19610
rect 27786 19558 27838 19610
rect 27850 19558 27902 19610
rect 27914 19558 27966 19610
rect 27978 19558 28030 19610
rect 2688 19456 2740 19508
rect 3056 19456 3108 19508
rect 3976 19456 4028 19508
rect 6184 19499 6236 19508
rect 6184 19465 6193 19499
rect 6193 19465 6227 19499
rect 6227 19465 6236 19499
rect 6184 19456 6236 19465
rect 6736 19456 6788 19508
rect 4528 19388 4580 19440
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 2688 19320 2740 19372
rect 2872 19320 2924 19372
rect 3424 19320 3476 19372
rect 4068 19320 4120 19372
rect 3056 19252 3108 19304
rect 3700 19252 3752 19304
rect 3792 19295 3844 19304
rect 3792 19261 3801 19295
rect 3801 19261 3835 19295
rect 3835 19261 3844 19295
rect 3792 19252 3844 19261
rect 3976 19252 4028 19304
rect 5632 19363 5684 19372
rect 5632 19329 5641 19363
rect 5641 19329 5675 19363
rect 5675 19329 5684 19363
rect 5632 19320 5684 19329
rect 5816 19363 5868 19372
rect 5816 19329 5825 19363
rect 5825 19329 5859 19363
rect 5859 19329 5868 19363
rect 5816 19320 5868 19329
rect 5908 19363 5960 19372
rect 5908 19329 5917 19363
rect 5917 19329 5951 19363
rect 5951 19329 5960 19363
rect 5908 19320 5960 19329
rect 6000 19363 6052 19372
rect 6000 19329 6009 19363
rect 6009 19329 6043 19363
rect 6043 19329 6052 19363
rect 6000 19320 6052 19329
rect 6368 19320 6420 19372
rect 6736 19363 6788 19372
rect 6736 19329 6745 19363
rect 6745 19329 6779 19363
rect 6779 19329 6788 19363
rect 6736 19320 6788 19329
rect 7472 19388 7524 19440
rect 8208 19499 8260 19508
rect 8208 19465 8217 19499
rect 8217 19465 8251 19499
rect 8251 19465 8260 19499
rect 8208 19456 8260 19465
rect 9404 19456 9456 19508
rect 9772 19456 9824 19508
rect 12532 19456 12584 19508
rect 23388 19456 23440 19508
rect 6828 19295 6880 19304
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 8024 19363 8076 19372
rect 8024 19329 8033 19363
rect 8033 19329 8067 19363
rect 8067 19329 8076 19363
rect 8024 19320 8076 19329
rect 9864 19388 9916 19440
rect 18144 19431 18196 19440
rect 18144 19397 18153 19431
rect 18153 19397 18187 19431
rect 18187 19397 18196 19431
rect 18144 19388 18196 19397
rect 18788 19388 18840 19440
rect 7932 19295 7984 19304
rect 6828 19252 6880 19261
rect 3240 19227 3292 19236
rect 3240 19193 3249 19227
rect 3249 19193 3283 19227
rect 3283 19193 3292 19227
rect 3240 19184 3292 19193
rect 3332 19184 3384 19236
rect 2136 19116 2188 19168
rect 2964 19116 3016 19168
rect 3424 19159 3476 19168
rect 3424 19125 3433 19159
rect 3433 19125 3467 19159
rect 3467 19125 3476 19159
rect 3424 19116 3476 19125
rect 3608 19116 3660 19168
rect 5632 19184 5684 19236
rect 7932 19261 7941 19295
rect 7941 19261 7975 19295
rect 7975 19261 7984 19295
rect 7932 19252 7984 19261
rect 10232 19320 10284 19372
rect 15108 19320 15160 19372
rect 15292 19363 15344 19372
rect 15292 19329 15301 19363
rect 15301 19329 15335 19363
rect 15335 19329 15344 19363
rect 15292 19320 15344 19329
rect 16856 19320 16908 19372
rect 22744 19363 22796 19372
rect 22744 19329 22753 19363
rect 22753 19329 22787 19363
rect 22787 19329 22796 19363
rect 22744 19320 22796 19329
rect 23296 19388 23348 19440
rect 24032 19388 24084 19440
rect 23020 19363 23072 19372
rect 23020 19329 23029 19363
rect 23029 19329 23063 19363
rect 23063 19329 23072 19363
rect 23020 19320 23072 19329
rect 12808 19295 12860 19304
rect 12808 19261 12817 19295
rect 12817 19261 12851 19295
rect 12851 19261 12860 19295
rect 12808 19252 12860 19261
rect 12900 19295 12952 19304
rect 12900 19261 12909 19295
rect 12909 19261 12943 19295
rect 12943 19261 12952 19295
rect 12900 19252 12952 19261
rect 5540 19116 5592 19168
rect 5908 19116 5960 19168
rect 8208 19116 8260 19168
rect 9220 19116 9272 19168
rect 15476 19159 15528 19168
rect 15476 19125 15485 19159
rect 15485 19125 15519 19159
rect 15519 19125 15528 19159
rect 15476 19116 15528 19125
rect 19340 19116 19392 19168
rect 20444 19116 20496 19168
rect 2918 19014 2970 19066
rect 2982 19014 3034 19066
rect 3046 19014 3098 19066
rect 3110 19014 3162 19066
rect 3174 19014 3226 19066
rect 3238 19014 3290 19066
rect 10918 19014 10970 19066
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 11238 19014 11290 19066
rect 18918 19014 18970 19066
rect 18982 19014 19034 19066
rect 19046 19014 19098 19066
rect 19110 19014 19162 19066
rect 19174 19014 19226 19066
rect 19238 19014 19290 19066
rect 26918 19014 26970 19066
rect 26982 19014 27034 19066
rect 27046 19014 27098 19066
rect 27110 19014 27162 19066
rect 27174 19014 27226 19066
rect 27238 19014 27290 19066
rect 3240 18912 3292 18964
rect 3424 18955 3476 18964
rect 3424 18921 3433 18955
rect 3433 18921 3467 18955
rect 3467 18921 3476 18955
rect 3424 18912 3476 18921
rect 4252 18912 4304 18964
rect 12808 18912 12860 18964
rect 14464 18955 14516 18964
rect 14464 18921 14473 18955
rect 14473 18921 14507 18955
rect 14507 18921 14516 18955
rect 14464 18912 14516 18921
rect 22192 18955 22244 18964
rect 22192 18921 22201 18955
rect 22201 18921 22235 18955
rect 22235 18921 22244 18955
rect 22192 18912 22244 18921
rect 22744 18912 22796 18964
rect 23388 18955 23440 18964
rect 23388 18921 23397 18955
rect 23397 18921 23431 18955
rect 23431 18921 23440 18955
rect 23388 18912 23440 18921
rect 24308 18912 24360 18964
rect 3608 18844 3660 18896
rect 1308 18708 1360 18760
rect 2596 18776 2648 18828
rect 3148 18776 3200 18828
rect 14188 18776 14240 18828
rect 2872 18708 2924 18760
rect 3240 18708 3292 18760
rect 3516 18708 3568 18760
rect 4528 18751 4580 18760
rect 4528 18717 4537 18751
rect 4537 18717 4571 18751
rect 4571 18717 4580 18751
rect 4528 18708 4580 18717
rect 11336 18708 11388 18760
rect 12808 18708 12860 18760
rect 16856 18708 16908 18760
rect 21824 18751 21876 18760
rect 21824 18717 21833 18751
rect 21833 18717 21867 18751
rect 21867 18717 21876 18751
rect 21824 18708 21876 18717
rect 24584 18751 24636 18760
rect 24584 18717 24593 18751
rect 24593 18717 24627 18751
rect 24627 18717 24636 18751
rect 24584 18708 24636 18717
rect 2228 18640 2280 18692
rect 2688 18683 2740 18692
rect 2688 18649 2697 18683
rect 2697 18649 2731 18683
rect 2731 18649 2740 18683
rect 2688 18640 2740 18649
rect 6736 18640 6788 18692
rect 3516 18572 3568 18624
rect 3792 18615 3844 18624
rect 3792 18581 3801 18615
rect 3801 18581 3835 18615
rect 3835 18581 3844 18615
rect 3792 18572 3844 18581
rect 4436 18615 4488 18624
rect 4436 18581 4445 18615
rect 4445 18581 4479 18615
rect 4479 18581 4488 18615
rect 4436 18572 4488 18581
rect 15936 18683 15988 18692
rect 15936 18649 15945 18683
rect 15945 18649 15979 18683
rect 15979 18649 15988 18683
rect 15936 18640 15988 18649
rect 23204 18640 23256 18692
rect 23480 18640 23532 18692
rect 24492 18640 24544 18692
rect 12072 18572 12124 18624
rect 15568 18572 15620 18624
rect 22100 18572 22152 18624
rect 22376 18615 22428 18624
rect 22376 18581 22385 18615
rect 22385 18581 22419 18615
rect 22419 18581 22428 18615
rect 22376 18572 22428 18581
rect 3658 18470 3710 18522
rect 3722 18470 3774 18522
rect 3786 18470 3838 18522
rect 3850 18470 3902 18522
rect 3914 18470 3966 18522
rect 3978 18470 4030 18522
rect 11658 18470 11710 18522
rect 11722 18470 11774 18522
rect 11786 18470 11838 18522
rect 11850 18470 11902 18522
rect 11914 18470 11966 18522
rect 11978 18470 12030 18522
rect 19658 18470 19710 18522
rect 19722 18470 19774 18522
rect 19786 18470 19838 18522
rect 19850 18470 19902 18522
rect 19914 18470 19966 18522
rect 19978 18470 20030 18522
rect 27658 18470 27710 18522
rect 27722 18470 27774 18522
rect 27786 18470 27838 18522
rect 27850 18470 27902 18522
rect 27914 18470 27966 18522
rect 27978 18470 28030 18522
rect 3148 18411 3200 18420
rect 3148 18377 3157 18411
rect 3157 18377 3191 18411
rect 3191 18377 3200 18411
rect 3148 18368 3200 18377
rect 2136 18300 2188 18352
rect 2596 18300 2648 18352
rect 1308 18232 1360 18284
rect 2320 18232 2372 18284
rect 4436 18368 4488 18420
rect 3516 18300 3568 18352
rect 3424 18232 3476 18284
rect 3976 18275 4028 18284
rect 3976 18241 3985 18275
rect 3985 18241 4019 18275
rect 4019 18241 4028 18275
rect 3976 18232 4028 18241
rect 9496 18300 9548 18352
rect 10140 18300 10192 18352
rect 12072 18368 12124 18420
rect 12716 18368 12768 18420
rect 15108 18368 15160 18420
rect 22100 18368 22152 18420
rect 24492 18368 24544 18420
rect 12440 18300 12492 18352
rect 23388 18300 23440 18352
rect 9404 18275 9456 18284
rect 9404 18241 9413 18275
rect 9413 18241 9447 18275
rect 9447 18241 9456 18275
rect 9404 18232 9456 18241
rect 9588 18232 9640 18284
rect 2136 18164 2188 18216
rect 2688 18207 2740 18216
rect 2688 18173 2697 18207
rect 2697 18173 2731 18207
rect 2731 18173 2740 18207
rect 2688 18164 2740 18173
rect 2872 18164 2924 18216
rect 5540 18164 5592 18216
rect 9220 18164 9272 18216
rect 9864 18232 9916 18284
rect 3056 18139 3108 18148
rect 3056 18105 3065 18139
rect 3065 18105 3099 18139
rect 3099 18105 3108 18139
rect 3056 18096 3108 18105
rect 8484 18096 8536 18148
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 3424 18071 3476 18080
rect 3424 18037 3433 18071
rect 3433 18037 3467 18071
rect 3467 18037 3476 18071
rect 3424 18028 3476 18037
rect 9496 18028 9548 18080
rect 14188 18275 14240 18284
rect 14188 18241 14197 18275
rect 14197 18241 14231 18275
rect 14231 18241 14240 18275
rect 14188 18232 14240 18241
rect 15568 18232 15620 18284
rect 12624 18207 12676 18216
rect 12624 18173 12633 18207
rect 12633 18173 12667 18207
rect 12667 18173 12676 18207
rect 12624 18164 12676 18173
rect 12164 18096 12216 18148
rect 14464 18207 14516 18216
rect 14464 18173 14473 18207
rect 14473 18173 14507 18207
rect 14507 18173 14516 18207
rect 14464 18164 14516 18173
rect 16488 18232 16540 18284
rect 20904 18275 20956 18284
rect 20904 18241 20913 18275
rect 20913 18241 20947 18275
rect 20947 18241 20956 18275
rect 20904 18232 20956 18241
rect 22376 18232 22428 18284
rect 23388 18207 23440 18216
rect 23388 18173 23397 18207
rect 23397 18173 23431 18207
rect 23431 18173 23440 18207
rect 23388 18164 23440 18173
rect 24584 18164 24636 18216
rect 23204 18096 23256 18148
rect 18236 18028 18288 18080
rect 20812 18028 20864 18080
rect 23112 18028 23164 18080
rect 2918 17926 2970 17978
rect 2982 17926 3034 17978
rect 3046 17926 3098 17978
rect 3110 17926 3162 17978
rect 3174 17926 3226 17978
rect 3238 17926 3290 17978
rect 10918 17926 10970 17978
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 11238 17926 11290 17978
rect 18918 17926 18970 17978
rect 18982 17926 19034 17978
rect 19046 17926 19098 17978
rect 19110 17926 19162 17978
rect 19174 17926 19226 17978
rect 19238 17926 19290 17978
rect 26918 17926 26970 17978
rect 26982 17926 27034 17978
rect 27046 17926 27098 17978
rect 27110 17926 27162 17978
rect 27174 17926 27226 17978
rect 27238 17926 27290 17978
rect 2320 17867 2372 17876
rect 2320 17833 2329 17867
rect 2329 17833 2363 17867
rect 2363 17833 2372 17867
rect 2320 17824 2372 17833
rect 4160 17824 4212 17876
rect 7380 17824 7432 17876
rect 14464 17824 14516 17876
rect 15936 17824 15988 17876
rect 16488 17824 16540 17876
rect 3424 17688 3476 17740
rect 6828 17731 6880 17740
rect 6828 17697 6837 17731
rect 6837 17697 6871 17731
rect 6871 17697 6880 17731
rect 6828 17688 6880 17697
rect 14740 17688 14792 17740
rect 15476 17688 15528 17740
rect 18880 17688 18932 17740
rect 20720 17688 20772 17740
rect 21180 17824 21232 17876
rect 21824 17824 21876 17876
rect 2228 17663 2280 17672
rect 2228 17629 2237 17663
rect 2237 17629 2271 17663
rect 2271 17629 2280 17663
rect 2228 17620 2280 17629
rect 3056 17663 3108 17672
rect 3056 17629 3065 17663
rect 3065 17629 3099 17663
rect 3099 17629 3108 17663
rect 3056 17620 3108 17629
rect 4160 17620 4212 17672
rect 5816 17663 5868 17672
rect 5816 17629 5825 17663
rect 5825 17629 5859 17663
rect 5859 17629 5868 17663
rect 5816 17620 5868 17629
rect 1216 17552 1268 17604
rect 4528 17552 4580 17604
rect 5724 17552 5776 17604
rect 6736 17663 6788 17672
rect 6736 17629 6745 17663
rect 6745 17629 6779 17663
rect 6779 17629 6788 17663
rect 6736 17620 6788 17629
rect 6920 17620 6972 17672
rect 7104 17663 7156 17672
rect 7104 17629 7113 17663
rect 7113 17629 7147 17663
rect 7147 17629 7156 17663
rect 7104 17620 7156 17629
rect 14556 17620 14608 17672
rect 24124 17688 24176 17740
rect 7748 17552 7800 17604
rect 15108 17595 15160 17604
rect 15108 17561 15117 17595
rect 15117 17561 15151 17595
rect 15151 17561 15160 17595
rect 15108 17552 15160 17561
rect 16212 17552 16264 17604
rect 18696 17552 18748 17604
rect 6368 17484 6420 17536
rect 15844 17527 15896 17536
rect 15844 17493 15853 17527
rect 15853 17493 15887 17527
rect 15887 17493 15896 17527
rect 15844 17484 15896 17493
rect 17684 17527 17736 17536
rect 17684 17493 17693 17527
rect 17693 17493 17727 17527
rect 17727 17493 17736 17527
rect 17684 17484 17736 17493
rect 18604 17484 18656 17536
rect 20812 17484 20864 17536
rect 3658 17382 3710 17434
rect 3722 17382 3774 17434
rect 3786 17382 3838 17434
rect 3850 17382 3902 17434
rect 3914 17382 3966 17434
rect 3978 17382 4030 17434
rect 11658 17382 11710 17434
rect 11722 17382 11774 17434
rect 11786 17382 11838 17434
rect 11850 17382 11902 17434
rect 11914 17382 11966 17434
rect 11978 17382 12030 17434
rect 19658 17382 19710 17434
rect 19722 17382 19774 17434
rect 19786 17382 19838 17434
rect 19850 17382 19902 17434
rect 19914 17382 19966 17434
rect 19978 17382 20030 17434
rect 27658 17382 27710 17434
rect 27722 17382 27774 17434
rect 27786 17382 27838 17434
rect 27850 17382 27902 17434
rect 27914 17382 27966 17434
rect 27978 17382 28030 17434
rect 7104 17323 7156 17332
rect 7104 17289 7113 17323
rect 7113 17289 7147 17323
rect 7147 17289 7156 17323
rect 7104 17280 7156 17289
rect 7748 17323 7800 17332
rect 7748 17289 7757 17323
rect 7757 17289 7791 17323
rect 7791 17289 7800 17323
rect 7748 17280 7800 17289
rect 9404 17280 9456 17332
rect 18604 17323 18656 17332
rect 18604 17289 18613 17323
rect 18613 17289 18647 17323
rect 18647 17289 18656 17323
rect 18604 17280 18656 17289
rect 1584 17212 1636 17264
rect 6276 17212 6328 17264
rect 1308 17144 1360 17196
rect 5448 17187 5500 17196
rect 5448 17153 5457 17187
rect 5457 17153 5491 17187
rect 5491 17153 5500 17187
rect 5448 17144 5500 17153
rect 6368 17187 6420 17196
rect 6368 17153 6377 17187
rect 6377 17153 6411 17187
rect 6411 17153 6420 17187
rect 6368 17144 6420 17153
rect 6828 17212 6880 17264
rect 5724 17119 5776 17128
rect 5724 17085 5733 17119
rect 5733 17085 5767 17119
rect 5767 17085 5776 17119
rect 5724 17076 5776 17085
rect 6644 17119 6696 17128
rect 6644 17085 6653 17119
rect 6653 17085 6687 17119
rect 6687 17085 6696 17119
rect 6644 17076 6696 17085
rect 6736 17119 6788 17128
rect 6736 17085 6745 17119
rect 6745 17085 6779 17119
rect 6779 17085 6788 17119
rect 7472 17187 7524 17196
rect 7472 17153 7481 17187
rect 7481 17153 7515 17187
rect 7515 17153 7524 17187
rect 7472 17144 7524 17153
rect 9036 17212 9088 17264
rect 9864 17212 9916 17264
rect 20904 17280 20956 17332
rect 24584 17323 24636 17332
rect 18880 17255 18932 17264
rect 18880 17221 18889 17255
rect 18889 17221 18923 17255
rect 18923 17221 18932 17255
rect 18880 17212 18932 17221
rect 8392 17144 8444 17196
rect 18236 17144 18288 17196
rect 21180 17187 21232 17196
rect 21180 17153 21189 17187
rect 21189 17153 21223 17187
rect 21223 17153 21232 17187
rect 21180 17144 21232 17153
rect 21824 17212 21876 17264
rect 24584 17289 24593 17323
rect 24593 17289 24627 17323
rect 24627 17289 24636 17323
rect 24584 17280 24636 17289
rect 23020 17212 23072 17264
rect 23112 17255 23164 17264
rect 23112 17221 23121 17255
rect 23121 17221 23155 17255
rect 23155 17221 23164 17255
rect 23112 17212 23164 17221
rect 6736 17076 6788 17085
rect 16856 17119 16908 17128
rect 16856 17085 16865 17119
rect 16865 17085 16899 17119
rect 16899 17085 16908 17119
rect 16856 17076 16908 17085
rect 19892 17076 19944 17128
rect 20628 17076 20680 17128
rect 24216 17144 24268 17196
rect 5816 17008 5868 17060
rect 7840 17008 7892 17060
rect 2596 16940 2648 16992
rect 3608 16940 3660 16992
rect 6828 16940 6880 16992
rect 9128 16983 9180 16992
rect 9128 16949 9137 16983
rect 9137 16949 9171 16983
rect 9171 16949 9180 16983
rect 9128 16940 9180 16949
rect 21180 16940 21232 16992
rect 23204 16940 23256 16992
rect 2918 16838 2970 16890
rect 2982 16838 3034 16890
rect 3046 16838 3098 16890
rect 3110 16838 3162 16890
rect 3174 16838 3226 16890
rect 3238 16838 3290 16890
rect 10918 16838 10970 16890
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 11238 16838 11290 16890
rect 18918 16838 18970 16890
rect 18982 16838 19034 16890
rect 19046 16838 19098 16890
rect 19110 16838 19162 16890
rect 19174 16838 19226 16890
rect 19238 16838 19290 16890
rect 26918 16838 26970 16890
rect 26982 16838 27034 16890
rect 27046 16838 27098 16890
rect 27110 16838 27162 16890
rect 27174 16838 27226 16890
rect 27238 16838 27290 16890
rect 2504 16736 2556 16788
rect 6644 16736 6696 16788
rect 1768 16668 1820 16720
rect 2596 16668 2648 16720
rect 6184 16711 6236 16720
rect 6184 16677 6193 16711
rect 6193 16677 6227 16711
rect 6227 16677 6236 16711
rect 6184 16668 6236 16677
rect 6736 16668 6788 16720
rect 7472 16736 7524 16788
rect 8576 16779 8628 16788
rect 8576 16745 8585 16779
rect 8585 16745 8619 16779
rect 8619 16745 8628 16779
rect 8576 16736 8628 16745
rect 12716 16736 12768 16788
rect 17684 16736 17736 16788
rect 18696 16779 18748 16788
rect 18696 16745 18705 16779
rect 18705 16745 18739 16779
rect 18739 16745 18748 16779
rect 18696 16736 18748 16745
rect 20720 16668 20772 16720
rect 23020 16668 23072 16720
rect 8300 16600 8352 16652
rect 9128 16600 9180 16652
rect 11336 16643 11388 16652
rect 11336 16609 11345 16643
rect 11345 16609 11379 16643
rect 11379 16609 11388 16643
rect 11336 16600 11388 16609
rect 12072 16600 12124 16652
rect 16856 16600 16908 16652
rect 17316 16600 17368 16652
rect 2780 16532 2832 16584
rect 1492 16507 1544 16516
rect 1492 16473 1501 16507
rect 1501 16473 1535 16507
rect 1535 16473 1544 16507
rect 1492 16464 1544 16473
rect 2320 16464 2372 16516
rect 3056 16507 3108 16516
rect 3056 16473 3065 16507
rect 3065 16473 3099 16507
rect 3099 16473 3108 16507
rect 3056 16464 3108 16473
rect 3424 16575 3476 16584
rect 3424 16541 3433 16575
rect 3433 16541 3467 16575
rect 3467 16541 3476 16575
rect 3424 16532 3476 16541
rect 3608 16575 3660 16584
rect 3608 16541 3617 16575
rect 3617 16541 3651 16575
rect 3651 16541 3660 16575
rect 3608 16532 3660 16541
rect 5908 16575 5960 16584
rect 5908 16541 5917 16575
rect 5917 16541 5951 16575
rect 5951 16541 5960 16575
rect 5908 16532 5960 16541
rect 6460 16575 6512 16584
rect 6460 16541 6469 16575
rect 6469 16541 6503 16575
rect 6503 16541 6512 16575
rect 6460 16532 6512 16541
rect 6552 16532 6604 16584
rect 6920 16575 6972 16584
rect 6920 16541 6929 16575
rect 6929 16541 6963 16575
rect 6963 16541 6972 16575
rect 6920 16532 6972 16541
rect 7104 16532 7156 16584
rect 8392 16575 8444 16584
rect 8392 16541 8406 16575
rect 8406 16541 8440 16575
rect 8440 16541 8444 16575
rect 8392 16532 8444 16541
rect 12716 16532 12768 16584
rect 19892 16575 19944 16584
rect 19892 16541 19901 16575
rect 19901 16541 19935 16575
rect 19935 16541 19944 16575
rect 19892 16532 19944 16541
rect 22008 16600 22060 16652
rect 23204 16600 23256 16652
rect 23480 16575 23532 16584
rect 23480 16541 23489 16575
rect 23489 16541 23523 16575
rect 23523 16541 23532 16575
rect 23480 16532 23532 16541
rect 6644 16464 6696 16516
rect 3332 16396 3384 16448
rect 8208 16507 8260 16516
rect 8208 16473 8217 16507
rect 8217 16473 8251 16507
rect 8251 16473 8260 16507
rect 8208 16464 8260 16473
rect 18236 16464 18288 16516
rect 12532 16396 12584 16448
rect 24124 16464 24176 16516
rect 3658 16294 3710 16346
rect 3722 16294 3774 16346
rect 3786 16294 3838 16346
rect 3850 16294 3902 16346
rect 3914 16294 3966 16346
rect 3978 16294 4030 16346
rect 11658 16294 11710 16346
rect 11722 16294 11774 16346
rect 11786 16294 11838 16346
rect 11850 16294 11902 16346
rect 11914 16294 11966 16346
rect 11978 16294 12030 16346
rect 19658 16294 19710 16346
rect 19722 16294 19774 16346
rect 19786 16294 19838 16346
rect 19850 16294 19902 16346
rect 19914 16294 19966 16346
rect 19978 16294 20030 16346
rect 27658 16294 27710 16346
rect 27722 16294 27774 16346
rect 27786 16294 27838 16346
rect 27850 16294 27902 16346
rect 27914 16294 27966 16346
rect 27978 16294 28030 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 2044 16192 2096 16244
rect 2596 16192 2648 16244
rect 3056 16192 3108 16244
rect 3424 16192 3476 16244
rect 3608 16192 3660 16244
rect 2320 16124 2372 16176
rect 1308 16056 1360 16108
rect 2504 16099 2556 16108
rect 2504 16065 2513 16099
rect 2513 16065 2547 16099
rect 2547 16065 2556 16099
rect 2504 16056 2556 16065
rect 2596 16099 2648 16108
rect 2596 16065 2605 16099
rect 2605 16065 2639 16099
rect 2639 16065 2648 16099
rect 2596 16056 2648 16065
rect 2688 16056 2740 16108
rect 3516 16056 3568 16108
rect 4252 16056 4304 16108
rect 6000 16124 6052 16176
rect 6092 16124 6144 16176
rect 2412 15920 2464 15972
rect 4068 15988 4120 16040
rect 3424 15920 3476 15972
rect 3884 15920 3936 15972
rect 5448 15852 5500 15904
rect 6736 15852 6788 15904
rect 7104 16235 7156 16244
rect 7104 16201 7113 16235
rect 7113 16201 7147 16235
rect 7147 16201 7156 16235
rect 7104 16192 7156 16201
rect 8208 16192 8260 16244
rect 9864 16235 9916 16244
rect 9864 16201 9873 16235
rect 9873 16201 9907 16235
rect 9907 16201 9916 16235
rect 9864 16192 9916 16201
rect 7196 16167 7248 16176
rect 7196 16133 7205 16167
rect 7205 16133 7239 16167
rect 7239 16133 7248 16167
rect 7196 16124 7248 16133
rect 7288 16124 7340 16176
rect 10140 16124 10192 16176
rect 12072 16235 12124 16244
rect 12072 16201 12081 16235
rect 12081 16201 12115 16235
rect 12115 16201 12124 16235
rect 12072 16192 12124 16201
rect 12532 16192 12584 16244
rect 8852 16099 8904 16108
rect 8852 16065 8861 16099
rect 8861 16065 8895 16099
rect 8895 16065 8904 16099
rect 8852 16056 8904 16065
rect 8944 16099 8996 16108
rect 8944 16065 8954 16099
rect 8954 16065 8988 16099
rect 8988 16065 8996 16099
rect 8944 16056 8996 16065
rect 9588 16056 9640 16108
rect 8300 15920 8352 15972
rect 16028 16192 16080 16244
rect 14556 16124 14608 16176
rect 14740 16124 14792 16176
rect 12532 16031 12584 16040
rect 12532 15997 12541 16031
rect 12541 15997 12575 16031
rect 12575 15997 12584 16031
rect 12532 15988 12584 15997
rect 18696 16056 18748 16108
rect 15016 16031 15068 16040
rect 15016 15997 15025 16031
rect 15025 15997 15059 16031
rect 15059 15997 15068 16031
rect 15016 15988 15068 15997
rect 10600 15852 10652 15904
rect 13544 15895 13596 15904
rect 13544 15861 13553 15895
rect 13553 15861 13587 15895
rect 13587 15861 13596 15895
rect 13544 15852 13596 15861
rect 15200 15852 15252 15904
rect 18788 15895 18840 15904
rect 18788 15861 18797 15895
rect 18797 15861 18831 15895
rect 18831 15861 18840 15895
rect 18788 15852 18840 15861
rect 2918 15750 2970 15802
rect 2982 15750 3034 15802
rect 3046 15750 3098 15802
rect 3110 15750 3162 15802
rect 3174 15750 3226 15802
rect 3238 15750 3290 15802
rect 10918 15750 10970 15802
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 11238 15750 11290 15802
rect 18918 15750 18970 15802
rect 18982 15750 19034 15802
rect 19046 15750 19098 15802
rect 19110 15750 19162 15802
rect 19174 15750 19226 15802
rect 19238 15750 19290 15802
rect 26918 15750 26970 15802
rect 26982 15750 27034 15802
rect 27046 15750 27098 15802
rect 27110 15750 27162 15802
rect 27174 15750 27226 15802
rect 27238 15750 27290 15802
rect 3332 15648 3384 15700
rect 3884 15691 3936 15700
rect 3884 15657 3893 15691
rect 3893 15657 3927 15691
rect 3927 15657 3936 15691
rect 3884 15648 3936 15657
rect 5724 15648 5776 15700
rect 2596 15580 2648 15632
rect 7196 15648 7248 15700
rect 9588 15691 9640 15700
rect 9588 15657 9597 15691
rect 9597 15657 9631 15691
rect 9631 15657 9640 15691
rect 9588 15648 9640 15657
rect 10140 15648 10192 15700
rect 10600 15691 10652 15700
rect 10600 15657 10609 15691
rect 10609 15657 10643 15691
rect 10643 15657 10652 15691
rect 10600 15648 10652 15657
rect 12532 15648 12584 15700
rect 15016 15648 15068 15700
rect 1676 15555 1728 15564
rect 1676 15521 1685 15555
rect 1685 15521 1719 15555
rect 1719 15521 1728 15555
rect 1676 15512 1728 15521
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 2320 15487 2372 15496
rect 2320 15453 2329 15487
rect 2329 15453 2363 15487
rect 2363 15453 2372 15487
rect 2320 15444 2372 15453
rect 2412 15487 2464 15496
rect 2412 15453 2422 15487
rect 2422 15453 2456 15487
rect 2456 15453 2464 15487
rect 2412 15444 2464 15453
rect 2504 15376 2556 15428
rect 2688 15419 2740 15428
rect 2688 15385 2697 15419
rect 2697 15385 2731 15419
rect 2731 15385 2740 15419
rect 2688 15376 2740 15385
rect 1860 15308 1912 15360
rect 3332 15487 3384 15496
rect 3332 15453 3340 15487
rect 3340 15453 3374 15487
rect 3374 15453 3384 15487
rect 3332 15444 3384 15453
rect 5724 15512 5776 15564
rect 6460 15512 6512 15564
rect 7288 15580 7340 15632
rect 8392 15580 8444 15632
rect 8852 15580 8904 15632
rect 8944 15512 8996 15564
rect 14556 15580 14608 15632
rect 15568 15580 15620 15632
rect 3608 15376 3660 15428
rect 6092 15444 6144 15496
rect 5448 15376 5500 15428
rect 6644 15487 6696 15496
rect 6644 15453 6654 15487
rect 6654 15453 6688 15487
rect 6688 15453 6696 15487
rect 6644 15444 6696 15453
rect 9772 15444 9824 15496
rect 13636 15512 13688 15564
rect 14740 15512 14792 15564
rect 15200 15512 15252 15564
rect 17316 15512 17368 15564
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 13084 15487 13136 15496
rect 13084 15453 13093 15487
rect 13093 15453 13127 15487
rect 13127 15453 13136 15487
rect 13084 15444 13136 15453
rect 13544 15444 13596 15496
rect 19340 15444 19392 15496
rect 3332 15308 3384 15360
rect 5908 15308 5960 15360
rect 13268 15308 13320 15360
rect 14372 15351 14424 15360
rect 14372 15317 14381 15351
rect 14381 15317 14415 15351
rect 14415 15317 14424 15351
rect 14372 15308 14424 15317
rect 20720 15308 20772 15360
rect 21364 15308 21416 15360
rect 3658 15206 3710 15258
rect 3722 15206 3774 15258
rect 3786 15206 3838 15258
rect 3850 15206 3902 15258
rect 3914 15206 3966 15258
rect 3978 15206 4030 15258
rect 11658 15206 11710 15258
rect 11722 15206 11774 15258
rect 11786 15206 11838 15258
rect 11850 15206 11902 15258
rect 11914 15206 11966 15258
rect 11978 15206 12030 15258
rect 19658 15206 19710 15258
rect 19722 15206 19774 15258
rect 19786 15206 19838 15258
rect 19850 15206 19902 15258
rect 19914 15206 19966 15258
rect 19978 15206 20030 15258
rect 27658 15206 27710 15258
rect 27722 15206 27774 15258
rect 27786 15206 27838 15258
rect 27850 15206 27902 15258
rect 27914 15206 27966 15258
rect 27978 15206 28030 15258
rect 1400 15104 1452 15156
rect 2320 15104 2372 15156
rect 2412 15036 2464 15088
rect 1308 14968 1360 15020
rect 3516 15104 3568 15156
rect 9220 15104 9272 15156
rect 9680 15104 9732 15156
rect 12624 15104 12676 15156
rect 13084 15147 13136 15156
rect 13084 15113 13093 15147
rect 13093 15113 13127 15147
rect 13127 15113 13136 15147
rect 13084 15104 13136 15113
rect 18788 15104 18840 15156
rect 4436 15036 4488 15088
rect 8024 15036 8076 15088
rect 18420 15036 18472 15088
rect 2964 15011 3016 15020
rect 2964 14977 2973 15011
rect 2973 14977 3007 15011
rect 3007 14977 3016 15011
rect 2964 14968 3016 14977
rect 2504 14900 2556 14952
rect 2596 14900 2648 14952
rect 6644 14968 6696 15020
rect 9588 14968 9640 15020
rect 10048 14968 10100 15020
rect 10416 14968 10468 15020
rect 18788 15011 18840 15020
rect 18788 14977 18797 15011
rect 18797 14977 18831 15011
rect 18831 14977 18840 15011
rect 18788 14968 18840 14977
rect 20720 15036 20772 15088
rect 3700 14943 3752 14952
rect 3700 14909 3709 14943
rect 3709 14909 3743 14943
rect 3743 14909 3752 14943
rect 3700 14900 3752 14909
rect 4068 14900 4120 14952
rect 6000 14900 6052 14952
rect 6184 14900 6236 14952
rect 1860 14832 1912 14884
rect 3240 14832 3292 14884
rect 5724 14832 5776 14884
rect 9772 14900 9824 14952
rect 13268 14900 13320 14952
rect 13360 14943 13412 14952
rect 13360 14909 13369 14943
rect 13369 14909 13403 14943
rect 13403 14909 13412 14943
rect 13360 14900 13412 14909
rect 19616 14968 19668 15020
rect 21180 15011 21232 15020
rect 21180 14977 21189 15011
rect 21189 14977 21223 15011
rect 21223 14977 21232 15011
rect 21180 14968 21232 14977
rect 23480 15036 23532 15088
rect 24216 15036 24268 15088
rect 20628 14900 20680 14952
rect 9864 14832 9916 14884
rect 17960 14764 18012 14816
rect 21916 14764 21968 14816
rect 2918 14662 2970 14714
rect 2982 14662 3034 14714
rect 3046 14662 3098 14714
rect 3110 14662 3162 14714
rect 3174 14662 3226 14714
rect 3238 14662 3290 14714
rect 10918 14662 10970 14714
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 11238 14662 11290 14714
rect 18918 14662 18970 14714
rect 18982 14662 19034 14714
rect 19046 14662 19098 14714
rect 19110 14662 19162 14714
rect 19174 14662 19226 14714
rect 19238 14662 19290 14714
rect 26918 14662 26970 14714
rect 26982 14662 27034 14714
rect 27046 14662 27098 14714
rect 27110 14662 27162 14714
rect 27174 14662 27226 14714
rect 27238 14662 27290 14714
rect 1308 14560 1360 14612
rect 4252 14603 4304 14612
rect 4252 14569 4261 14603
rect 4261 14569 4295 14603
rect 4295 14569 4304 14603
rect 4252 14560 4304 14569
rect 15844 14560 15896 14612
rect 16212 14603 16264 14612
rect 16212 14569 16221 14603
rect 16221 14569 16255 14603
rect 16255 14569 16264 14603
rect 16212 14560 16264 14569
rect 2596 14492 2648 14544
rect 1308 14356 1360 14408
rect 2412 14356 2464 14408
rect 2688 14356 2740 14408
rect 3700 14424 3752 14476
rect 15200 14424 15252 14476
rect 16120 14424 16172 14476
rect 17316 14467 17368 14476
rect 17316 14433 17325 14467
rect 17325 14433 17359 14467
rect 17359 14433 17368 14467
rect 17316 14424 17368 14433
rect 19524 14424 19576 14476
rect 3516 14356 3568 14408
rect 3148 14331 3200 14340
rect 3148 14297 3157 14331
rect 3157 14297 3191 14331
rect 3191 14297 3200 14331
rect 3148 14288 3200 14297
rect 3424 14288 3476 14340
rect 18696 14356 18748 14408
rect 15936 14288 15988 14340
rect 4068 14220 4120 14272
rect 15200 14263 15252 14272
rect 15200 14229 15209 14263
rect 15209 14229 15243 14263
rect 15243 14229 15252 14263
rect 15200 14220 15252 14229
rect 16580 14263 16632 14272
rect 16580 14229 16589 14263
rect 16589 14229 16623 14263
rect 16623 14229 16632 14263
rect 16580 14220 16632 14229
rect 18880 14220 18932 14272
rect 19616 14399 19668 14408
rect 19616 14365 19625 14399
rect 19625 14365 19659 14399
rect 19659 14365 19668 14399
rect 19616 14356 19668 14365
rect 21364 14467 21416 14476
rect 21364 14433 21373 14467
rect 21373 14433 21407 14467
rect 21407 14433 21416 14467
rect 21364 14424 21416 14433
rect 23204 14424 23256 14476
rect 21088 14399 21140 14408
rect 21088 14365 21097 14399
rect 21097 14365 21131 14399
rect 21131 14365 21140 14399
rect 21088 14356 21140 14365
rect 20628 14220 20680 14272
rect 23480 14288 23532 14340
rect 23112 14263 23164 14272
rect 23112 14229 23121 14263
rect 23121 14229 23155 14263
rect 23155 14229 23164 14263
rect 23112 14220 23164 14229
rect 3658 14118 3710 14170
rect 3722 14118 3774 14170
rect 3786 14118 3838 14170
rect 3850 14118 3902 14170
rect 3914 14118 3966 14170
rect 3978 14118 4030 14170
rect 11658 14118 11710 14170
rect 11722 14118 11774 14170
rect 11786 14118 11838 14170
rect 11850 14118 11902 14170
rect 11914 14118 11966 14170
rect 11978 14118 12030 14170
rect 19658 14118 19710 14170
rect 19722 14118 19774 14170
rect 19786 14118 19838 14170
rect 19850 14118 19902 14170
rect 19914 14118 19966 14170
rect 19978 14118 20030 14170
rect 27658 14118 27710 14170
rect 27722 14118 27774 14170
rect 27786 14118 27838 14170
rect 27850 14118 27902 14170
rect 27914 14118 27966 14170
rect 27978 14118 28030 14170
rect 3516 14059 3568 14068
rect 3516 14025 3525 14059
rect 3525 14025 3559 14059
rect 3559 14025 3568 14059
rect 3516 14016 3568 14025
rect 4068 14016 4120 14068
rect 3148 13948 3200 14000
rect 1308 13880 1360 13932
rect 2964 13923 3016 13932
rect 2964 13889 2973 13923
rect 2973 13889 3007 13923
rect 3007 13889 3016 13923
rect 2964 13880 3016 13889
rect 3792 13923 3844 13932
rect 3792 13889 3801 13923
rect 3801 13889 3835 13923
rect 3835 13889 3844 13923
rect 3792 13880 3844 13889
rect 3884 13923 3936 13932
rect 3884 13889 3893 13923
rect 3893 13889 3927 13923
rect 3927 13889 3936 13923
rect 3884 13880 3936 13889
rect 3976 13880 4028 13932
rect 4160 13923 4212 13932
rect 4160 13889 4169 13923
rect 4169 13889 4203 13923
rect 4203 13889 4212 13923
rect 4160 13880 4212 13889
rect 6000 13948 6052 14000
rect 2412 13744 2464 13796
rect 6092 13812 6144 13864
rect 6460 13923 6512 13932
rect 6460 13889 6469 13923
rect 6469 13889 6503 13923
rect 6503 13889 6512 13923
rect 6460 13880 6512 13889
rect 8024 13991 8076 14000
rect 8024 13957 8033 13991
rect 8033 13957 8067 13991
rect 8067 13957 8076 13991
rect 8024 13948 8076 13957
rect 7012 13880 7064 13932
rect 8116 13923 8168 13932
rect 8116 13889 8125 13923
rect 8125 13889 8159 13923
rect 8159 13889 8168 13923
rect 8116 13880 8168 13889
rect 8484 14016 8536 14068
rect 9588 14059 9640 14068
rect 9588 14025 9597 14059
rect 9597 14025 9631 14059
rect 9631 14025 9640 14059
rect 9588 14016 9640 14025
rect 12164 14016 12216 14068
rect 15108 14016 15160 14068
rect 18788 14016 18840 14068
rect 22284 14016 22336 14068
rect 22376 14016 22428 14068
rect 9220 13991 9272 14000
rect 9220 13957 9229 13991
rect 9229 13957 9263 13991
rect 9263 13957 9272 13991
rect 9220 13948 9272 13957
rect 9496 13948 9548 14000
rect 13268 13880 13320 13932
rect 14740 13948 14792 14000
rect 17960 13991 18012 14000
rect 17960 13957 17969 13991
rect 17969 13957 18003 13991
rect 18003 13957 18012 13991
rect 17960 13948 18012 13957
rect 18512 13948 18564 14000
rect 21364 13948 21416 14000
rect 15568 13880 15620 13932
rect 2596 13676 2648 13728
rect 3332 13744 3384 13796
rect 7104 13744 7156 13796
rect 8944 13812 8996 13864
rect 10048 13812 10100 13864
rect 12532 13855 12584 13864
rect 12532 13821 12541 13855
rect 12541 13821 12575 13855
rect 12575 13821 12584 13855
rect 12532 13812 12584 13821
rect 12164 13744 12216 13796
rect 14464 13855 14516 13864
rect 14464 13821 14473 13855
rect 14473 13821 14507 13855
rect 14507 13821 14516 13855
rect 14464 13812 14516 13821
rect 15936 13855 15988 13864
rect 15936 13821 15945 13855
rect 15945 13821 15979 13855
rect 15979 13821 15988 13855
rect 15936 13812 15988 13821
rect 16120 13855 16172 13864
rect 16120 13821 16129 13855
rect 16129 13821 16163 13855
rect 16163 13821 16172 13855
rect 16120 13812 16172 13821
rect 17316 13880 17368 13932
rect 21088 13880 21140 13932
rect 23112 13880 23164 13932
rect 24216 13948 24268 14000
rect 24676 13948 24728 14000
rect 18512 13812 18564 13864
rect 21916 13812 21968 13864
rect 22376 13855 22428 13864
rect 22376 13821 22385 13855
rect 22385 13821 22419 13855
rect 22419 13821 22428 13855
rect 22376 13812 22428 13821
rect 3056 13719 3108 13728
rect 3056 13685 3065 13719
rect 3065 13685 3099 13719
rect 3099 13685 3108 13719
rect 3056 13676 3108 13685
rect 3792 13676 3844 13728
rect 8392 13676 8444 13728
rect 9404 13719 9456 13728
rect 9404 13685 9413 13719
rect 9413 13685 9447 13719
rect 9447 13685 9456 13719
rect 9404 13676 9456 13685
rect 12072 13719 12124 13728
rect 12072 13685 12081 13719
rect 12081 13685 12115 13719
rect 12115 13685 12124 13719
rect 12072 13676 12124 13685
rect 23204 13855 23256 13864
rect 23204 13821 23213 13855
rect 23213 13821 23247 13855
rect 23247 13821 23256 13855
rect 23204 13812 23256 13821
rect 24216 13855 24268 13864
rect 24216 13821 24225 13855
rect 24225 13821 24259 13855
rect 24259 13821 24268 13855
rect 24216 13812 24268 13821
rect 24768 13812 24820 13864
rect 23664 13676 23716 13728
rect 23848 13719 23900 13728
rect 23848 13685 23857 13719
rect 23857 13685 23891 13719
rect 23891 13685 23900 13719
rect 23848 13676 23900 13685
rect 2918 13574 2970 13626
rect 2982 13574 3034 13626
rect 3046 13574 3098 13626
rect 3110 13574 3162 13626
rect 3174 13574 3226 13626
rect 3238 13574 3290 13626
rect 10918 13574 10970 13626
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 11238 13574 11290 13626
rect 18918 13574 18970 13626
rect 18982 13574 19034 13626
rect 19046 13574 19098 13626
rect 19110 13574 19162 13626
rect 19174 13574 19226 13626
rect 19238 13574 19290 13626
rect 26918 13574 26970 13626
rect 26982 13574 27034 13626
rect 27046 13574 27098 13626
rect 27110 13574 27162 13626
rect 27174 13574 27226 13626
rect 27238 13574 27290 13626
rect 3516 13515 3568 13524
rect 3516 13481 3525 13515
rect 3525 13481 3559 13515
rect 3559 13481 3568 13515
rect 3516 13472 3568 13481
rect 4160 13472 4212 13524
rect 6092 13472 6144 13524
rect 6460 13472 6512 13524
rect 7012 13515 7064 13524
rect 7012 13481 7021 13515
rect 7021 13481 7055 13515
rect 7055 13481 7064 13515
rect 7012 13472 7064 13481
rect 2872 13404 2924 13456
rect 3976 13404 4028 13456
rect 8116 13472 8168 13524
rect 8944 13515 8996 13524
rect 8944 13481 8953 13515
rect 8953 13481 8987 13515
rect 8987 13481 8996 13515
rect 8944 13472 8996 13481
rect 14464 13515 14516 13524
rect 14464 13481 14473 13515
rect 14473 13481 14507 13515
rect 14507 13481 14516 13515
rect 14464 13472 14516 13481
rect 24216 13472 24268 13524
rect 2780 13336 2832 13388
rect 3516 13336 3568 13388
rect 4252 13379 4304 13388
rect 4252 13345 4261 13379
rect 4261 13345 4295 13379
rect 4295 13345 4304 13379
rect 4252 13336 4304 13345
rect 6276 13336 6328 13388
rect 1216 13268 1268 13320
rect 2504 13268 2556 13320
rect 3240 13268 3292 13320
rect 3424 13200 3476 13252
rect 4068 13200 4120 13252
rect 4436 13311 4488 13320
rect 4436 13277 4445 13311
rect 4445 13277 4479 13311
rect 4479 13277 4488 13311
rect 4436 13268 4488 13277
rect 6000 13311 6052 13320
rect 6000 13277 6009 13311
rect 6009 13277 6043 13311
rect 6043 13277 6052 13311
rect 6000 13268 6052 13277
rect 6552 13268 6604 13320
rect 8024 13404 8076 13456
rect 14832 13404 14884 13456
rect 6920 13336 6972 13388
rect 7840 13336 7892 13388
rect 4528 13132 4580 13184
rect 6552 13132 6604 13184
rect 8392 13311 8444 13320
rect 8392 13277 8401 13311
rect 8401 13277 8435 13311
rect 8435 13277 8444 13311
rect 8392 13268 8444 13277
rect 9404 13336 9456 13388
rect 24492 13404 24544 13456
rect 23848 13336 23900 13388
rect 8852 13268 8904 13320
rect 9496 13268 9548 13320
rect 9864 13311 9916 13320
rect 9864 13277 9903 13311
rect 9903 13277 9916 13311
rect 9864 13268 9916 13277
rect 10048 13311 10100 13320
rect 10048 13277 10057 13311
rect 10057 13277 10091 13311
rect 10091 13277 10100 13311
rect 10048 13268 10100 13277
rect 11336 13311 11388 13320
rect 11336 13277 11345 13311
rect 11345 13277 11379 13311
rect 11379 13277 11388 13311
rect 11336 13268 11388 13277
rect 15936 13268 15988 13320
rect 24768 13311 24820 13320
rect 24768 13277 24777 13311
rect 24777 13277 24811 13311
rect 24811 13277 24820 13311
rect 24768 13268 24820 13277
rect 7104 13243 7156 13252
rect 7104 13209 7113 13243
rect 7113 13209 7147 13243
rect 7147 13209 7156 13243
rect 7104 13200 7156 13209
rect 11520 13200 11572 13252
rect 13820 13200 13872 13252
rect 7196 13132 7248 13184
rect 9220 13132 9272 13184
rect 13452 13175 13504 13184
rect 13452 13141 13461 13175
rect 13461 13141 13495 13175
rect 13495 13141 13504 13175
rect 13452 13132 13504 13141
rect 3658 13030 3710 13082
rect 3722 13030 3774 13082
rect 3786 13030 3838 13082
rect 3850 13030 3902 13082
rect 3914 13030 3966 13082
rect 3978 13030 4030 13082
rect 11658 13030 11710 13082
rect 11722 13030 11774 13082
rect 11786 13030 11838 13082
rect 11850 13030 11902 13082
rect 11914 13030 11966 13082
rect 11978 13030 12030 13082
rect 19658 13030 19710 13082
rect 19722 13030 19774 13082
rect 19786 13030 19838 13082
rect 19850 13030 19902 13082
rect 19914 13030 19966 13082
rect 19978 13030 20030 13082
rect 27658 13030 27710 13082
rect 27722 13030 27774 13082
rect 27786 13030 27838 13082
rect 27850 13030 27902 13082
rect 27914 13030 27966 13082
rect 27978 13030 28030 13082
rect 1216 12928 1268 12980
rect 2780 12928 2832 12980
rect 3424 12971 3476 12980
rect 3424 12937 3433 12971
rect 3433 12937 3467 12971
rect 3467 12937 3476 12971
rect 3424 12928 3476 12937
rect 3608 12928 3660 12980
rect 6552 12928 6604 12980
rect 7196 12928 7248 12980
rect 9220 12971 9272 12980
rect 9220 12937 9229 12971
rect 9229 12937 9263 12971
rect 9263 12937 9272 12971
rect 9220 12928 9272 12937
rect 11428 12928 11480 12980
rect 4068 12860 4120 12912
rect 8392 12860 8444 12912
rect 1308 12792 1360 12844
rect 2596 12835 2648 12844
rect 2596 12801 2635 12835
rect 2635 12801 2648 12835
rect 2596 12792 2648 12801
rect 2964 12792 3016 12844
rect 3332 12792 3384 12844
rect 6276 12792 6328 12844
rect 8852 12835 8904 12844
rect 8852 12801 8861 12835
rect 8861 12801 8895 12835
rect 8895 12801 8904 12835
rect 8852 12792 8904 12801
rect 12072 12860 12124 12912
rect 12716 12928 12768 12980
rect 13268 12971 13320 12980
rect 13268 12937 13277 12971
rect 13277 12937 13311 12971
rect 13311 12937 13320 12971
rect 13268 12928 13320 12937
rect 14832 12928 14884 12980
rect 15844 12971 15896 12980
rect 15844 12937 15853 12971
rect 15853 12937 15887 12971
rect 15887 12937 15896 12971
rect 15844 12928 15896 12937
rect 18788 12928 18840 12980
rect 15292 12860 15344 12912
rect 16948 12860 17000 12912
rect 18696 12860 18748 12912
rect 11336 12792 11388 12844
rect 13452 12792 13504 12844
rect 13636 12835 13688 12844
rect 13636 12801 13645 12835
rect 13645 12801 13679 12835
rect 13679 12801 13688 12835
rect 13636 12792 13688 12801
rect 2412 12724 2464 12776
rect 3240 12724 3292 12776
rect 3424 12724 3476 12776
rect 6460 12767 6512 12776
rect 6460 12733 6469 12767
rect 6469 12733 6503 12767
rect 6503 12733 6512 12767
rect 6460 12724 6512 12733
rect 18788 12724 18840 12776
rect 19524 12724 19576 12776
rect 20536 12724 20588 12776
rect 21180 12724 21232 12776
rect 2872 12656 2924 12708
rect 2964 12656 3016 12708
rect 3608 12656 3660 12708
rect 2044 12588 2096 12640
rect 6276 12588 6328 12640
rect 11428 12588 11480 12640
rect 16764 12631 16816 12640
rect 16764 12597 16773 12631
rect 16773 12597 16807 12631
rect 16807 12597 16816 12631
rect 16764 12588 16816 12597
rect 18696 12631 18748 12640
rect 18696 12597 18705 12631
rect 18705 12597 18739 12631
rect 18739 12597 18748 12631
rect 18696 12588 18748 12597
rect 22008 12588 22060 12640
rect 2918 12486 2970 12538
rect 2982 12486 3034 12538
rect 3046 12486 3098 12538
rect 3110 12486 3162 12538
rect 3174 12486 3226 12538
rect 3238 12486 3290 12538
rect 10918 12486 10970 12538
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 11238 12486 11290 12538
rect 18918 12486 18970 12538
rect 18982 12486 19034 12538
rect 19046 12486 19098 12538
rect 19110 12486 19162 12538
rect 19174 12486 19226 12538
rect 19238 12486 19290 12538
rect 26918 12486 26970 12538
rect 26982 12486 27034 12538
rect 27046 12486 27098 12538
rect 27110 12486 27162 12538
rect 27174 12486 27226 12538
rect 27238 12486 27290 12538
rect 3332 12384 3384 12436
rect 12532 12384 12584 12436
rect 13636 12384 13688 12436
rect 20812 12384 20864 12436
rect 3608 12316 3660 12368
rect 1952 12291 2004 12300
rect 1952 12257 1961 12291
rect 1961 12257 1995 12291
rect 1995 12257 2004 12291
rect 1952 12248 2004 12257
rect 12532 12248 12584 12300
rect 13820 12316 13872 12368
rect 21916 12359 21968 12368
rect 21916 12325 21925 12359
rect 21925 12325 21959 12359
rect 21959 12325 21968 12359
rect 21916 12316 21968 12325
rect 13360 12248 13412 12300
rect 13728 12248 13780 12300
rect 14740 12248 14792 12300
rect 22008 12248 22060 12300
rect 24492 12316 24544 12368
rect 24676 12359 24728 12368
rect 24676 12325 24685 12359
rect 24685 12325 24719 12359
rect 24719 12325 24728 12359
rect 24676 12316 24728 12325
rect 1308 12180 1360 12232
rect 5724 12180 5776 12232
rect 10692 12180 10744 12232
rect 2596 12155 2648 12164
rect 2596 12121 2605 12155
rect 2605 12121 2639 12155
rect 2639 12121 2648 12155
rect 2596 12112 2648 12121
rect 4160 12087 4212 12096
rect 4160 12053 4169 12087
rect 4169 12053 4203 12087
rect 4203 12053 4212 12087
rect 4160 12044 4212 12053
rect 11152 12044 11204 12096
rect 16764 12223 16816 12232
rect 16764 12189 16773 12223
rect 16773 12189 16807 12223
rect 16807 12189 16816 12223
rect 16764 12180 16816 12189
rect 12532 12112 12584 12164
rect 13636 12112 13688 12164
rect 15292 12112 15344 12164
rect 16212 12112 16264 12164
rect 16488 12112 16540 12164
rect 16948 12112 17000 12164
rect 21824 12112 21876 12164
rect 13268 12044 13320 12096
rect 16672 12087 16724 12096
rect 16672 12053 16681 12087
rect 16681 12053 16715 12087
rect 16715 12053 16724 12087
rect 16672 12044 16724 12053
rect 23296 12044 23348 12096
rect 23572 12087 23624 12096
rect 23572 12053 23581 12087
rect 23581 12053 23615 12087
rect 23615 12053 23624 12087
rect 23572 12044 23624 12053
rect 3658 11942 3710 11994
rect 3722 11942 3774 11994
rect 3786 11942 3838 11994
rect 3850 11942 3902 11994
rect 3914 11942 3966 11994
rect 3978 11942 4030 11994
rect 11658 11942 11710 11994
rect 11722 11942 11774 11994
rect 11786 11942 11838 11994
rect 11850 11942 11902 11994
rect 11914 11942 11966 11994
rect 11978 11942 12030 11994
rect 19658 11942 19710 11994
rect 19722 11942 19774 11994
rect 19786 11942 19838 11994
rect 19850 11942 19902 11994
rect 19914 11942 19966 11994
rect 19978 11942 20030 11994
rect 27658 11942 27710 11994
rect 27722 11942 27774 11994
rect 27786 11942 27838 11994
rect 27850 11942 27902 11994
rect 27914 11942 27966 11994
rect 27978 11942 28030 11994
rect 2412 11883 2464 11892
rect 2412 11849 2421 11883
rect 2421 11849 2455 11883
rect 2455 11849 2464 11883
rect 2412 11840 2464 11849
rect 8852 11840 8904 11892
rect 15292 11883 15344 11892
rect 15292 11849 15301 11883
rect 15301 11849 15335 11883
rect 15335 11849 15344 11883
rect 15292 11840 15344 11849
rect 15568 11840 15620 11892
rect 16212 11883 16264 11892
rect 16212 11849 16221 11883
rect 16221 11849 16255 11883
rect 16255 11849 16264 11883
rect 16212 11840 16264 11849
rect 18696 11840 18748 11892
rect 22284 11883 22336 11892
rect 22284 11849 22293 11883
rect 22293 11849 22327 11883
rect 22327 11849 22336 11883
rect 22284 11840 22336 11849
rect 23572 11840 23624 11892
rect 24768 11883 24820 11892
rect 24768 11849 24777 11883
rect 24777 11849 24811 11883
rect 24811 11849 24820 11883
rect 24768 11840 24820 11849
rect 11428 11772 11480 11824
rect 16672 11772 16724 11824
rect 23296 11815 23348 11824
rect 23296 11781 23305 11815
rect 23305 11781 23339 11815
rect 23339 11781 23348 11815
rect 23296 11772 23348 11781
rect 24584 11772 24636 11824
rect 1952 11747 2004 11756
rect 1952 11713 1961 11747
rect 1961 11713 1995 11747
rect 1995 11713 2004 11747
rect 1952 11704 2004 11713
rect 2320 11747 2372 11756
rect 2320 11713 2329 11747
rect 2329 11713 2363 11747
rect 2363 11713 2372 11747
rect 2320 11704 2372 11713
rect 2780 11704 2832 11756
rect 1308 11636 1360 11688
rect 2688 11636 2740 11688
rect 9404 11679 9456 11688
rect 9404 11645 9413 11679
rect 9413 11645 9447 11679
rect 9447 11645 9456 11679
rect 9404 11636 9456 11645
rect 9680 11679 9732 11688
rect 9680 11645 9689 11679
rect 9689 11645 9723 11679
rect 9723 11645 9732 11679
rect 9680 11636 9732 11645
rect 1032 11568 1084 11620
rect 15016 11704 15068 11756
rect 16120 11704 16172 11756
rect 16488 11704 16540 11756
rect 15752 11679 15804 11688
rect 15752 11645 15761 11679
rect 15761 11645 15795 11679
rect 15795 11645 15804 11679
rect 15752 11636 15804 11645
rect 15844 11636 15896 11688
rect 16672 11679 16724 11688
rect 16672 11645 16681 11679
rect 16681 11645 16715 11679
rect 16715 11645 16724 11679
rect 16672 11636 16724 11645
rect 16948 11747 17000 11756
rect 16948 11713 16957 11747
rect 16957 11713 16991 11747
rect 16991 11713 17000 11747
rect 16948 11704 17000 11713
rect 19432 11704 19484 11756
rect 20720 11704 20772 11756
rect 21916 11636 21968 11688
rect 3332 11500 3384 11552
rect 3608 11500 3660 11552
rect 4252 11500 4304 11552
rect 10784 11500 10836 11552
rect 11152 11543 11204 11552
rect 11152 11509 11161 11543
rect 11161 11509 11195 11543
rect 11195 11509 11204 11543
rect 11152 11500 11204 11509
rect 11428 11500 11480 11552
rect 19340 11568 19392 11620
rect 22008 11568 22060 11620
rect 17592 11500 17644 11552
rect 22100 11500 22152 11552
rect 2918 11398 2970 11450
rect 2982 11398 3034 11450
rect 3046 11398 3098 11450
rect 3110 11398 3162 11450
rect 3174 11398 3226 11450
rect 3238 11398 3290 11450
rect 10918 11398 10970 11450
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 11238 11398 11290 11450
rect 18918 11398 18970 11450
rect 18982 11398 19034 11450
rect 19046 11398 19098 11450
rect 19110 11398 19162 11450
rect 19174 11398 19226 11450
rect 19238 11398 19290 11450
rect 26918 11398 26970 11450
rect 26982 11398 27034 11450
rect 27046 11398 27098 11450
rect 27110 11398 27162 11450
rect 27174 11398 27226 11450
rect 27238 11398 27290 11450
rect 2136 11296 2188 11348
rect 2688 11296 2740 11348
rect 3700 11296 3752 11348
rect 3792 11339 3844 11348
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 3884 11296 3936 11348
rect 2044 11203 2096 11212
rect 2044 11169 2053 11203
rect 2053 11169 2087 11203
rect 2087 11169 2096 11203
rect 2044 11160 2096 11169
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 1584 11092 1636 11144
rect 2320 11092 2372 11144
rect 3516 11092 3568 11144
rect 4344 11228 4396 11280
rect 4160 11160 4212 11212
rect 14372 11296 14424 11348
rect 15752 11296 15804 11348
rect 13728 11228 13780 11280
rect 15016 11203 15068 11212
rect 4252 11135 4304 11144
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 4344 11135 4396 11144
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 4436 11135 4488 11144
rect 4436 11101 4445 11135
rect 4445 11101 4479 11135
rect 4479 11101 4488 11135
rect 4436 11092 4488 11101
rect 4804 11135 4856 11144
rect 4804 11101 4813 11135
rect 4813 11101 4847 11135
rect 4847 11101 4856 11135
rect 4804 11092 4856 11101
rect 9404 11092 9456 11144
rect 11428 11024 11480 11076
rect 14004 11024 14056 11076
rect 15016 11169 15025 11203
rect 15025 11169 15059 11203
rect 15059 11169 15068 11203
rect 15016 11160 15068 11169
rect 15200 11092 15252 11144
rect 17592 11203 17644 11212
rect 17592 11169 17601 11203
rect 17601 11169 17635 11203
rect 17635 11169 17644 11203
rect 17592 11160 17644 11169
rect 15568 11092 15620 11144
rect 16028 11092 16080 11144
rect 16488 11092 16540 11144
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 19432 11296 19484 11348
rect 20628 11228 20680 11280
rect 23480 11228 23532 11280
rect 24584 11228 24636 11280
rect 22008 11160 22060 11212
rect 24768 11160 24820 11212
rect 14280 11067 14332 11076
rect 14280 11033 14289 11067
rect 14289 11033 14323 11067
rect 14323 11033 14332 11067
rect 14280 11024 14332 11033
rect 15384 11024 15436 11076
rect 18052 11024 18104 11076
rect 3516 10999 3568 11008
rect 3516 10965 3525 10999
rect 3525 10965 3559 10999
rect 3559 10965 3568 10999
rect 3516 10956 3568 10965
rect 3884 10956 3936 11008
rect 9404 10999 9456 11008
rect 9404 10965 9413 10999
rect 9413 10965 9447 10999
rect 9447 10965 9456 10999
rect 9404 10956 9456 10965
rect 15292 10956 15344 11008
rect 19524 10999 19576 11008
rect 19524 10965 19533 10999
rect 19533 10965 19567 10999
rect 19567 10965 19576 10999
rect 19524 10956 19576 10965
rect 21640 11024 21692 11076
rect 22100 11067 22152 11076
rect 22100 11033 22109 11067
rect 22109 11033 22143 11067
rect 22143 11033 22152 11067
rect 22100 11024 22152 11033
rect 24676 11024 24728 11076
rect 20720 10956 20772 11008
rect 24400 10999 24452 11008
rect 24400 10965 24409 10999
rect 24409 10965 24443 10999
rect 24443 10965 24452 10999
rect 24400 10956 24452 10965
rect 3658 10854 3710 10906
rect 3722 10854 3774 10906
rect 3786 10854 3838 10906
rect 3850 10854 3902 10906
rect 3914 10854 3966 10906
rect 3978 10854 4030 10906
rect 11658 10854 11710 10906
rect 11722 10854 11774 10906
rect 11786 10854 11838 10906
rect 11850 10854 11902 10906
rect 11914 10854 11966 10906
rect 11978 10854 12030 10906
rect 19658 10854 19710 10906
rect 19722 10854 19774 10906
rect 19786 10854 19838 10906
rect 19850 10854 19902 10906
rect 19914 10854 19966 10906
rect 19978 10854 20030 10906
rect 27658 10854 27710 10906
rect 27722 10854 27774 10906
rect 27786 10854 27838 10906
rect 27850 10854 27902 10906
rect 27914 10854 27966 10906
rect 27978 10854 28030 10906
rect 1400 10752 1452 10804
rect 3516 10752 3568 10804
rect 4804 10752 4856 10804
rect 9680 10795 9732 10804
rect 9680 10761 9689 10795
rect 9689 10761 9723 10795
rect 9723 10761 9732 10795
rect 9680 10752 9732 10761
rect 10784 10752 10836 10804
rect 1308 10616 1360 10668
rect 3332 10659 3384 10668
rect 3332 10625 3342 10659
rect 3342 10625 3376 10659
rect 3376 10625 3384 10659
rect 6920 10684 6972 10736
rect 7288 10684 7340 10736
rect 3332 10616 3384 10625
rect 9588 10684 9640 10736
rect 10692 10684 10744 10736
rect 2780 10548 2832 10600
rect 6368 10591 6420 10600
rect 6368 10557 6377 10591
rect 6377 10557 6411 10591
rect 6411 10557 6420 10591
rect 6368 10548 6420 10557
rect 7104 10548 7156 10600
rect 8944 10591 8996 10600
rect 8944 10557 8953 10591
rect 8953 10557 8987 10591
rect 8987 10557 8996 10591
rect 8944 10548 8996 10557
rect 2228 10480 2280 10532
rect 8116 10455 8168 10464
rect 8116 10421 8125 10455
rect 8125 10421 8159 10455
rect 8159 10421 8168 10455
rect 11336 10616 11388 10668
rect 12440 10684 12492 10736
rect 20628 10752 20680 10804
rect 18052 10684 18104 10736
rect 20720 10684 20772 10736
rect 24768 10684 24820 10736
rect 17960 10616 18012 10668
rect 8116 10412 8168 10421
rect 11796 10591 11848 10600
rect 11796 10557 11805 10591
rect 11805 10557 11839 10591
rect 11839 10557 11848 10591
rect 11796 10548 11848 10557
rect 14096 10591 14148 10600
rect 14096 10557 14105 10591
rect 14105 10557 14139 10591
rect 14139 10557 14148 10591
rect 14096 10548 14148 10557
rect 15292 10548 15344 10600
rect 20812 10548 20864 10600
rect 23664 10548 23716 10600
rect 24216 10548 24268 10600
rect 25044 10616 25096 10668
rect 24676 10548 24728 10600
rect 24492 10480 24544 10532
rect 12164 10412 12216 10464
rect 13268 10455 13320 10464
rect 13268 10421 13277 10455
rect 13277 10421 13311 10455
rect 13311 10421 13320 10455
rect 13268 10412 13320 10421
rect 19892 10412 19944 10464
rect 23388 10455 23440 10464
rect 23388 10421 23397 10455
rect 23397 10421 23431 10455
rect 23431 10421 23440 10455
rect 23388 10412 23440 10421
rect 23664 10412 23716 10464
rect 2918 10310 2970 10362
rect 2982 10310 3034 10362
rect 3046 10310 3098 10362
rect 3110 10310 3162 10362
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 10918 10310 10970 10362
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 11238 10310 11290 10362
rect 18918 10310 18970 10362
rect 18982 10310 19034 10362
rect 19046 10310 19098 10362
rect 19110 10310 19162 10362
rect 19174 10310 19226 10362
rect 19238 10310 19290 10362
rect 26918 10310 26970 10362
rect 26982 10310 27034 10362
rect 27046 10310 27098 10362
rect 27110 10310 27162 10362
rect 27174 10310 27226 10362
rect 27238 10310 27290 10362
rect 2596 10208 2648 10260
rect 7012 10208 7064 10260
rect 7104 10251 7156 10260
rect 7104 10217 7113 10251
rect 7113 10217 7147 10251
rect 7147 10217 7156 10251
rect 7104 10208 7156 10217
rect 11796 10208 11848 10260
rect 14096 10251 14148 10260
rect 14096 10217 14105 10251
rect 14105 10217 14139 10251
rect 14139 10217 14148 10251
rect 14096 10208 14148 10217
rect 6368 10072 6420 10124
rect 1308 10004 1360 10056
rect 7564 10115 7616 10124
rect 7564 10081 7573 10115
rect 7573 10081 7607 10115
rect 7607 10081 7616 10115
rect 7564 10072 7616 10081
rect 7656 10115 7708 10124
rect 7656 10081 7665 10115
rect 7665 10081 7699 10115
rect 7699 10081 7708 10115
rect 7656 10072 7708 10081
rect 10784 10140 10836 10192
rect 13452 10140 13504 10192
rect 12164 10115 12216 10124
rect 12164 10081 12173 10115
rect 12173 10081 12207 10115
rect 12207 10081 12216 10115
rect 12164 10072 12216 10081
rect 17868 10072 17920 10124
rect 19524 10072 19576 10124
rect 19892 10115 19944 10124
rect 19892 10081 19901 10115
rect 19901 10081 19935 10115
rect 19935 10081 19944 10115
rect 19892 10072 19944 10081
rect 24492 10072 24544 10124
rect 9404 10004 9456 10056
rect 13268 10004 13320 10056
rect 15292 10004 15344 10056
rect 6276 9936 6328 9988
rect 7288 9936 7340 9988
rect 8116 9936 8168 9988
rect 6736 9868 6788 9920
rect 8944 9868 8996 9920
rect 12072 9911 12124 9920
rect 12072 9877 12081 9911
rect 12081 9877 12115 9911
rect 12115 9877 12124 9911
rect 12072 9868 12124 9877
rect 18144 9868 18196 9920
rect 19524 9868 19576 9920
rect 3658 9766 3710 9818
rect 3722 9766 3774 9818
rect 3786 9766 3838 9818
rect 3850 9766 3902 9818
rect 3914 9766 3966 9818
rect 3978 9766 4030 9818
rect 11658 9766 11710 9818
rect 11722 9766 11774 9818
rect 11786 9766 11838 9818
rect 11850 9766 11902 9818
rect 11914 9766 11966 9818
rect 11978 9766 12030 9818
rect 19658 9766 19710 9818
rect 19722 9766 19774 9818
rect 19786 9766 19838 9818
rect 19850 9766 19902 9818
rect 19914 9766 19966 9818
rect 19978 9766 20030 9818
rect 27658 9766 27710 9818
rect 27722 9766 27774 9818
rect 27786 9766 27838 9818
rect 27850 9766 27902 9818
rect 27914 9766 27966 9818
rect 27978 9766 28030 9818
rect 1584 9707 1636 9716
rect 1584 9673 1593 9707
rect 1593 9673 1627 9707
rect 1627 9673 1636 9707
rect 1584 9664 1636 9673
rect 7012 9664 7064 9716
rect 12072 9664 12124 9716
rect 18052 9664 18104 9716
rect 6736 9639 6788 9648
rect 6736 9605 6745 9639
rect 6745 9605 6779 9639
rect 6779 9605 6788 9639
rect 6736 9596 6788 9605
rect 18144 9639 18196 9648
rect 18144 9605 18153 9639
rect 18153 9605 18187 9639
rect 18187 9605 18196 9639
rect 18144 9596 18196 9605
rect 19524 9664 19576 9716
rect 23388 9664 23440 9716
rect 23664 9639 23716 9648
rect 23664 9605 23673 9639
rect 23673 9605 23707 9639
rect 23707 9605 23716 9639
rect 23664 9596 23716 9605
rect 25136 9596 25188 9648
rect 1308 9528 1360 9580
rect 5448 9460 5500 9512
rect 7656 9528 7708 9580
rect 11520 9528 11572 9580
rect 15384 9528 15436 9580
rect 15844 9528 15896 9580
rect 17316 9528 17368 9580
rect 22376 9571 22428 9580
rect 22376 9537 22385 9571
rect 22385 9537 22419 9571
rect 22419 9537 22428 9571
rect 22376 9528 22428 9537
rect 6644 9503 6696 9512
rect 6644 9469 6653 9503
rect 6653 9469 6687 9503
rect 6687 9469 6696 9503
rect 6644 9460 6696 9469
rect 7840 9324 7892 9376
rect 11980 9460 12032 9512
rect 12532 9392 12584 9444
rect 14188 9460 14240 9512
rect 22008 9460 22060 9512
rect 22744 9460 22796 9512
rect 14832 9392 14884 9444
rect 21824 9392 21876 9444
rect 25044 9460 25096 9512
rect 14372 9324 14424 9376
rect 22100 9324 22152 9376
rect 2918 9222 2970 9274
rect 2982 9222 3034 9274
rect 3046 9222 3098 9274
rect 3110 9222 3162 9274
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 10918 9222 10970 9274
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 11238 9222 11290 9274
rect 18918 9222 18970 9274
rect 18982 9222 19034 9274
rect 19046 9222 19098 9274
rect 19110 9222 19162 9274
rect 19174 9222 19226 9274
rect 19238 9222 19290 9274
rect 26918 9222 26970 9274
rect 26982 9222 27034 9274
rect 27046 9222 27098 9274
rect 27110 9222 27162 9274
rect 27174 9222 27226 9274
rect 27238 9222 27290 9274
rect 4252 9120 4304 9172
rect 5448 9120 5500 9172
rect 7564 9120 7616 9172
rect 3516 9095 3568 9104
rect 3516 9061 3525 9095
rect 3525 9061 3559 9095
rect 3559 9061 3568 9095
rect 11980 9120 12032 9172
rect 14188 9120 14240 9172
rect 15844 9163 15896 9172
rect 15844 9129 15853 9163
rect 15853 9129 15887 9163
rect 15887 9129 15896 9163
rect 15844 9120 15896 9129
rect 19340 9120 19392 9172
rect 3516 9052 3568 9061
rect 6276 8984 6328 9036
rect 7840 9027 7892 9036
rect 7840 8993 7849 9027
rect 7849 8993 7883 9027
rect 7883 8993 7892 9027
rect 7840 8984 7892 8993
rect 9404 8984 9456 9036
rect 11336 8984 11388 9036
rect 11980 9027 12032 9036
rect 11980 8993 11989 9027
rect 11989 8993 12023 9027
rect 12023 8993 12032 9027
rect 11980 8984 12032 8993
rect 14372 9027 14424 9036
rect 14372 8993 14381 9027
rect 14381 8993 14415 9027
rect 14415 8993 14424 9027
rect 14372 8984 14424 8993
rect 1584 8916 1636 8968
rect 3148 8916 3200 8968
rect 3424 8916 3476 8968
rect 11244 8916 11296 8968
rect 12440 8916 12492 8968
rect 14096 8959 14148 8968
rect 14096 8925 14105 8959
rect 14105 8925 14139 8959
rect 14139 8925 14148 8959
rect 14096 8916 14148 8925
rect 21272 8916 21324 8968
rect 2044 8891 2096 8900
rect 2044 8857 2053 8891
rect 2053 8857 2087 8891
rect 2087 8857 2096 8891
rect 2044 8848 2096 8857
rect 4712 8848 4764 8900
rect 1308 8780 1360 8832
rect 4344 8823 4396 8832
rect 4344 8789 4353 8823
rect 4353 8789 4387 8823
rect 4387 8789 4396 8823
rect 4344 8780 4396 8789
rect 6092 8780 6144 8832
rect 7656 8823 7708 8832
rect 7656 8789 7665 8823
rect 7665 8789 7699 8823
rect 7699 8789 7708 8823
rect 7656 8780 7708 8789
rect 7748 8823 7800 8832
rect 7748 8789 7757 8823
rect 7757 8789 7791 8823
rect 7791 8789 7800 8823
rect 7748 8780 7800 8789
rect 10232 8848 10284 8900
rect 11060 8780 11112 8832
rect 11520 8780 11572 8832
rect 15384 8848 15436 8900
rect 21824 8780 21876 8832
rect 23388 8780 23440 8832
rect 3658 8678 3710 8730
rect 3722 8678 3774 8730
rect 3786 8678 3838 8730
rect 3850 8678 3902 8730
rect 3914 8678 3966 8730
rect 3978 8678 4030 8730
rect 11658 8678 11710 8730
rect 11722 8678 11774 8730
rect 11786 8678 11838 8730
rect 11850 8678 11902 8730
rect 11914 8678 11966 8730
rect 11978 8678 12030 8730
rect 19658 8678 19710 8730
rect 19722 8678 19774 8730
rect 19786 8678 19838 8730
rect 19850 8678 19902 8730
rect 19914 8678 19966 8730
rect 19978 8678 20030 8730
rect 27658 8678 27710 8730
rect 27722 8678 27774 8730
rect 27786 8678 27838 8730
rect 27850 8678 27902 8730
rect 27914 8678 27966 8730
rect 27978 8678 28030 8730
rect 2044 8576 2096 8628
rect 3516 8576 3568 8628
rect 6644 8576 6696 8628
rect 7748 8576 7800 8628
rect 10232 8619 10284 8628
rect 10232 8585 10241 8619
rect 10241 8585 10275 8619
rect 10275 8585 10284 8619
rect 10232 8576 10284 8585
rect 11520 8576 11572 8628
rect 17316 8576 17368 8628
rect 24400 8576 24452 8628
rect 7656 8508 7708 8560
rect 19432 8508 19484 8560
rect 22100 8551 22152 8560
rect 22100 8517 22109 8551
rect 22109 8517 22143 8551
rect 22143 8517 22152 8551
rect 22100 8508 22152 8517
rect 23388 8508 23440 8560
rect 25136 8508 25188 8560
rect 1308 8440 1360 8492
rect 3700 8440 3752 8492
rect 3792 8483 3844 8492
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 3884 8483 3936 8492
rect 3884 8449 3893 8483
rect 3893 8449 3927 8483
rect 3927 8449 3936 8483
rect 3884 8440 3936 8449
rect 4160 8440 4212 8492
rect 2780 8372 2832 8424
rect 3148 8304 3200 8356
rect 4252 8304 4304 8356
rect 7196 8372 7248 8424
rect 11336 8440 11388 8492
rect 18052 8440 18104 8492
rect 24768 8440 24820 8492
rect 6920 8304 6972 8356
rect 11060 8372 11112 8424
rect 12164 8372 12216 8424
rect 18788 8372 18840 8424
rect 21824 8415 21876 8424
rect 21824 8381 21833 8415
rect 21833 8381 21867 8415
rect 21867 8381 21876 8415
rect 21824 8372 21876 8381
rect 24492 8372 24544 8424
rect 19524 8304 19576 8356
rect 23388 8304 23440 8356
rect 2780 8236 2832 8288
rect 14556 8236 14608 8288
rect 16764 8236 16816 8288
rect 24676 8236 24728 8288
rect 2918 8134 2970 8186
rect 2982 8134 3034 8186
rect 3046 8134 3098 8186
rect 3110 8134 3162 8186
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 10918 8134 10970 8186
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 11238 8134 11290 8186
rect 18918 8134 18970 8186
rect 18982 8134 19034 8186
rect 19046 8134 19098 8186
rect 19110 8134 19162 8186
rect 19174 8134 19226 8186
rect 19238 8134 19290 8186
rect 26918 8134 26970 8186
rect 26982 8134 27034 8186
rect 27046 8134 27098 8186
rect 27110 8134 27162 8186
rect 27174 8134 27226 8186
rect 27238 8134 27290 8186
rect 3700 8032 3752 8084
rect 7748 8032 7800 8084
rect 4160 7964 4212 8016
rect 1308 7896 1360 7948
rect 4436 7964 4488 8016
rect 4344 7939 4396 7948
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 7104 7896 7156 7948
rect 1216 7828 1268 7880
rect 4068 7828 4120 7880
rect 18052 8032 18104 8084
rect 19340 8075 19392 8084
rect 19340 8041 19349 8075
rect 19349 8041 19383 8075
rect 19383 8041 19392 8075
rect 19340 8032 19392 8041
rect 19524 8075 19576 8084
rect 19524 8041 19533 8075
rect 19533 8041 19567 8075
rect 19567 8041 19576 8075
rect 19524 8032 19576 8041
rect 20444 8032 20496 8084
rect 17868 7964 17920 8016
rect 19892 7964 19944 8016
rect 17316 7939 17368 7948
rect 17316 7905 17325 7939
rect 17325 7905 17359 7939
rect 17359 7905 17368 7939
rect 17316 7896 17368 7905
rect 3516 7760 3568 7812
rect 3792 7760 3844 7812
rect 3884 7692 3936 7744
rect 4160 7735 4212 7744
rect 4160 7701 4169 7735
rect 4169 7701 4203 7735
rect 4203 7701 4212 7735
rect 4160 7692 4212 7701
rect 17960 7828 18012 7880
rect 18696 7896 18748 7948
rect 20076 7939 20128 7948
rect 20076 7905 20085 7939
rect 20085 7905 20119 7939
rect 20119 7905 20128 7939
rect 20076 7896 20128 7905
rect 20536 7964 20588 8016
rect 24676 7939 24728 7948
rect 24676 7905 24685 7939
rect 24685 7905 24719 7939
rect 24719 7905 24728 7939
rect 24676 7896 24728 7905
rect 19616 7828 19668 7880
rect 21824 7828 21876 7880
rect 24400 7871 24452 7880
rect 24400 7837 24409 7871
rect 24409 7837 24443 7871
rect 24443 7837 24452 7871
rect 24400 7828 24452 7837
rect 6736 7803 6788 7812
rect 6736 7769 6745 7803
rect 6745 7769 6779 7803
rect 6779 7769 6788 7803
rect 6736 7760 6788 7769
rect 7288 7760 7340 7812
rect 17040 7803 17092 7812
rect 17040 7769 17049 7803
rect 17049 7769 17083 7803
rect 17083 7769 17092 7803
rect 17040 7760 17092 7769
rect 17500 7803 17552 7812
rect 17500 7769 17509 7803
rect 17509 7769 17543 7803
rect 17543 7769 17552 7803
rect 17500 7760 17552 7769
rect 6920 7692 6972 7744
rect 16948 7692 17000 7744
rect 18788 7692 18840 7744
rect 19524 7692 19576 7744
rect 22376 7760 22428 7812
rect 23388 7760 23440 7812
rect 25136 7760 25188 7812
rect 28356 7803 28408 7812
rect 28356 7769 28365 7803
rect 28365 7769 28399 7803
rect 28399 7769 28408 7803
rect 28356 7760 28408 7769
rect 21272 7692 21324 7744
rect 22284 7692 22336 7744
rect 24768 7692 24820 7744
rect 3658 7590 3710 7642
rect 3722 7590 3774 7642
rect 3786 7590 3838 7642
rect 3850 7590 3902 7642
rect 3914 7590 3966 7642
rect 3978 7590 4030 7642
rect 11658 7590 11710 7642
rect 11722 7590 11774 7642
rect 11786 7590 11838 7642
rect 11850 7590 11902 7642
rect 11914 7590 11966 7642
rect 11978 7590 12030 7642
rect 19658 7590 19710 7642
rect 19722 7590 19774 7642
rect 19786 7590 19838 7642
rect 19850 7590 19902 7642
rect 19914 7590 19966 7642
rect 19978 7590 20030 7642
rect 27658 7590 27710 7642
rect 27722 7590 27774 7642
rect 27786 7590 27838 7642
rect 27850 7590 27902 7642
rect 27914 7590 27966 7642
rect 27978 7590 28030 7642
rect 1308 7488 1360 7540
rect 1584 7488 1636 7540
rect 3332 7488 3384 7540
rect 4068 7488 4120 7540
rect 2596 7420 2648 7472
rect 3608 7420 3660 7472
rect 1584 7395 1636 7404
rect 1584 7361 1593 7395
rect 1593 7361 1627 7395
rect 1627 7361 1636 7395
rect 1584 7352 1636 7361
rect 3516 7352 3568 7404
rect 6736 7488 6788 7540
rect 7748 7488 7800 7540
rect 8852 7531 8904 7540
rect 8852 7497 8861 7531
rect 8861 7497 8895 7531
rect 8895 7497 8904 7531
rect 8852 7488 8904 7497
rect 5632 7420 5684 7472
rect 14832 7463 14884 7472
rect 14832 7429 14841 7463
rect 14841 7429 14875 7463
rect 14875 7429 14884 7463
rect 14832 7420 14884 7429
rect 15384 7531 15436 7540
rect 15384 7497 15393 7531
rect 15393 7497 15427 7531
rect 15427 7497 15436 7531
rect 15384 7488 15436 7497
rect 17040 7488 17092 7540
rect 18788 7488 18840 7540
rect 24768 7488 24820 7540
rect 17500 7420 17552 7472
rect 21640 7420 21692 7472
rect 14556 7395 14608 7404
rect 4620 7327 4672 7336
rect 4620 7293 4629 7327
rect 4629 7293 4663 7327
rect 4663 7293 4672 7327
rect 4620 7284 4672 7293
rect 7656 7327 7708 7336
rect 7656 7293 7665 7327
rect 7665 7293 7699 7327
rect 7699 7293 7708 7327
rect 7656 7284 7708 7293
rect 7840 7327 7892 7336
rect 7840 7293 7849 7327
rect 7849 7293 7883 7327
rect 7883 7293 7892 7327
rect 7840 7284 7892 7293
rect 6000 7148 6052 7200
rect 6092 7191 6144 7200
rect 6092 7157 6101 7191
rect 6101 7157 6135 7191
rect 6135 7157 6144 7191
rect 6092 7148 6144 7157
rect 14188 7148 14240 7200
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 15568 7395 15620 7404
rect 15568 7361 15577 7395
rect 15577 7361 15611 7395
rect 15611 7361 15620 7395
rect 15568 7352 15620 7361
rect 16948 7352 17000 7404
rect 19616 7352 19668 7404
rect 25044 7488 25096 7540
rect 17868 7284 17920 7336
rect 18696 7284 18748 7336
rect 21364 7284 21416 7336
rect 21824 7327 21876 7336
rect 21824 7293 21833 7327
rect 21833 7293 21867 7327
rect 21867 7293 21876 7327
rect 21824 7284 21876 7293
rect 22100 7327 22152 7336
rect 22100 7293 22109 7327
rect 22109 7293 22143 7327
rect 22143 7293 22152 7327
rect 22100 7284 22152 7293
rect 24216 7327 24268 7336
rect 24216 7293 24225 7327
rect 24225 7293 24259 7327
rect 24259 7293 24268 7327
rect 24216 7284 24268 7293
rect 24584 7284 24636 7336
rect 24768 7284 24820 7336
rect 17960 7216 18012 7268
rect 22560 7148 22612 7200
rect 23664 7191 23716 7200
rect 23664 7157 23673 7191
rect 23673 7157 23707 7191
rect 23707 7157 23716 7191
rect 23664 7148 23716 7157
rect 24676 7148 24728 7200
rect 2918 7046 2970 7098
rect 2982 7046 3034 7098
rect 3046 7046 3098 7098
rect 3110 7046 3162 7098
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 10918 7046 10970 7098
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 11238 7046 11290 7098
rect 18918 7046 18970 7098
rect 18982 7046 19034 7098
rect 19046 7046 19098 7098
rect 19110 7046 19162 7098
rect 19174 7046 19226 7098
rect 19238 7046 19290 7098
rect 26918 7046 26970 7098
rect 26982 7046 27034 7098
rect 27046 7046 27098 7098
rect 27110 7046 27162 7098
rect 27174 7046 27226 7098
rect 27238 7046 27290 7098
rect 4620 6944 4672 6996
rect 22100 6944 22152 6996
rect 2688 6876 2740 6928
rect 2780 6876 2832 6928
rect 3424 6808 3476 6860
rect 5448 6851 5500 6860
rect 5448 6817 5457 6851
rect 5457 6817 5491 6851
rect 5491 6817 5500 6851
rect 5448 6808 5500 6817
rect 6920 6808 6972 6860
rect 1308 6740 1360 6792
rect 6092 6740 6144 6792
rect 13820 6808 13872 6860
rect 14096 6851 14148 6860
rect 14096 6817 14105 6851
rect 14105 6817 14139 6851
rect 14139 6817 14148 6851
rect 14096 6808 14148 6817
rect 19524 6808 19576 6860
rect 11336 6740 11388 6792
rect 19340 6740 19392 6792
rect 20536 6808 20588 6860
rect 22008 6808 22060 6860
rect 22744 6851 22796 6860
rect 22744 6817 22753 6851
rect 22753 6817 22787 6851
rect 22787 6817 22796 6851
rect 22744 6808 22796 6817
rect 22560 6783 22612 6792
rect 22560 6749 22569 6783
rect 22569 6749 22603 6783
rect 22603 6749 22612 6783
rect 22560 6740 22612 6749
rect 23664 6740 23716 6792
rect 1216 6672 1268 6724
rect 3424 6672 3476 6724
rect 8760 6715 8812 6724
rect 8760 6681 8769 6715
rect 8769 6681 8803 6715
rect 8803 6681 8812 6715
rect 8760 6672 8812 6681
rect 8852 6672 8904 6724
rect 10324 6672 10376 6724
rect 11520 6672 11572 6724
rect 12808 6715 12860 6724
rect 12808 6681 12817 6715
rect 12817 6681 12851 6715
rect 12851 6681 12860 6715
rect 12808 6672 12860 6681
rect 13728 6715 13780 6724
rect 13728 6681 13737 6715
rect 13737 6681 13771 6715
rect 13771 6681 13780 6715
rect 13728 6672 13780 6681
rect 14372 6715 14424 6724
rect 14372 6681 14381 6715
rect 14381 6681 14415 6715
rect 14415 6681 14424 6715
rect 14372 6672 14424 6681
rect 15384 6672 15436 6724
rect 19616 6715 19668 6724
rect 19616 6681 19625 6715
rect 19625 6681 19659 6715
rect 19659 6681 19668 6715
rect 19616 6672 19668 6681
rect 5540 6604 5592 6656
rect 8024 6604 8076 6656
rect 11336 6647 11388 6656
rect 11336 6613 11345 6647
rect 11345 6613 11379 6647
rect 11379 6613 11388 6647
rect 11336 6604 11388 6613
rect 14096 6604 14148 6656
rect 14740 6604 14792 6656
rect 18512 6604 18564 6656
rect 3658 6502 3710 6554
rect 3722 6502 3774 6554
rect 3786 6502 3838 6554
rect 3850 6502 3902 6554
rect 3914 6502 3966 6554
rect 3978 6502 4030 6554
rect 11658 6502 11710 6554
rect 11722 6502 11774 6554
rect 11786 6502 11838 6554
rect 11850 6502 11902 6554
rect 11914 6502 11966 6554
rect 11978 6502 12030 6554
rect 19658 6502 19710 6554
rect 19722 6502 19774 6554
rect 19786 6502 19838 6554
rect 19850 6502 19902 6554
rect 19914 6502 19966 6554
rect 19978 6502 20030 6554
rect 27658 6502 27710 6554
rect 27722 6502 27774 6554
rect 27786 6502 27838 6554
rect 27850 6502 27902 6554
rect 27914 6502 27966 6554
rect 27978 6502 28030 6554
rect 7656 6400 7708 6452
rect 8760 6400 8812 6452
rect 11428 6400 11480 6452
rect 6920 6332 6972 6384
rect 7196 6332 7248 6384
rect 8116 6332 8168 6384
rect 9588 6332 9640 6384
rect 14372 6443 14424 6452
rect 14372 6409 14381 6443
rect 14381 6409 14415 6443
rect 14415 6409 14424 6443
rect 14372 6400 14424 6409
rect 14740 6443 14792 6452
rect 14740 6409 14749 6443
rect 14749 6409 14783 6443
rect 14783 6409 14792 6443
rect 14740 6400 14792 6409
rect 16948 6400 17000 6452
rect 20904 6400 20956 6452
rect 21640 6400 21692 6452
rect 1308 6264 1360 6316
rect 8208 6307 8260 6316
rect 8208 6273 8217 6307
rect 8217 6273 8251 6307
rect 8251 6273 8260 6307
rect 8208 6264 8260 6273
rect 3608 6196 3660 6248
rect 6184 6128 6236 6180
rect 3700 6103 3752 6112
rect 3700 6069 3709 6103
rect 3709 6069 3743 6103
rect 3743 6069 3752 6103
rect 3700 6060 3752 6069
rect 8024 6196 8076 6248
rect 10692 6264 10744 6316
rect 7104 6128 7156 6180
rect 8852 6060 8904 6112
rect 9772 6239 9824 6248
rect 9772 6205 9781 6239
rect 9781 6205 9815 6239
rect 9815 6205 9824 6239
rect 9772 6196 9824 6205
rect 10324 6171 10376 6180
rect 10324 6137 10333 6171
rect 10333 6137 10367 6171
rect 10367 6137 10376 6171
rect 10324 6128 10376 6137
rect 13820 6264 13872 6316
rect 13912 6307 13964 6316
rect 13912 6273 13921 6307
rect 13921 6273 13955 6307
rect 13955 6273 13964 6307
rect 13912 6264 13964 6273
rect 14096 6264 14148 6316
rect 13728 6196 13780 6248
rect 14832 6196 14884 6248
rect 11336 6128 11388 6180
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 17040 6264 17092 6273
rect 21272 6375 21324 6384
rect 21272 6341 21281 6375
rect 21281 6341 21315 6375
rect 21315 6341 21324 6375
rect 21272 6332 21324 6341
rect 18696 6196 18748 6248
rect 10784 6060 10836 6112
rect 12716 6060 12768 6112
rect 16672 6060 16724 6112
rect 2918 5958 2970 6010
rect 2982 5958 3034 6010
rect 3046 5958 3098 6010
rect 3110 5958 3162 6010
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 10918 5958 10970 6010
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 11238 5958 11290 6010
rect 18918 5958 18970 6010
rect 18982 5958 19034 6010
rect 19046 5958 19098 6010
rect 19110 5958 19162 6010
rect 19174 5958 19226 6010
rect 19238 5958 19290 6010
rect 26918 5958 26970 6010
rect 26982 5958 27034 6010
rect 27046 5958 27098 6010
rect 27110 5958 27162 6010
rect 27174 5958 27226 6010
rect 27238 5958 27290 6010
rect 3056 5856 3108 5908
rect 3608 5856 3660 5908
rect 5540 5899 5592 5908
rect 5540 5865 5549 5899
rect 5549 5865 5583 5899
rect 5583 5865 5592 5899
rect 5540 5856 5592 5865
rect 6000 5856 6052 5908
rect 9772 5856 9824 5908
rect 12164 5899 12216 5908
rect 12164 5865 12173 5899
rect 12173 5865 12207 5899
rect 12207 5865 12216 5899
rect 12164 5856 12216 5865
rect 12808 5856 12860 5908
rect 17960 5856 18012 5908
rect 1308 5652 1360 5704
rect 2504 5695 2556 5704
rect 2504 5661 2513 5695
rect 2513 5661 2547 5695
rect 2547 5661 2556 5695
rect 2504 5652 2556 5661
rect 6092 5788 6144 5840
rect 5724 5720 5776 5772
rect 11612 5788 11664 5840
rect 3700 5652 3752 5704
rect 8024 5763 8076 5772
rect 8024 5729 8033 5763
rect 8033 5729 8067 5763
rect 8067 5729 8076 5763
rect 8024 5720 8076 5729
rect 8116 5763 8168 5772
rect 8116 5729 8125 5763
rect 8125 5729 8159 5763
rect 8159 5729 8168 5763
rect 8116 5720 8168 5729
rect 10784 5763 10836 5772
rect 10784 5729 10793 5763
rect 10793 5729 10827 5763
rect 10827 5729 10836 5763
rect 10784 5720 10836 5729
rect 14096 5831 14148 5840
rect 14096 5797 14105 5831
rect 14105 5797 14139 5831
rect 14139 5797 14148 5831
rect 14096 5788 14148 5797
rect 14740 5788 14792 5840
rect 14832 5788 14884 5840
rect 17224 5788 17276 5840
rect 16672 5763 16724 5772
rect 16672 5729 16681 5763
rect 16681 5729 16715 5763
rect 16715 5729 16724 5763
rect 16672 5720 16724 5729
rect 8208 5652 8260 5704
rect 11336 5695 11388 5704
rect 11336 5661 11345 5695
rect 11345 5661 11379 5695
rect 11379 5661 11388 5695
rect 11336 5652 11388 5661
rect 12716 5695 12768 5704
rect 12716 5661 12725 5695
rect 12725 5661 12759 5695
rect 12759 5661 12768 5695
rect 12716 5652 12768 5661
rect 13912 5652 13964 5704
rect 16948 5652 17000 5704
rect 18512 5763 18564 5772
rect 18512 5729 18521 5763
rect 18521 5729 18555 5763
rect 18555 5729 18564 5763
rect 18512 5720 18564 5729
rect 21364 5720 21416 5772
rect 19340 5652 19392 5704
rect 3240 5516 3292 5568
rect 4988 5516 5040 5568
rect 5172 5559 5224 5568
rect 5172 5525 5181 5559
rect 5181 5525 5215 5559
rect 5215 5525 5224 5559
rect 5172 5516 5224 5525
rect 5724 5559 5776 5568
rect 5724 5525 5733 5559
rect 5733 5525 5767 5559
rect 5767 5525 5776 5559
rect 5724 5516 5776 5525
rect 6092 5584 6144 5636
rect 14188 5584 14240 5636
rect 17040 5584 17092 5636
rect 9772 5516 9824 5568
rect 10876 5559 10928 5568
rect 10876 5525 10885 5559
rect 10885 5525 10919 5559
rect 10919 5525 10928 5559
rect 10876 5516 10928 5525
rect 10968 5516 11020 5568
rect 11336 5516 11388 5568
rect 11612 5516 11664 5568
rect 15568 5516 15620 5568
rect 16028 5559 16080 5568
rect 16028 5525 16037 5559
rect 16037 5525 16071 5559
rect 16071 5525 16080 5559
rect 16028 5516 16080 5525
rect 17960 5516 18012 5568
rect 18420 5559 18472 5568
rect 18420 5525 18429 5559
rect 18429 5525 18463 5559
rect 18463 5525 18472 5559
rect 18420 5516 18472 5525
rect 20904 5584 20956 5636
rect 21456 5584 21508 5636
rect 22008 5627 22060 5636
rect 22008 5593 22017 5627
rect 22017 5593 22051 5627
rect 22051 5593 22060 5627
rect 22008 5584 22060 5593
rect 21180 5516 21232 5568
rect 3658 5414 3710 5466
rect 3722 5414 3774 5466
rect 3786 5414 3838 5466
rect 3850 5414 3902 5466
rect 3914 5414 3966 5466
rect 3978 5414 4030 5466
rect 11658 5414 11710 5466
rect 11722 5414 11774 5466
rect 11786 5414 11838 5466
rect 11850 5414 11902 5466
rect 11914 5414 11966 5466
rect 11978 5414 12030 5466
rect 19658 5414 19710 5466
rect 19722 5414 19774 5466
rect 19786 5414 19838 5466
rect 19850 5414 19902 5466
rect 19914 5414 19966 5466
rect 19978 5414 20030 5466
rect 27658 5414 27710 5466
rect 27722 5414 27774 5466
rect 27786 5414 27838 5466
rect 27850 5414 27902 5466
rect 27914 5414 27966 5466
rect 27978 5414 28030 5466
rect 2504 5312 2556 5364
rect 2688 5312 2740 5364
rect 3700 5355 3752 5364
rect 3700 5321 3709 5355
rect 3709 5321 3743 5355
rect 3743 5321 3752 5355
rect 3700 5312 3752 5321
rect 1308 5176 1360 5228
rect 2596 5040 2648 5092
rect 2780 5040 2832 5092
rect 3056 5219 3108 5228
rect 3056 5185 3065 5219
rect 3065 5185 3099 5219
rect 3099 5185 3108 5219
rect 3056 5176 3108 5185
rect 3240 5176 3292 5228
rect 4712 5244 4764 5296
rect 4252 5176 4304 5228
rect 3516 5108 3568 5160
rect 10876 5312 10928 5364
rect 15384 5312 15436 5364
rect 6184 5287 6236 5296
rect 4988 5176 5040 5228
rect 6184 5253 6193 5287
rect 6193 5253 6227 5287
rect 6227 5253 6236 5287
rect 6184 5244 6236 5253
rect 5356 5151 5408 5160
rect 3424 5040 3476 5092
rect 5356 5117 5365 5151
rect 5365 5117 5399 5151
rect 5399 5117 5408 5151
rect 5356 5108 5408 5117
rect 14004 5244 14056 5296
rect 17960 5244 18012 5296
rect 18420 5312 18472 5364
rect 21180 5355 21232 5364
rect 21180 5321 21189 5355
rect 21189 5321 21223 5355
rect 21223 5321 21232 5355
rect 21180 5312 21232 5321
rect 21456 5312 21508 5364
rect 24400 5312 24452 5364
rect 20904 5244 20956 5296
rect 21824 5244 21876 5296
rect 17316 5176 17368 5228
rect 20720 5108 20772 5160
rect 21916 5108 21968 5160
rect 25136 5108 25188 5160
rect 3056 4972 3108 5024
rect 3608 4972 3660 5024
rect 4620 4972 4672 5024
rect 4712 5015 4764 5024
rect 4712 4981 4721 5015
rect 4721 4981 4755 5015
rect 4755 4981 4764 5015
rect 4712 4972 4764 4981
rect 5724 5015 5776 5024
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 6828 4972 6880 5024
rect 8300 4972 8352 5024
rect 23296 5015 23348 5024
rect 23296 4981 23305 5015
rect 23305 4981 23339 5015
rect 23339 4981 23348 5015
rect 23296 4972 23348 4981
rect 2918 4870 2970 4922
rect 2982 4870 3034 4922
rect 3046 4870 3098 4922
rect 3110 4870 3162 4922
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 10918 4870 10970 4922
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 11238 4870 11290 4922
rect 18918 4870 18970 4922
rect 18982 4870 19034 4922
rect 19046 4870 19098 4922
rect 19110 4870 19162 4922
rect 19174 4870 19226 4922
rect 19238 4870 19290 4922
rect 26918 4870 26970 4922
rect 26982 4870 27034 4922
rect 27046 4870 27098 4922
rect 27110 4870 27162 4922
rect 27174 4870 27226 4922
rect 27238 4870 27290 4922
rect 2964 4768 3016 4820
rect 4068 4768 4120 4820
rect 4252 4768 4304 4820
rect 3516 4743 3568 4752
rect 3516 4709 3525 4743
rect 3525 4709 3559 4743
rect 3559 4709 3568 4743
rect 3516 4700 3568 4709
rect 3332 4632 3384 4684
rect 4712 4632 4764 4684
rect 6920 4675 6972 4684
rect 6920 4641 6929 4675
rect 6929 4641 6963 4675
rect 6963 4641 6972 4675
rect 6920 4632 6972 4641
rect 8208 4768 8260 4820
rect 12532 4768 12584 4820
rect 9680 4632 9732 4684
rect 11520 4632 11572 4684
rect 14832 4675 14884 4684
rect 14832 4641 14841 4675
rect 14841 4641 14875 4675
rect 14875 4641 14884 4675
rect 14832 4632 14884 4641
rect 2780 4564 2832 4616
rect 3608 4564 3660 4616
rect 16028 4564 16080 4616
rect 18512 4811 18564 4820
rect 18512 4777 18521 4811
rect 18521 4777 18555 4811
rect 18555 4777 18564 4811
rect 18512 4768 18564 4777
rect 21916 4811 21968 4820
rect 21916 4777 21925 4811
rect 21925 4777 21959 4811
rect 21959 4777 21968 4811
rect 21916 4768 21968 4777
rect 25136 4811 25188 4820
rect 25136 4777 25145 4811
rect 25145 4777 25179 4811
rect 25179 4777 25188 4811
rect 25136 4768 25188 4777
rect 22008 4700 22060 4752
rect 18512 4632 18564 4684
rect 24216 4632 24268 4684
rect 24676 4675 24728 4684
rect 24676 4641 24685 4675
rect 24685 4641 24719 4675
rect 24719 4641 24728 4675
rect 24676 4632 24728 4641
rect 23296 4564 23348 4616
rect 1676 4539 1728 4548
rect 1676 4505 1685 4539
rect 1685 4505 1719 4539
rect 1719 4505 1728 4539
rect 1676 4496 1728 4505
rect 7196 4539 7248 4548
rect 7196 4505 7205 4539
rect 7205 4505 7239 4539
rect 7239 4505 7248 4539
rect 7196 4496 7248 4505
rect 5448 4428 5500 4480
rect 5632 4428 5684 4480
rect 13912 4496 13964 4548
rect 14372 4428 14424 4480
rect 14740 4428 14792 4480
rect 17868 4496 17920 4548
rect 15660 4428 15712 4480
rect 22376 4471 22428 4480
rect 22376 4437 22385 4471
rect 22385 4437 22419 4471
rect 22419 4437 22428 4471
rect 22376 4428 22428 4437
rect 3658 4326 3710 4378
rect 3722 4326 3774 4378
rect 3786 4326 3838 4378
rect 3850 4326 3902 4378
rect 3914 4326 3966 4378
rect 3978 4326 4030 4378
rect 11658 4326 11710 4378
rect 11722 4326 11774 4378
rect 11786 4326 11838 4378
rect 11850 4326 11902 4378
rect 11914 4326 11966 4378
rect 11978 4326 12030 4378
rect 19658 4326 19710 4378
rect 19722 4326 19774 4378
rect 19786 4326 19838 4378
rect 19850 4326 19902 4378
rect 19914 4326 19966 4378
rect 19978 4326 20030 4378
rect 27658 4326 27710 4378
rect 27722 4326 27774 4378
rect 27786 4326 27838 4378
rect 27850 4326 27902 4378
rect 27914 4326 27966 4378
rect 27978 4326 28030 4378
rect 1676 4224 1728 4276
rect 2964 4267 3016 4276
rect 2964 4233 2973 4267
rect 2973 4233 3007 4267
rect 3007 4233 3016 4267
rect 2964 4224 3016 4233
rect 4988 4224 5040 4276
rect 5448 4224 5500 4276
rect 7196 4224 7248 4276
rect 8208 4224 8260 4276
rect 17868 4267 17920 4276
rect 17868 4233 17877 4267
rect 17877 4233 17911 4267
rect 17911 4233 17920 4267
rect 17868 4224 17920 4233
rect 18420 4224 18472 4276
rect 22376 4224 22428 4276
rect 23296 4224 23348 4276
rect 5172 4156 5224 4208
rect 9312 4156 9364 4208
rect 11336 4156 11388 4208
rect 11796 4156 11848 4208
rect 12164 4156 12216 4208
rect 15384 4156 15436 4208
rect 15660 4199 15712 4208
rect 15660 4165 15669 4199
rect 15669 4165 15703 4199
rect 15703 4165 15712 4199
rect 15660 4156 15712 4165
rect 20444 4156 20496 4208
rect 22836 4156 22888 4208
rect 4620 4088 4672 4140
rect 5356 3952 5408 4004
rect 8116 4063 8168 4072
rect 8116 4029 8125 4063
rect 8125 4029 8159 4063
rect 8159 4029 8168 4063
rect 8116 4020 8168 4029
rect 8760 4063 8812 4072
rect 8760 4029 8769 4063
rect 8769 4029 8803 4063
rect 8803 4029 8812 4063
rect 8760 4020 8812 4029
rect 8944 4063 8996 4072
rect 8944 4029 8953 4063
rect 8953 4029 8987 4063
rect 8987 4029 8996 4063
rect 8944 4020 8996 4029
rect 10784 4063 10836 4072
rect 10784 4029 10793 4063
rect 10793 4029 10827 4063
rect 10827 4029 10836 4063
rect 10784 4020 10836 4029
rect 12072 4063 12124 4072
rect 12072 4029 12081 4063
rect 12081 4029 12115 4063
rect 12115 4029 12124 4063
rect 12072 4020 12124 4029
rect 11428 3884 11480 3936
rect 11888 3884 11940 3936
rect 12532 4088 12584 4140
rect 17316 4088 17368 4140
rect 22284 4131 22336 4140
rect 22284 4097 22293 4131
rect 22293 4097 22327 4131
rect 22327 4097 22336 4131
rect 22284 4088 22336 4097
rect 13912 4020 13964 4072
rect 18512 4063 18564 4072
rect 18512 4029 18521 4063
rect 18521 4029 18555 4063
rect 18555 4029 18564 4063
rect 18512 4020 18564 4029
rect 18604 3952 18656 4004
rect 20720 4020 20772 4072
rect 22008 4020 22060 4072
rect 24768 4020 24820 4072
rect 12808 3884 12860 3936
rect 17408 3884 17460 3936
rect 21456 3884 21508 3936
rect 22652 3927 22704 3936
rect 22652 3893 22661 3927
rect 22661 3893 22695 3927
rect 22695 3893 22704 3927
rect 22652 3884 22704 3893
rect 2918 3782 2970 3834
rect 2982 3782 3034 3834
rect 3046 3782 3098 3834
rect 3110 3782 3162 3834
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 10918 3782 10970 3834
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 11238 3782 11290 3834
rect 18918 3782 18970 3834
rect 18982 3782 19034 3834
rect 19046 3782 19098 3834
rect 19110 3782 19162 3834
rect 19174 3782 19226 3834
rect 19238 3782 19290 3834
rect 26918 3782 26970 3834
rect 26982 3782 27034 3834
rect 27046 3782 27098 3834
rect 27110 3782 27162 3834
rect 27174 3782 27226 3834
rect 27238 3782 27290 3834
rect 5172 3680 5224 3732
rect 8944 3680 8996 3732
rect 11796 3680 11848 3732
rect 12164 3680 12216 3732
rect 14740 3680 14792 3732
rect 18604 3723 18656 3732
rect 18604 3689 18613 3723
rect 18613 3689 18647 3723
rect 18647 3689 18656 3723
rect 18604 3680 18656 3689
rect 22836 3723 22888 3732
rect 22836 3689 22845 3723
rect 22845 3689 22879 3723
rect 22879 3689 22888 3723
rect 22836 3680 22888 3689
rect 3332 3544 3384 3596
rect 6828 3544 6880 3596
rect 8300 3544 8352 3596
rect 11520 3544 11572 3596
rect 11888 3587 11940 3596
rect 11888 3553 11897 3587
rect 11897 3553 11931 3587
rect 11931 3553 11940 3587
rect 11888 3544 11940 3553
rect 12716 3587 12768 3596
rect 12716 3553 12725 3587
rect 12725 3553 12759 3587
rect 12759 3553 12768 3587
rect 12716 3544 12768 3553
rect 12808 3587 12860 3596
rect 12808 3553 12817 3587
rect 12817 3553 12851 3587
rect 12851 3553 12860 3587
rect 12808 3544 12860 3553
rect 13820 3544 13872 3596
rect 14372 3587 14424 3596
rect 14372 3553 14381 3587
rect 14381 3553 14415 3587
rect 14415 3553 14424 3587
rect 14372 3544 14424 3553
rect 17316 3544 17368 3596
rect 21364 3544 21416 3596
rect 9312 3519 9364 3528
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 12164 3519 12216 3528
rect 12164 3485 12173 3519
rect 12173 3485 12207 3519
rect 12207 3485 12216 3519
rect 12164 3476 12216 3485
rect 15476 3476 15528 3528
rect 4068 3451 4120 3460
rect 4068 3417 4077 3451
rect 4077 3417 4111 3451
rect 4111 3417 4120 3451
rect 4068 3408 4120 3417
rect 5632 3408 5684 3460
rect 6828 3451 6880 3460
rect 6828 3417 6837 3451
rect 6837 3417 6871 3451
rect 6871 3417 6880 3451
rect 6828 3408 6880 3417
rect 7288 3408 7340 3460
rect 8760 3408 8812 3460
rect 9680 3408 9732 3460
rect 17868 3408 17920 3460
rect 8300 3383 8352 3392
rect 8300 3349 8309 3383
rect 8309 3349 8343 3383
rect 8343 3349 8352 3383
rect 8300 3340 8352 3349
rect 8944 3383 8996 3392
rect 8944 3349 8953 3383
rect 8953 3349 8987 3383
rect 8987 3349 8996 3383
rect 8944 3340 8996 3349
rect 12624 3383 12676 3392
rect 12624 3349 12633 3383
rect 12633 3349 12667 3383
rect 12667 3349 12676 3383
rect 12624 3340 12676 3349
rect 16304 3383 16356 3392
rect 16304 3349 16313 3383
rect 16313 3349 16347 3383
rect 16347 3349 16356 3383
rect 16304 3340 16356 3349
rect 17132 3340 17184 3392
rect 19524 3451 19576 3460
rect 19524 3417 19533 3451
rect 19533 3417 19567 3451
rect 19567 3417 19576 3451
rect 19524 3408 19576 3417
rect 20444 3340 20496 3392
rect 21456 3408 21508 3460
rect 21824 3408 21876 3460
rect 3658 3238 3710 3290
rect 3722 3238 3774 3290
rect 3786 3238 3838 3290
rect 3850 3238 3902 3290
rect 3914 3238 3966 3290
rect 3978 3238 4030 3290
rect 11658 3238 11710 3290
rect 11722 3238 11774 3290
rect 11786 3238 11838 3290
rect 11850 3238 11902 3290
rect 11914 3238 11966 3290
rect 11978 3238 12030 3290
rect 19658 3238 19710 3290
rect 19722 3238 19774 3290
rect 19786 3238 19838 3290
rect 19850 3238 19902 3290
rect 19914 3238 19966 3290
rect 19978 3238 20030 3290
rect 27658 3238 27710 3290
rect 27722 3238 27774 3290
rect 27786 3238 27838 3290
rect 27850 3238 27902 3290
rect 27914 3238 27966 3290
rect 27978 3238 28030 3290
rect 4068 3136 4120 3188
rect 5172 3136 5224 3188
rect 6828 3136 6880 3188
rect 8300 3136 8352 3188
rect 9312 3136 9364 3188
rect 10784 3136 10836 3188
rect 12624 3136 12676 3188
rect 16304 3136 16356 3188
rect 17868 3179 17920 3188
rect 17868 3145 17877 3179
rect 17877 3145 17911 3179
rect 17911 3145 17920 3179
rect 17868 3136 17920 3145
rect 19524 3136 19576 3188
rect 20444 3179 20496 3188
rect 20444 3145 20453 3179
rect 20453 3145 20487 3179
rect 20487 3145 20496 3179
rect 20444 3136 20496 3145
rect 22652 3136 22704 3188
rect 8944 3068 8996 3120
rect 9680 3068 9732 3120
rect 11428 3068 11480 3120
rect 5356 2932 5408 2984
rect 8116 2975 8168 2984
rect 8116 2941 8125 2975
rect 8125 2941 8159 2975
rect 8159 2941 8168 2975
rect 8116 2932 8168 2941
rect 12164 3000 12216 3052
rect 12716 3068 12768 3120
rect 17408 3111 17460 3120
rect 17408 3077 17417 3111
rect 17417 3077 17451 3111
rect 17451 3077 17460 3111
rect 17408 3068 17460 3077
rect 11520 2932 11572 2984
rect 17132 2932 17184 2984
rect 17224 2975 17276 2984
rect 17224 2941 17233 2975
rect 17233 2941 17267 2975
rect 17267 2941 17276 2975
rect 17224 2932 17276 2941
rect 20720 2975 20772 2984
rect 20720 2941 20729 2975
rect 20729 2941 20763 2975
rect 20763 2941 20772 2975
rect 20720 2932 20772 2941
rect 14096 2864 14148 2916
rect 2918 2694 2970 2746
rect 2982 2694 3034 2746
rect 3046 2694 3098 2746
rect 3110 2694 3162 2746
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 10918 2694 10970 2746
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 11238 2694 11290 2746
rect 18918 2694 18970 2746
rect 18982 2694 19034 2746
rect 19046 2694 19098 2746
rect 19110 2694 19162 2746
rect 19174 2694 19226 2746
rect 19238 2694 19290 2746
rect 26918 2694 26970 2746
rect 26982 2694 27034 2746
rect 27046 2694 27098 2746
rect 27110 2694 27162 2746
rect 27174 2694 27226 2746
rect 27238 2694 27290 2746
rect 3658 2150 3710 2202
rect 3722 2150 3774 2202
rect 3786 2150 3838 2202
rect 3850 2150 3902 2202
rect 3914 2150 3966 2202
rect 3978 2150 4030 2202
rect 11658 2150 11710 2202
rect 11722 2150 11774 2202
rect 11786 2150 11838 2202
rect 11850 2150 11902 2202
rect 11914 2150 11966 2202
rect 11978 2150 12030 2202
rect 19658 2150 19710 2202
rect 19722 2150 19774 2202
rect 19786 2150 19838 2202
rect 19850 2150 19902 2202
rect 19914 2150 19966 2202
rect 19978 2150 20030 2202
rect 27658 2150 27710 2202
rect 27722 2150 27774 2202
rect 27786 2150 27838 2202
rect 27850 2150 27902 2202
rect 27914 2150 27966 2202
rect 27978 2150 28030 2202
<< metal2 >>
rect 2916 27772 3292 27781
rect 2972 27770 2996 27772
rect 3052 27770 3076 27772
rect 3132 27770 3156 27772
rect 3212 27770 3236 27772
rect 2972 27718 2982 27770
rect 3226 27718 3236 27770
rect 2972 27716 2996 27718
rect 3052 27716 3076 27718
rect 3132 27716 3156 27718
rect 3212 27716 3236 27718
rect 2916 27707 3292 27716
rect 10916 27772 11292 27781
rect 10972 27770 10996 27772
rect 11052 27770 11076 27772
rect 11132 27770 11156 27772
rect 11212 27770 11236 27772
rect 10972 27718 10982 27770
rect 11226 27718 11236 27770
rect 10972 27716 10996 27718
rect 11052 27716 11076 27718
rect 11132 27716 11156 27718
rect 11212 27716 11236 27718
rect 10916 27707 11292 27716
rect 18916 27772 19292 27781
rect 18972 27770 18996 27772
rect 19052 27770 19076 27772
rect 19132 27770 19156 27772
rect 19212 27770 19236 27772
rect 18972 27718 18982 27770
rect 19226 27718 19236 27770
rect 18972 27716 18996 27718
rect 19052 27716 19076 27718
rect 19132 27716 19156 27718
rect 19212 27716 19236 27718
rect 18916 27707 19292 27716
rect 26916 27772 27292 27781
rect 26972 27770 26996 27772
rect 27052 27770 27076 27772
rect 27132 27770 27156 27772
rect 27212 27770 27236 27772
rect 26972 27718 26982 27770
rect 27226 27718 27236 27770
rect 26972 27716 26996 27718
rect 27052 27716 27076 27718
rect 27132 27716 27156 27718
rect 27212 27716 27236 27718
rect 26916 27707 27292 27716
rect 3656 27228 4032 27237
rect 3712 27226 3736 27228
rect 3792 27226 3816 27228
rect 3872 27226 3896 27228
rect 3952 27226 3976 27228
rect 3712 27174 3722 27226
rect 3966 27174 3976 27226
rect 3712 27172 3736 27174
rect 3792 27172 3816 27174
rect 3872 27172 3896 27174
rect 3952 27172 3976 27174
rect 3656 27163 4032 27172
rect 11656 27228 12032 27237
rect 11712 27226 11736 27228
rect 11792 27226 11816 27228
rect 11872 27226 11896 27228
rect 11952 27226 11976 27228
rect 11712 27174 11722 27226
rect 11966 27174 11976 27226
rect 11712 27172 11736 27174
rect 11792 27172 11816 27174
rect 11872 27172 11896 27174
rect 11952 27172 11976 27174
rect 11656 27163 12032 27172
rect 19656 27228 20032 27237
rect 19712 27226 19736 27228
rect 19792 27226 19816 27228
rect 19872 27226 19896 27228
rect 19952 27226 19976 27228
rect 19712 27174 19722 27226
rect 19966 27174 19976 27226
rect 19712 27172 19736 27174
rect 19792 27172 19816 27174
rect 19872 27172 19896 27174
rect 19952 27172 19976 27174
rect 19656 27163 20032 27172
rect 27656 27228 28032 27237
rect 27712 27226 27736 27228
rect 27792 27226 27816 27228
rect 27872 27226 27896 27228
rect 27952 27226 27976 27228
rect 27712 27174 27722 27226
rect 27966 27174 27976 27226
rect 27712 27172 27736 27174
rect 27792 27172 27816 27174
rect 27872 27172 27896 27174
rect 27952 27172 27976 27174
rect 27656 27163 28032 27172
rect 2916 26684 3292 26693
rect 2972 26682 2996 26684
rect 3052 26682 3076 26684
rect 3132 26682 3156 26684
rect 3212 26682 3236 26684
rect 2972 26630 2982 26682
rect 3226 26630 3236 26682
rect 2972 26628 2996 26630
rect 3052 26628 3076 26630
rect 3132 26628 3156 26630
rect 3212 26628 3236 26630
rect 2916 26619 3292 26628
rect 10916 26684 11292 26693
rect 10972 26682 10996 26684
rect 11052 26682 11076 26684
rect 11132 26682 11156 26684
rect 11212 26682 11236 26684
rect 10972 26630 10982 26682
rect 11226 26630 11236 26682
rect 10972 26628 10996 26630
rect 11052 26628 11076 26630
rect 11132 26628 11156 26630
rect 11212 26628 11236 26630
rect 10916 26619 11292 26628
rect 18916 26684 19292 26693
rect 18972 26682 18996 26684
rect 19052 26682 19076 26684
rect 19132 26682 19156 26684
rect 19212 26682 19236 26684
rect 18972 26630 18982 26682
rect 19226 26630 19236 26682
rect 18972 26628 18996 26630
rect 19052 26628 19076 26630
rect 19132 26628 19156 26630
rect 19212 26628 19236 26630
rect 18916 26619 19292 26628
rect 26916 26684 27292 26693
rect 26972 26682 26996 26684
rect 27052 26682 27076 26684
rect 27132 26682 27156 26684
rect 27212 26682 27236 26684
rect 26972 26630 26982 26682
rect 27226 26630 27236 26682
rect 26972 26628 26996 26630
rect 27052 26628 27076 26630
rect 27132 26628 27156 26630
rect 27212 26628 27236 26630
rect 26916 26619 27292 26628
rect 3656 26140 4032 26149
rect 3712 26138 3736 26140
rect 3792 26138 3816 26140
rect 3872 26138 3896 26140
rect 3952 26138 3976 26140
rect 3712 26086 3722 26138
rect 3966 26086 3976 26138
rect 3712 26084 3736 26086
rect 3792 26084 3816 26086
rect 3872 26084 3896 26086
rect 3952 26084 3976 26086
rect 3656 26075 4032 26084
rect 11656 26140 12032 26149
rect 11712 26138 11736 26140
rect 11792 26138 11816 26140
rect 11872 26138 11896 26140
rect 11952 26138 11976 26140
rect 11712 26086 11722 26138
rect 11966 26086 11976 26138
rect 11712 26084 11736 26086
rect 11792 26084 11816 26086
rect 11872 26084 11896 26086
rect 11952 26084 11976 26086
rect 11656 26075 12032 26084
rect 19656 26140 20032 26149
rect 19712 26138 19736 26140
rect 19792 26138 19816 26140
rect 19872 26138 19896 26140
rect 19952 26138 19976 26140
rect 19712 26086 19722 26138
rect 19966 26086 19976 26138
rect 19712 26084 19736 26086
rect 19792 26084 19816 26086
rect 19872 26084 19896 26086
rect 19952 26084 19976 26086
rect 19656 26075 20032 26084
rect 27656 26140 28032 26149
rect 27712 26138 27736 26140
rect 27792 26138 27816 26140
rect 27872 26138 27896 26140
rect 27952 26138 27976 26140
rect 27712 26086 27722 26138
rect 27966 26086 27976 26138
rect 27712 26084 27736 26086
rect 27792 26084 27816 26086
rect 27872 26084 27896 26086
rect 27952 26084 27976 26086
rect 27656 26075 28032 26084
rect 2916 25596 3292 25605
rect 2972 25594 2996 25596
rect 3052 25594 3076 25596
rect 3132 25594 3156 25596
rect 3212 25594 3236 25596
rect 2972 25542 2982 25594
rect 3226 25542 3236 25594
rect 2972 25540 2996 25542
rect 3052 25540 3076 25542
rect 3132 25540 3156 25542
rect 3212 25540 3236 25542
rect 2916 25531 3292 25540
rect 10916 25596 11292 25605
rect 10972 25594 10996 25596
rect 11052 25594 11076 25596
rect 11132 25594 11156 25596
rect 11212 25594 11236 25596
rect 10972 25542 10982 25594
rect 11226 25542 11236 25594
rect 10972 25540 10996 25542
rect 11052 25540 11076 25542
rect 11132 25540 11156 25542
rect 11212 25540 11236 25542
rect 10916 25531 11292 25540
rect 18916 25596 19292 25605
rect 18972 25594 18996 25596
rect 19052 25594 19076 25596
rect 19132 25594 19156 25596
rect 19212 25594 19236 25596
rect 18972 25542 18982 25594
rect 19226 25542 19236 25594
rect 18972 25540 18996 25542
rect 19052 25540 19076 25542
rect 19132 25540 19156 25542
rect 19212 25540 19236 25542
rect 18916 25531 19292 25540
rect 26916 25596 27292 25605
rect 26972 25594 26996 25596
rect 27052 25594 27076 25596
rect 27132 25594 27156 25596
rect 27212 25594 27236 25596
rect 26972 25542 26982 25594
rect 27226 25542 27236 25594
rect 26972 25540 26996 25542
rect 27052 25540 27076 25542
rect 27132 25540 27156 25542
rect 27212 25540 27236 25542
rect 26916 25531 27292 25540
rect 1216 25220 1268 25226
rect 1216 25162 1268 25168
rect 1228 25129 1256 25162
rect 2504 25152 2556 25158
rect 1214 25120 1270 25129
rect 2504 25094 2556 25100
rect 1214 25055 1270 25064
rect 1308 24812 1360 24818
rect 1308 24754 1360 24760
rect 1320 24585 1348 24754
rect 1306 24576 1362 24585
rect 1306 24511 1362 24520
rect 1308 24200 1360 24206
rect 1308 24142 1360 24148
rect 1320 24041 1348 24142
rect 2044 24064 2096 24070
rect 1306 24032 1362 24041
rect 2044 24006 2096 24012
rect 1306 23967 1362 23976
rect 1308 23724 1360 23730
rect 1308 23666 1360 23672
rect 1320 23497 1348 23666
rect 1400 23588 1452 23594
rect 1400 23530 1452 23536
rect 1306 23488 1362 23497
rect 1306 23423 1362 23432
rect 1412 23118 1440 23530
rect 1952 23520 2004 23526
rect 1952 23462 2004 23468
rect 1768 23316 1820 23322
rect 1768 23258 1820 23264
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1412 22953 1440 23054
rect 1398 22944 1454 22953
rect 1398 22879 1454 22888
rect 1216 22636 1268 22642
rect 1216 22578 1268 22584
rect 1228 22409 1256 22578
rect 1214 22400 1270 22409
rect 1214 22335 1270 22344
rect 1216 21956 1268 21962
rect 1216 21898 1268 21904
rect 1228 21865 1256 21898
rect 1214 21856 1270 21865
rect 1214 21791 1270 21800
rect 1308 21548 1360 21554
rect 1308 21490 1360 21496
rect 1216 21412 1268 21418
rect 1216 21354 1268 21360
rect 1228 20924 1256 21354
rect 1320 21321 1348 21490
rect 1584 21344 1636 21350
rect 1306 21312 1362 21321
rect 1584 21286 1636 21292
rect 1306 21247 1362 21256
rect 1308 20936 1360 20942
rect 1228 20896 1308 20924
rect 1308 20878 1360 20884
rect 1320 20777 1348 20878
rect 1596 20777 1624 21286
rect 1306 20768 1362 20777
rect 1306 20703 1362 20712
rect 1582 20768 1638 20777
rect 1582 20703 1638 20712
rect 1308 20460 1360 20466
rect 1308 20402 1360 20408
rect 1320 20233 1348 20402
rect 1676 20324 1728 20330
rect 1676 20266 1728 20272
rect 1306 20224 1362 20233
rect 1306 20159 1362 20168
rect 1308 19848 1360 19854
rect 1308 19790 1360 19796
rect 1320 19689 1348 19790
rect 1306 19680 1362 19689
rect 1306 19615 1362 19624
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1412 19145 1440 19314
rect 1398 19136 1454 19145
rect 1398 19071 1454 19080
rect 1308 18760 1360 18766
rect 1308 18702 1360 18708
rect 1320 18601 1348 18702
rect 1306 18592 1362 18601
rect 1306 18527 1362 18536
rect 1308 18284 1360 18290
rect 1308 18226 1360 18232
rect 1320 18057 1348 18226
rect 1584 18080 1636 18086
rect 1306 18048 1362 18057
rect 1584 18022 1636 18028
rect 1306 17983 1362 17992
rect 1216 17604 1268 17610
rect 1216 17546 1268 17552
rect 1228 17513 1256 17546
rect 1214 17504 1270 17513
rect 1214 17439 1270 17448
rect 1596 17270 1624 18022
rect 1584 17264 1636 17270
rect 1584 17206 1636 17212
rect 1308 17196 1360 17202
rect 1308 17138 1360 17144
rect 1320 16969 1348 17138
rect 1306 16960 1362 16969
rect 1306 16895 1362 16904
rect 1492 16516 1544 16522
rect 1492 16458 1544 16464
rect 1504 16425 1532 16458
rect 1490 16416 1546 16425
rect 1490 16351 1546 16360
rect 1582 16280 1638 16289
rect 1582 16215 1584 16224
rect 1636 16215 1638 16224
rect 1584 16186 1636 16192
rect 1308 16108 1360 16114
rect 1308 16050 1360 16056
rect 1320 15881 1348 16050
rect 1306 15872 1362 15881
rect 1306 15807 1362 15816
rect 1688 15570 1716 20266
rect 1780 16726 1808 23258
rect 1964 22642 1992 23462
rect 1952 22636 2004 22642
rect 1952 22578 2004 22584
rect 1860 21888 1912 21894
rect 1860 21830 1912 21836
rect 1768 16720 1820 16726
rect 1768 16662 1820 16668
rect 1676 15564 1728 15570
rect 1676 15506 1728 15512
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15337 1440 15438
rect 1872 15366 1900 21830
rect 1964 20874 1992 22578
rect 2056 22574 2084 24006
rect 2516 23594 2544 25094
rect 3656 25052 4032 25061
rect 3712 25050 3736 25052
rect 3792 25050 3816 25052
rect 3872 25050 3896 25052
rect 3952 25050 3976 25052
rect 3712 24998 3722 25050
rect 3966 24998 3976 25050
rect 3712 24996 3736 24998
rect 3792 24996 3816 24998
rect 3872 24996 3896 24998
rect 3952 24996 3976 24998
rect 3656 24987 4032 24996
rect 11656 25052 12032 25061
rect 11712 25050 11736 25052
rect 11792 25050 11816 25052
rect 11872 25050 11896 25052
rect 11952 25050 11976 25052
rect 11712 24998 11722 25050
rect 11966 24998 11976 25050
rect 11712 24996 11736 24998
rect 11792 24996 11816 24998
rect 11872 24996 11896 24998
rect 11952 24996 11976 24998
rect 11656 24987 12032 24996
rect 19656 25052 20032 25061
rect 19712 25050 19736 25052
rect 19792 25050 19816 25052
rect 19872 25050 19896 25052
rect 19952 25050 19976 25052
rect 19712 24998 19722 25050
rect 19966 24998 19976 25050
rect 19712 24996 19736 24998
rect 19792 24996 19816 24998
rect 19872 24996 19896 24998
rect 19952 24996 19976 24998
rect 19656 24987 20032 24996
rect 27656 25052 28032 25061
rect 27712 25050 27736 25052
rect 27792 25050 27816 25052
rect 27872 25050 27896 25052
rect 27952 25050 27976 25052
rect 27712 24998 27722 25050
rect 27966 24998 27976 25050
rect 27712 24996 27736 24998
rect 27792 24996 27816 24998
rect 27872 24996 27896 24998
rect 27952 24996 27976 24998
rect 27656 24987 28032 24996
rect 2688 24608 2740 24614
rect 2688 24550 2740 24556
rect 2700 23730 2728 24550
rect 2916 24508 3292 24517
rect 2972 24506 2996 24508
rect 3052 24506 3076 24508
rect 3132 24506 3156 24508
rect 3212 24506 3236 24508
rect 2972 24454 2982 24506
rect 3226 24454 3236 24506
rect 2972 24452 2996 24454
rect 3052 24452 3076 24454
rect 3132 24452 3156 24454
rect 3212 24452 3236 24454
rect 2916 24443 3292 24452
rect 10916 24508 11292 24517
rect 10972 24506 10996 24508
rect 11052 24506 11076 24508
rect 11132 24506 11156 24508
rect 11212 24506 11236 24508
rect 10972 24454 10982 24506
rect 11226 24454 11236 24506
rect 10972 24452 10996 24454
rect 11052 24452 11076 24454
rect 11132 24452 11156 24454
rect 11212 24452 11236 24454
rect 10916 24443 11292 24452
rect 18916 24508 19292 24517
rect 18972 24506 18996 24508
rect 19052 24506 19076 24508
rect 19132 24506 19156 24508
rect 19212 24506 19236 24508
rect 18972 24454 18982 24506
rect 19226 24454 19236 24506
rect 18972 24452 18996 24454
rect 19052 24452 19076 24454
rect 19132 24452 19156 24454
rect 19212 24452 19236 24454
rect 18916 24443 19292 24452
rect 26916 24508 27292 24517
rect 26972 24506 26996 24508
rect 27052 24506 27076 24508
rect 27132 24506 27156 24508
rect 27212 24506 27236 24508
rect 26972 24454 26982 24506
rect 27226 24454 27236 24506
rect 26972 24452 26996 24454
rect 27052 24452 27076 24454
rect 27132 24452 27156 24454
rect 27212 24452 27236 24454
rect 26916 24443 27292 24452
rect 5448 24268 5500 24274
rect 5448 24210 5500 24216
rect 3656 23964 4032 23973
rect 3712 23962 3736 23964
rect 3792 23962 3816 23964
rect 3872 23962 3896 23964
rect 3952 23962 3976 23964
rect 3712 23910 3722 23962
rect 3966 23910 3976 23962
rect 3712 23908 3736 23910
rect 3792 23908 3816 23910
rect 3872 23908 3896 23910
rect 3952 23908 3976 23910
rect 3656 23899 4032 23908
rect 5460 23730 5488 24210
rect 6828 24200 6880 24206
rect 6828 24142 6880 24148
rect 6840 23866 6868 24142
rect 6920 24132 6972 24138
rect 6920 24074 6972 24080
rect 7104 24132 7156 24138
rect 7104 24074 7156 24080
rect 6828 23860 6880 23866
rect 6828 23802 6880 23808
rect 2688 23724 2740 23730
rect 2688 23666 2740 23672
rect 3424 23724 3476 23730
rect 3424 23666 3476 23672
rect 3792 23724 3844 23730
rect 3792 23666 3844 23672
rect 5448 23724 5500 23730
rect 5448 23666 5500 23672
rect 2780 23656 2832 23662
rect 2780 23598 2832 23604
rect 2504 23588 2556 23594
rect 2504 23530 2556 23536
rect 2516 23186 2544 23530
rect 2596 23520 2648 23526
rect 2596 23462 2648 23468
rect 2504 23180 2556 23186
rect 2504 23122 2556 23128
rect 2608 23118 2636 23462
rect 2320 23112 2372 23118
rect 2320 23054 2372 23060
rect 2412 23112 2464 23118
rect 2412 23054 2464 23060
rect 2596 23112 2648 23118
rect 2792 23100 2820 23598
rect 3436 23526 3464 23666
rect 3700 23656 3752 23662
rect 3700 23598 3752 23604
rect 3424 23520 3476 23526
rect 3424 23462 3476 23468
rect 2916 23420 3292 23429
rect 2972 23418 2996 23420
rect 3052 23418 3076 23420
rect 3132 23418 3156 23420
rect 3212 23418 3236 23420
rect 2972 23366 2982 23418
rect 3226 23366 3236 23418
rect 2972 23364 2996 23366
rect 3052 23364 3076 23366
rect 3132 23364 3156 23366
rect 3212 23364 3236 23366
rect 2916 23355 3292 23364
rect 3436 23254 3464 23462
rect 3332 23248 3384 23254
rect 3332 23190 3384 23196
rect 3424 23248 3476 23254
rect 3424 23190 3476 23196
rect 2872 23112 2924 23118
rect 2792 23072 2872 23100
rect 2596 23054 2648 23060
rect 2872 23054 2924 23060
rect 2228 22636 2280 22642
rect 2228 22578 2280 22584
rect 2044 22568 2096 22574
rect 2096 22528 2176 22556
rect 2044 22510 2096 22516
rect 2044 22432 2096 22438
rect 2044 22374 2096 22380
rect 1952 20868 2004 20874
rect 1952 20810 2004 20816
rect 1952 19780 2004 19786
rect 1952 19722 2004 19728
rect 1860 15360 1912 15366
rect 1398 15328 1454 15337
rect 1860 15302 1912 15308
rect 1398 15263 1454 15272
rect 1412 15162 1440 15263
rect 1400 15156 1452 15162
rect 1400 15098 1452 15104
rect 1308 15020 1360 15026
rect 1308 14962 1360 14968
rect 1320 14793 1348 14962
rect 1872 14890 1900 15302
rect 1860 14884 1912 14890
rect 1860 14826 1912 14832
rect 1306 14784 1362 14793
rect 1306 14719 1362 14728
rect 1320 14618 1348 14719
rect 1308 14612 1360 14618
rect 1308 14554 1360 14560
rect 1308 14408 1360 14414
rect 1308 14350 1360 14356
rect 1320 14249 1348 14350
rect 1306 14240 1362 14249
rect 1306 14175 1362 14184
rect 1308 13932 1360 13938
rect 1308 13874 1360 13880
rect 1320 13705 1348 13874
rect 1306 13696 1362 13705
rect 1306 13631 1362 13640
rect 1216 13320 1268 13326
rect 1216 13262 1268 13268
rect 1228 13161 1256 13262
rect 1214 13152 1270 13161
rect 1214 13087 1270 13096
rect 1228 12986 1256 13087
rect 1216 12980 1268 12986
rect 1216 12922 1268 12928
rect 1308 12844 1360 12850
rect 1308 12786 1360 12792
rect 1320 12617 1348 12786
rect 1306 12608 1362 12617
rect 1306 12543 1362 12552
rect 1964 12306 1992 19722
rect 2056 16250 2084 22374
rect 2148 21690 2176 22528
rect 2136 21684 2188 21690
rect 2136 21626 2188 21632
rect 2240 20466 2268 22578
rect 2332 20482 2360 23054
rect 2424 22234 2452 23054
rect 2504 22976 2556 22982
rect 2504 22918 2556 22924
rect 2412 22228 2464 22234
rect 2412 22170 2464 22176
rect 2516 22114 2544 22918
rect 2884 22778 2912 23054
rect 2872 22772 2924 22778
rect 2872 22714 2924 22720
rect 2688 22636 2740 22642
rect 2688 22578 2740 22584
rect 2596 22432 2648 22438
rect 2596 22374 2648 22380
rect 2424 22086 2544 22114
rect 2424 21350 2452 22086
rect 2608 22030 2636 22374
rect 2596 22024 2648 22030
rect 2596 21966 2648 21972
rect 2700 21978 2728 22578
rect 2780 22500 2832 22506
rect 2780 22442 2832 22448
rect 2792 22098 2820 22442
rect 2916 22332 3292 22341
rect 2972 22330 2996 22332
rect 3052 22330 3076 22332
rect 3132 22330 3156 22332
rect 3212 22330 3236 22332
rect 2972 22278 2982 22330
rect 3226 22278 3236 22330
rect 2972 22276 2996 22278
rect 3052 22276 3076 22278
rect 3132 22276 3156 22278
rect 3212 22276 3236 22278
rect 2916 22267 3292 22276
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 2780 22092 2832 22098
rect 2780 22034 2832 22040
rect 2700 21962 2820 21978
rect 2700 21956 2832 21962
rect 2700 21950 2780 21956
rect 2504 21888 2556 21894
rect 2504 21830 2556 21836
rect 2412 21344 2464 21350
rect 2410 21312 2412 21321
rect 2464 21312 2466 21321
rect 2410 21247 2466 21256
rect 2228 20460 2280 20466
rect 2332 20454 2452 20482
rect 2228 20402 2280 20408
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 2240 19122 2268 20402
rect 2148 18358 2176 19110
rect 2240 19094 2360 19122
rect 2228 18692 2280 18698
rect 2228 18634 2280 18640
rect 2136 18352 2188 18358
rect 2136 18294 2188 18300
rect 2136 18216 2188 18222
rect 2136 18158 2188 18164
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 1952 12300 2004 12306
rect 1952 12242 2004 12248
rect 1308 12232 1360 12238
rect 1308 12174 1360 12180
rect 1320 12073 1348 12174
rect 1306 12064 1362 12073
rect 1306 11999 1362 12008
rect 1950 12064 2006 12073
rect 1950 11999 2006 12008
rect 1964 11762 1992 11999
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 1308 11688 1360 11694
rect 1308 11630 1360 11636
rect 1032 11620 1084 11626
rect 1032 11562 1084 11568
rect 1044 4457 1072 11562
rect 1320 11529 1348 11630
rect 1306 11520 1362 11529
rect 1306 11455 1362 11464
rect 2056 11218 2084 12582
rect 2148 11354 2176 18158
rect 2240 17678 2268 18634
rect 2332 18290 2360 19094
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2332 17882 2360 18226
rect 2320 17876 2372 17882
rect 2320 17818 2372 17824
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1412 10985 1440 11086
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1412 10810 1440 10911
rect 1400 10804 1452 10810
rect 1400 10746 1452 10752
rect 1308 10668 1360 10674
rect 1308 10610 1360 10616
rect 1320 10441 1348 10610
rect 1306 10432 1362 10441
rect 1306 10367 1362 10376
rect 1308 10056 1360 10062
rect 1308 9998 1360 10004
rect 1320 9897 1348 9998
rect 1306 9888 1362 9897
rect 1306 9823 1362 9832
rect 1596 9722 1624 11086
rect 2240 10538 2268 17614
rect 2332 16522 2360 17818
rect 2320 16516 2372 16522
rect 2320 16458 2372 16464
rect 2332 16182 2360 16458
rect 2320 16176 2372 16182
rect 2320 16118 2372 16124
rect 2424 15978 2452 20454
rect 2516 16794 2544 21830
rect 2700 21554 2728 21950
rect 2780 21898 2832 21904
rect 3252 21622 3280 22170
rect 3240 21616 3292 21622
rect 3240 21558 3292 21564
rect 2688 21548 2740 21554
rect 2688 21490 2740 21496
rect 2596 21480 2648 21486
rect 2596 21422 2648 21428
rect 2608 20330 2636 21422
rect 2700 20466 2728 21490
rect 2780 21344 2832 21350
rect 2780 21286 2832 21292
rect 2792 21010 2820 21286
rect 2916 21244 3292 21253
rect 2972 21242 2996 21244
rect 3052 21242 3076 21244
rect 3132 21242 3156 21244
rect 3212 21242 3236 21244
rect 2972 21190 2982 21242
rect 3226 21190 3236 21242
rect 2972 21188 2996 21190
rect 3052 21188 3076 21190
rect 3132 21188 3156 21190
rect 3212 21188 3236 21190
rect 2916 21179 3292 21188
rect 2780 21004 2832 21010
rect 2780 20946 2832 20952
rect 2964 20936 3016 20942
rect 2964 20878 3016 20884
rect 2780 20868 2832 20874
rect 2780 20810 2832 20816
rect 2688 20460 2740 20466
rect 2688 20402 2740 20408
rect 2596 20324 2648 20330
rect 2596 20266 2648 20272
rect 2608 19854 2636 20266
rect 2596 19848 2648 19854
rect 2596 19790 2648 19796
rect 2700 19514 2728 20402
rect 2688 19508 2740 19514
rect 2688 19450 2740 19456
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 2594 19272 2650 19281
rect 2594 19207 2650 19216
rect 2608 18834 2636 19207
rect 2596 18828 2648 18834
rect 2596 18770 2648 18776
rect 2700 18698 2728 19314
rect 2688 18692 2740 18698
rect 2688 18634 2740 18640
rect 2596 18352 2648 18358
rect 2596 18294 2648 18300
rect 2608 17082 2636 18294
rect 2700 18222 2728 18634
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 2792 17898 2820 20810
rect 2976 20369 3004 20878
rect 3056 20868 3108 20874
rect 3056 20810 3108 20816
rect 3068 20602 3096 20810
rect 3344 20806 3372 23190
rect 3712 23050 3740 23598
rect 3804 23118 3832 23666
rect 4252 23588 4304 23594
rect 4252 23530 4304 23536
rect 4264 23118 4292 23530
rect 4712 23316 4764 23322
rect 4712 23258 4764 23264
rect 4724 23118 4752 23258
rect 3792 23112 3844 23118
rect 3790 23080 3792 23089
rect 4068 23112 4120 23118
rect 3844 23080 3846 23089
rect 3700 23044 3752 23050
rect 4068 23054 4120 23060
rect 4252 23112 4304 23118
rect 4252 23054 4304 23060
rect 4712 23112 4764 23118
rect 4712 23054 4764 23060
rect 3790 23015 3846 23024
rect 3700 22986 3752 22992
rect 3516 22976 3568 22982
rect 3516 22918 3568 22924
rect 3424 22772 3476 22778
rect 3424 22714 3476 22720
rect 3436 22234 3464 22714
rect 3424 22228 3476 22234
rect 3424 22170 3476 22176
rect 3424 21888 3476 21894
rect 3424 21830 3476 21836
rect 3332 20800 3384 20806
rect 3332 20742 3384 20748
rect 3056 20596 3108 20602
rect 3056 20538 3108 20544
rect 2962 20360 3018 20369
rect 2962 20295 3018 20304
rect 3332 20256 3384 20262
rect 3332 20198 3384 20204
rect 2916 20156 3292 20165
rect 2972 20154 2996 20156
rect 3052 20154 3076 20156
rect 3132 20154 3156 20156
rect 3212 20154 3236 20156
rect 2972 20102 2982 20154
rect 3226 20102 3236 20154
rect 2972 20100 2996 20102
rect 3052 20100 3076 20102
rect 3132 20100 3156 20102
rect 3212 20100 3236 20102
rect 2916 20091 3292 20100
rect 2962 19952 3018 19961
rect 2962 19887 3018 19896
rect 2870 19408 2926 19417
rect 2870 19343 2872 19352
rect 2924 19343 2926 19352
rect 2872 19314 2924 19320
rect 2976 19174 3004 19887
rect 3056 19712 3108 19718
rect 3056 19654 3108 19660
rect 3068 19514 3096 19654
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 3068 19310 3096 19450
rect 3344 19334 3372 20198
rect 3436 19378 3464 21830
rect 3528 21146 3556 22918
rect 3656 22876 4032 22885
rect 3712 22874 3736 22876
rect 3792 22874 3816 22876
rect 3872 22874 3896 22876
rect 3952 22874 3976 22876
rect 3712 22822 3722 22874
rect 3966 22822 3976 22874
rect 3712 22820 3736 22822
rect 3792 22820 3816 22822
rect 3872 22820 3896 22822
rect 3952 22820 3976 22822
rect 3656 22811 4032 22820
rect 3976 22636 4028 22642
rect 4080 22624 4108 23054
rect 4160 22976 4212 22982
rect 4160 22918 4212 22924
rect 4252 22976 4304 22982
rect 4252 22918 4304 22924
rect 4028 22596 4108 22624
rect 3976 22578 4028 22584
rect 3988 22001 4016 22578
rect 4066 22536 4122 22545
rect 4066 22471 4122 22480
rect 3974 21992 4030 22001
rect 4080 21962 4108 22471
rect 4172 22098 4200 22918
rect 4160 22092 4212 22098
rect 4160 22034 4212 22040
rect 3974 21927 4030 21936
rect 4068 21956 4120 21962
rect 3988 21894 4016 21927
rect 4068 21898 4120 21904
rect 3976 21888 4028 21894
rect 3976 21830 4028 21836
rect 3656 21788 4032 21797
rect 3712 21786 3736 21788
rect 3792 21786 3816 21788
rect 3872 21786 3896 21788
rect 3952 21786 3976 21788
rect 3712 21734 3722 21786
rect 3966 21734 3976 21786
rect 3712 21732 3736 21734
rect 3792 21732 3816 21734
rect 3872 21732 3896 21734
rect 3952 21732 3976 21734
rect 3656 21723 4032 21732
rect 3608 21548 3660 21554
rect 3608 21490 3660 21496
rect 3516 21140 3568 21146
rect 3516 21082 3568 21088
rect 3620 21026 3648 21490
rect 3528 21010 3648 21026
rect 3516 21004 3648 21010
rect 3568 20998 3648 21004
rect 3516 20946 3568 20952
rect 3528 19990 3556 20946
rect 3656 20700 4032 20709
rect 3712 20698 3736 20700
rect 3792 20698 3816 20700
rect 3872 20698 3896 20700
rect 3952 20698 3976 20700
rect 3712 20646 3722 20698
rect 3966 20646 3976 20698
rect 3712 20644 3736 20646
rect 3792 20644 3816 20646
rect 3872 20644 3896 20646
rect 3952 20644 3976 20646
rect 3656 20635 4032 20644
rect 3516 19984 3568 19990
rect 3516 19926 3568 19932
rect 4080 19786 4108 21898
rect 4264 20942 4292 22918
rect 5460 22234 5488 23666
rect 6736 23656 6788 23662
rect 6736 23598 6788 23604
rect 5632 23520 5684 23526
rect 5632 23462 5684 23468
rect 5644 23254 5672 23462
rect 5632 23248 5684 23254
rect 5632 23190 5684 23196
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 4896 22092 4948 22098
rect 4896 22034 4948 22040
rect 4908 21962 4936 22034
rect 5460 22030 5488 22170
rect 5644 22030 5672 23190
rect 6368 23180 6420 23186
rect 6368 23122 6420 23128
rect 6184 22704 6236 22710
rect 6184 22646 6236 22652
rect 5724 22092 5776 22098
rect 5724 22034 5776 22040
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 5632 22024 5684 22030
rect 5632 21966 5684 21972
rect 4896 21956 4948 21962
rect 4896 21898 4948 21904
rect 4908 21690 4936 21898
rect 5356 21888 5408 21894
rect 5356 21830 5408 21836
rect 4896 21684 4948 21690
rect 4896 21626 4948 21632
rect 5368 21146 5396 21830
rect 5736 21622 5764 22034
rect 6196 22030 6224 22646
rect 6380 22438 6408 23122
rect 6368 22432 6420 22438
rect 6368 22374 6420 22380
rect 6380 22030 6408 22374
rect 5908 22024 5960 22030
rect 5908 21966 5960 21972
rect 6184 22024 6236 22030
rect 6184 21966 6236 21972
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 5816 21888 5868 21894
rect 5816 21830 5868 21836
rect 5828 21622 5856 21830
rect 5724 21616 5776 21622
rect 5724 21558 5776 21564
rect 5816 21616 5868 21622
rect 5816 21558 5868 21564
rect 5920 21468 5948 21966
rect 6092 21956 6144 21962
rect 6092 21898 6144 21904
rect 6472 21950 6684 21978
rect 6104 21690 6132 21898
rect 6092 21684 6144 21690
rect 6092 21626 6144 21632
rect 5736 21440 5948 21468
rect 5356 21140 5408 21146
rect 5356 21082 5408 21088
rect 4252 20936 4304 20942
rect 4252 20878 4304 20884
rect 5448 20936 5500 20942
rect 5448 20878 5500 20884
rect 4160 20800 4212 20806
rect 4160 20742 4212 20748
rect 4528 20800 4580 20806
rect 4528 20742 4580 20748
rect 4068 19780 4120 19786
rect 4068 19722 4120 19728
rect 3516 19712 3568 19718
rect 3516 19654 3568 19660
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 3252 19306 3372 19334
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3252 19242 3280 19306
rect 3240 19236 3292 19242
rect 3240 19178 3292 19184
rect 3332 19236 3384 19242
rect 3332 19178 3384 19184
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 2916 19068 3292 19077
rect 2972 19066 2996 19068
rect 3052 19066 3076 19068
rect 3132 19066 3156 19068
rect 3212 19066 3236 19068
rect 2972 19014 2982 19066
rect 3226 19014 3236 19066
rect 2972 19012 2996 19014
rect 3052 19012 3076 19014
rect 3132 19012 3156 19014
rect 3212 19012 3236 19014
rect 2916 19003 3292 19012
rect 3240 18964 3292 18970
rect 3344 18952 3372 19178
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 3436 18970 3464 19110
rect 3292 18924 3372 18952
rect 3424 18964 3476 18970
rect 3240 18906 3292 18912
rect 3424 18906 3476 18912
rect 3054 18864 3110 18873
rect 3054 18799 3110 18808
rect 3148 18828 3200 18834
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 2884 18222 2912 18702
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 3068 18154 3096 18799
rect 3148 18770 3200 18776
rect 3160 18426 3188 18770
rect 3252 18766 3280 18906
rect 3528 18766 3556 19654
rect 3656 19612 4032 19621
rect 3712 19610 3736 19612
rect 3792 19610 3816 19612
rect 3872 19610 3896 19612
rect 3952 19610 3976 19612
rect 3712 19558 3722 19610
rect 3966 19558 3976 19610
rect 3712 19556 3736 19558
rect 3792 19556 3816 19558
rect 3872 19556 3896 19558
rect 3952 19556 3976 19558
rect 3656 19547 4032 19556
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 3882 19408 3938 19417
rect 3882 19343 3938 19352
rect 3700 19304 3752 19310
rect 3700 19246 3752 19252
rect 3792 19304 3844 19310
rect 3792 19246 3844 19252
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3620 18902 3648 19110
rect 3608 18896 3660 18902
rect 3712 18873 3740 19246
rect 3608 18838 3660 18844
rect 3698 18864 3754 18873
rect 3698 18799 3754 18808
rect 3240 18760 3292 18766
rect 3516 18760 3568 18766
rect 3240 18702 3292 18708
rect 3330 18728 3386 18737
rect 3330 18663 3386 18672
rect 3436 18720 3516 18748
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 3344 18170 3372 18663
rect 3436 18290 3464 18720
rect 3516 18702 3568 18708
rect 3804 18630 3832 19246
rect 3896 18737 3924 19343
rect 3988 19310 4016 19450
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3882 18728 3938 18737
rect 3882 18663 3938 18672
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 3528 18358 3556 18566
rect 3656 18524 4032 18533
rect 3712 18522 3736 18524
rect 3792 18522 3816 18524
rect 3872 18522 3896 18524
rect 3952 18522 3976 18524
rect 3712 18470 3722 18522
rect 3966 18470 3976 18522
rect 3712 18468 3736 18470
rect 3792 18468 3816 18470
rect 3872 18468 3896 18470
rect 3952 18468 3976 18470
rect 3656 18459 4032 18468
rect 3516 18352 3568 18358
rect 3516 18294 3568 18300
rect 3424 18284 3476 18290
rect 3424 18226 3476 18232
rect 3976 18284 4028 18290
rect 4080 18272 4108 19314
rect 4028 18244 4108 18272
rect 3976 18226 4028 18232
rect 3056 18148 3108 18154
rect 3344 18142 3556 18170
rect 3056 18090 3108 18096
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 2916 17980 3292 17989
rect 2972 17978 2996 17980
rect 3052 17978 3076 17980
rect 3132 17978 3156 17980
rect 3212 17978 3236 17980
rect 2972 17926 2982 17978
rect 3226 17926 3236 17978
rect 2972 17924 2996 17926
rect 3052 17924 3076 17926
rect 3132 17924 3156 17926
rect 3212 17924 3236 17926
rect 2916 17915 3292 17924
rect 2700 17870 2820 17898
rect 2700 17728 2728 17870
rect 3436 17746 3464 18022
rect 3424 17740 3476 17746
rect 2700 17700 2820 17728
rect 2608 17054 2728 17082
rect 2596 16992 2648 16998
rect 2596 16934 2648 16940
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2608 16726 2636 16934
rect 2596 16720 2648 16726
rect 2596 16662 2648 16668
rect 2596 16244 2648 16250
rect 2596 16186 2648 16192
rect 2608 16114 2636 16186
rect 2700 16114 2728 17054
rect 2792 16590 2820 17700
rect 3424 17682 3476 17688
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 3068 17105 3096 17614
rect 3054 17096 3110 17105
rect 3054 17031 3110 17040
rect 2916 16892 3292 16901
rect 2972 16890 2996 16892
rect 3052 16890 3076 16892
rect 3132 16890 3156 16892
rect 3212 16890 3236 16892
rect 2972 16838 2982 16890
rect 3226 16838 3236 16890
rect 2972 16836 2996 16838
rect 3052 16836 3076 16838
rect 3132 16836 3156 16838
rect 3212 16836 3236 16838
rect 2916 16827 3292 16836
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 3424 16584 3476 16590
rect 3424 16526 3476 16532
rect 3056 16516 3108 16522
rect 3056 16458 3108 16464
rect 3068 16250 3096 16458
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3056 16244 3108 16250
rect 3056 16186 3108 16192
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 2412 15972 2464 15978
rect 2412 15914 2464 15920
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2332 15162 2360 15438
rect 2320 15156 2372 15162
rect 2320 15098 2372 15104
rect 2424 15094 2452 15438
rect 2516 15434 2544 16050
rect 2608 15638 2636 16050
rect 2916 15804 3292 15813
rect 2972 15802 2996 15804
rect 3052 15802 3076 15804
rect 3132 15802 3156 15804
rect 3212 15802 3236 15804
rect 2972 15750 2982 15802
rect 3226 15750 3236 15802
rect 2972 15748 2996 15750
rect 3052 15748 3076 15750
rect 3132 15748 3156 15750
rect 3212 15748 3236 15750
rect 2916 15739 3292 15748
rect 3344 15706 3372 16390
rect 3436 16250 3464 16526
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3528 16114 3556 18142
rect 4172 17882 4200 20742
rect 4252 20528 4304 20534
rect 4252 20470 4304 20476
rect 4264 19417 4292 20470
rect 4540 19990 4568 20742
rect 5460 20534 5488 20878
rect 5448 20528 5500 20534
rect 5448 20470 5500 20476
rect 5460 20262 5488 20470
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 4528 19984 4580 19990
rect 4528 19926 4580 19932
rect 4528 19440 4580 19446
rect 4250 19408 4306 19417
rect 4528 19382 4580 19388
rect 4250 19343 4306 19352
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 4160 17672 4212 17678
rect 4264 17660 4292 18906
rect 4540 18766 4568 19382
rect 5632 19372 5684 19378
rect 5736 19360 5764 21440
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 5920 21146 5948 21286
rect 5908 21140 5960 21146
rect 5908 21082 5960 21088
rect 6104 21026 6132 21626
rect 6472 21554 6500 21950
rect 6656 21894 6684 21950
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 6460 21548 6512 21554
rect 6460 21490 6512 21496
rect 6564 21350 6592 21830
rect 6552 21344 6604 21350
rect 6552 21286 6604 21292
rect 5920 20998 6132 21026
rect 5816 19916 5868 19922
rect 5816 19858 5868 19864
rect 5828 19417 5856 19858
rect 5684 19332 5764 19360
rect 5814 19408 5870 19417
rect 5920 19378 5948 20998
rect 6748 20398 6776 23598
rect 6840 23118 6868 23802
rect 6932 23730 6960 24074
rect 6920 23724 6972 23730
rect 6920 23666 6972 23672
rect 6932 23186 6960 23666
rect 7116 23526 7144 24074
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 8404 23730 8432 24006
rect 11656 23964 12032 23973
rect 11712 23962 11736 23964
rect 11792 23962 11816 23964
rect 11872 23962 11896 23964
rect 11952 23962 11976 23964
rect 11712 23910 11722 23962
rect 11966 23910 11976 23962
rect 11712 23908 11736 23910
rect 11792 23908 11816 23910
rect 11872 23908 11896 23910
rect 11952 23908 11976 23910
rect 11656 23899 12032 23908
rect 19656 23964 20032 23973
rect 19712 23962 19736 23964
rect 19792 23962 19816 23964
rect 19872 23962 19896 23964
rect 19952 23962 19976 23964
rect 19712 23910 19722 23962
rect 19966 23910 19976 23962
rect 19712 23908 19736 23910
rect 19792 23908 19816 23910
rect 19872 23908 19896 23910
rect 19952 23908 19976 23910
rect 19656 23899 20032 23908
rect 27656 23964 28032 23973
rect 27712 23962 27736 23964
rect 27792 23962 27816 23964
rect 27872 23962 27896 23964
rect 27952 23962 27976 23964
rect 27712 23910 27722 23962
rect 27966 23910 27976 23962
rect 27712 23908 27736 23910
rect 27792 23908 27816 23910
rect 27872 23908 27896 23910
rect 27952 23908 27976 23910
rect 27656 23899 28032 23908
rect 7840 23724 7892 23730
rect 7840 23666 7892 23672
rect 7932 23724 7984 23730
rect 7932 23666 7984 23672
rect 8392 23724 8444 23730
rect 8392 23666 8444 23672
rect 7656 23656 7708 23662
rect 7656 23598 7708 23604
rect 7104 23520 7156 23526
rect 7104 23462 7156 23468
rect 7668 23322 7696 23598
rect 7748 23520 7800 23526
rect 7748 23462 7800 23468
rect 7656 23316 7708 23322
rect 7656 23258 7708 23264
rect 6920 23180 6972 23186
rect 6920 23122 6972 23128
rect 7760 23118 7788 23462
rect 6828 23112 6880 23118
rect 6828 23054 6880 23060
rect 7104 23112 7156 23118
rect 7104 23054 7156 23060
rect 7196 23112 7248 23118
rect 7196 23054 7248 23060
rect 7748 23112 7800 23118
rect 7748 23054 7800 23060
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 6840 20058 6868 23054
rect 7116 22778 7144 23054
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 7208 22710 7236 23054
rect 7564 23044 7616 23050
rect 7564 22986 7616 22992
rect 7472 22772 7524 22778
rect 7472 22714 7524 22720
rect 7196 22704 7248 22710
rect 7196 22646 7248 22652
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 6932 21690 6960 21966
rect 6920 21684 6972 21690
rect 6920 21626 6972 21632
rect 7012 21412 7064 21418
rect 7012 21354 7064 21360
rect 7024 20942 7052 21354
rect 7196 21344 7248 21350
rect 7196 21286 7248 21292
rect 7208 20942 7236 21286
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 7196 20936 7248 20942
rect 7196 20878 7248 20884
rect 7380 20936 7432 20942
rect 7380 20878 7432 20884
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 6012 19378 6040 19790
rect 6184 19780 6236 19786
rect 6184 19722 6236 19728
rect 6196 19514 6224 19722
rect 6184 19508 6236 19514
rect 6184 19450 6236 19456
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 6748 19378 6776 19450
rect 5814 19343 5816 19352
rect 5632 19314 5684 19320
rect 5868 19343 5870 19352
rect 5908 19372 5960 19378
rect 5816 19314 5868 19320
rect 5908 19314 5960 19320
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 6368 19372 6420 19378
rect 6736 19372 6788 19378
rect 6420 19332 6736 19360
rect 6368 19314 6420 19320
rect 6736 19314 6788 19320
rect 5644 19281 5672 19314
rect 5630 19272 5686 19281
rect 5630 19207 5632 19216
rect 5684 19207 5686 19216
rect 5632 19178 5684 19184
rect 5920 19174 5948 19314
rect 6840 19310 6868 19994
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 4436 18624 4488 18630
rect 4436 18566 4488 18572
rect 4448 18426 4476 18566
rect 4436 18420 4488 18426
rect 4436 18362 4488 18368
rect 5552 18222 5580 19110
rect 6736 18692 6788 18698
rect 6736 18634 6788 18640
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 6748 17678 6776 18634
rect 7392 17882 7420 20878
rect 7484 20058 7512 22714
rect 7576 22166 7604 22986
rect 7748 22636 7800 22642
rect 7748 22578 7800 22584
rect 7564 22160 7616 22166
rect 7564 22102 7616 22108
rect 7760 21554 7788 22578
rect 7852 22506 7880 23666
rect 7944 23322 7972 23666
rect 9036 23588 9088 23594
rect 9036 23530 9088 23536
rect 8760 23520 8812 23526
rect 8760 23462 8812 23468
rect 7932 23316 7984 23322
rect 7932 23258 7984 23264
rect 8116 23248 8168 23254
rect 8116 23190 8168 23196
rect 7932 22636 7984 22642
rect 8128 22624 8156 23190
rect 8484 23180 8536 23186
rect 8484 23122 8536 23128
rect 7984 22596 8156 22624
rect 7932 22578 7984 22584
rect 7840 22500 7892 22506
rect 7840 22442 7892 22448
rect 7944 22234 7972 22578
rect 7932 22228 7984 22234
rect 7932 22170 7984 22176
rect 8496 21622 8524 23122
rect 8772 22098 8800 23462
rect 8944 22976 8996 22982
rect 8944 22918 8996 22924
rect 8760 22092 8812 22098
rect 8760 22034 8812 22040
rect 8576 21888 8628 21894
rect 8576 21830 8628 21836
rect 8484 21616 8536 21622
rect 8484 21558 8536 21564
rect 7748 21548 7800 21554
rect 7748 21490 7800 21496
rect 7932 21548 7984 21554
rect 7932 21490 7984 21496
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 7484 19446 7512 19994
rect 7472 19440 7524 19446
rect 7472 19382 7524 19388
rect 7944 19310 7972 21490
rect 8300 21412 8352 21418
rect 8300 21354 8352 21360
rect 8312 21078 8340 21354
rect 8300 21072 8352 21078
rect 8300 21014 8352 21020
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 8208 19916 8260 19922
rect 8208 19858 8260 19864
rect 8036 19378 8064 19858
rect 8220 19514 8248 19858
rect 8208 19508 8260 19514
rect 8208 19450 8260 19456
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 7932 19304 7984 19310
rect 7932 19246 7984 19252
rect 8220 19174 8248 19450
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 8484 18148 8536 18154
rect 8484 18090 8536 18096
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 4212 17632 4292 17660
rect 5816 17672 5868 17678
rect 4160 17614 4212 17620
rect 5816 17614 5868 17620
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 3656 17436 4032 17445
rect 3712 17434 3736 17436
rect 3792 17434 3816 17436
rect 3872 17434 3896 17436
rect 3952 17434 3976 17436
rect 3712 17382 3722 17434
rect 3966 17382 3976 17434
rect 3712 17380 3736 17382
rect 3792 17380 3816 17382
rect 3872 17380 3896 17382
rect 3952 17380 3976 17382
rect 3656 17371 4032 17380
rect 3608 16992 3660 16998
rect 3608 16934 3660 16940
rect 3620 16590 3648 16934
rect 3608 16584 3660 16590
rect 3608 16526 3660 16532
rect 3656 16348 4032 16357
rect 3712 16346 3736 16348
rect 3792 16346 3816 16348
rect 3872 16346 3896 16348
rect 3952 16346 3976 16348
rect 3712 16294 3722 16346
rect 3966 16294 3976 16346
rect 3712 16292 3736 16294
rect 3792 16292 3816 16294
rect 3872 16292 3896 16294
rect 3952 16292 3976 16294
rect 3656 16283 4032 16292
rect 3608 16244 3660 16250
rect 3608 16186 3660 16192
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3424 15972 3476 15978
rect 3424 15914 3476 15920
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 3332 15496 3384 15502
rect 3252 15456 3332 15484
rect 2504 15428 2556 15434
rect 2504 15370 2556 15376
rect 2688 15428 2740 15434
rect 2688 15370 2740 15376
rect 2412 15088 2464 15094
rect 2412 15030 2464 15036
rect 2504 14952 2556 14958
rect 2504 14894 2556 14900
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2424 13802 2452 14350
rect 2412 13796 2464 13802
rect 2412 13738 2464 13744
rect 2424 12782 2452 13738
rect 2516 13326 2544 14894
rect 2608 14550 2636 14894
rect 2596 14544 2648 14550
rect 2596 14486 2648 14492
rect 2700 14414 2728 15370
rect 2962 15056 3018 15065
rect 2962 14991 2964 15000
rect 3016 14991 3018 15000
rect 2964 14962 3016 14968
rect 3252 14890 3280 15456
rect 3332 15438 3384 15444
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 2916 14716 3292 14725
rect 2972 14714 2996 14716
rect 3052 14714 3076 14716
rect 3132 14714 3156 14716
rect 3212 14714 3236 14716
rect 2972 14662 2982 14714
rect 3226 14662 3236 14714
rect 2972 14660 2996 14662
rect 3052 14660 3076 14662
rect 3132 14660 3156 14662
rect 3212 14660 3236 14662
rect 2916 14651 3292 14660
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 3148 14340 3200 14346
rect 3148 14282 3200 14288
rect 3160 14006 3188 14282
rect 3148 14000 3200 14006
rect 2962 13968 3018 13977
rect 3148 13942 3200 13948
rect 2962 13903 2964 13912
rect 3016 13903 3018 13912
rect 2964 13874 3016 13880
rect 3344 13802 3372 15302
rect 3436 14346 3464 15914
rect 3528 15162 3556 16050
rect 3620 15434 3648 16186
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 3896 15706 3924 15914
rect 3884 15700 3936 15706
rect 3884 15642 3936 15648
rect 3608 15428 3660 15434
rect 3608 15370 3660 15376
rect 3656 15260 4032 15269
rect 3712 15258 3736 15260
rect 3792 15258 3816 15260
rect 3872 15258 3896 15260
rect 3952 15258 3976 15260
rect 3712 15206 3722 15258
rect 3966 15206 3976 15258
rect 3712 15204 3736 15206
rect 3792 15204 3816 15206
rect 3872 15204 3896 15206
rect 3952 15204 3976 15206
rect 3656 15195 4032 15204
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 4080 14958 4108 15982
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3712 14482 3740 14894
rect 4172 14498 4200 17614
rect 4528 17604 4580 17610
rect 4528 17546 4580 17552
rect 5724 17604 5776 17610
rect 5724 17546 5776 17552
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 4264 14618 4292 16050
rect 4436 15088 4488 15094
rect 4436 15030 4488 15036
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 3700 14476 3752 14482
rect 4172 14470 4292 14498
rect 3700 14418 3752 14424
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 3424 14340 3476 14346
rect 3424 14282 3476 14288
rect 3528 14074 3556 14350
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 3656 14172 4032 14181
rect 3712 14170 3736 14172
rect 3792 14170 3816 14172
rect 3872 14170 3896 14172
rect 3952 14170 3976 14172
rect 3712 14118 3722 14170
rect 3966 14118 3976 14170
rect 3712 14116 3736 14118
rect 3792 14116 3816 14118
rect 3872 14116 3896 14118
rect 3952 14116 3976 14118
rect 3656 14107 4032 14116
rect 4080 14074 4108 14214
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 3514 13968 3570 13977
rect 3882 13968 3938 13977
rect 3514 13903 3570 13912
rect 3792 13932 3844 13938
rect 3332 13796 3384 13802
rect 3332 13738 3384 13744
rect 2596 13728 2648 13734
rect 3056 13728 3108 13734
rect 2596 13670 2648 13676
rect 2792 13688 3056 13716
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2608 12850 2636 13670
rect 2792 13394 2820 13688
rect 3056 13670 3108 13676
rect 2916 13628 3292 13637
rect 2972 13626 2996 13628
rect 3052 13626 3076 13628
rect 3132 13626 3156 13628
rect 3212 13626 3236 13628
rect 2972 13574 2982 13626
rect 3226 13574 3236 13626
rect 2972 13572 2996 13574
rect 3052 13572 3076 13574
rect 3132 13572 3156 13574
rect 3212 13572 3236 13574
rect 2916 13563 3292 13572
rect 3528 13530 3556 13903
rect 3882 13903 3884 13912
rect 3792 13874 3844 13880
rect 3936 13903 3938 13912
rect 3976 13932 4028 13938
rect 3884 13874 3936 13880
rect 3976 13874 4028 13880
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 3804 13734 3832 13874
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3988 13462 4016 13874
rect 4172 13530 4200 13874
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 2872 13456 2924 13462
rect 2872 13398 2924 13404
rect 3976 13456 4028 13462
rect 3976 13398 4028 13404
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 2424 11898 2452 12718
rect 2608 12170 2636 12786
rect 2596 12164 2648 12170
rect 2596 12106 2648 12112
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2332 11150 2360 11698
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2228 10532 2280 10538
rect 2228 10474 2280 10480
rect 2608 10266 2636 12106
rect 2792 11762 2820 12922
rect 2884 12714 2912 13398
rect 4264 13394 4292 14470
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2976 12714 3004 12786
rect 3252 12782 3280 13262
rect 3424 13252 3476 13258
rect 3424 13194 3476 13200
rect 3436 12986 3464 13194
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 2916 12540 3292 12549
rect 2972 12538 2996 12540
rect 3052 12538 3076 12540
rect 3132 12538 3156 12540
rect 3212 12538 3236 12540
rect 2972 12486 2982 12538
rect 3226 12486 3236 12538
rect 2972 12484 2996 12486
rect 3052 12484 3076 12486
rect 3132 12484 3156 12486
rect 3212 12484 3236 12486
rect 2916 12475 3292 12484
rect 3344 12442 3372 12786
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2700 11354 2728 11630
rect 3344 11558 3372 12378
rect 3436 11642 3464 12718
rect 3528 11744 3556 13330
rect 4448 13326 4476 15030
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 3656 13084 4032 13093
rect 3712 13082 3736 13084
rect 3792 13082 3816 13084
rect 3872 13082 3896 13084
rect 3952 13082 3976 13084
rect 3712 13030 3722 13082
rect 3966 13030 3976 13082
rect 3712 13028 3736 13030
rect 3792 13028 3816 13030
rect 3872 13028 3896 13030
rect 3952 13028 3976 13030
rect 3656 13019 4032 13028
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 3620 12714 3648 12922
rect 4080 12918 4108 13194
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 3608 12708 3660 12714
rect 3608 12650 3660 12656
rect 3620 12374 3648 12650
rect 3608 12368 3660 12374
rect 3608 12310 3660 12316
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 3656 11996 4032 12005
rect 3712 11994 3736 11996
rect 3792 11994 3816 11996
rect 3872 11994 3896 11996
rect 3952 11994 3976 11996
rect 3712 11942 3722 11994
rect 3966 11942 3976 11994
rect 3712 11940 3736 11942
rect 3792 11940 3816 11942
rect 3872 11940 3896 11942
rect 3952 11940 3976 11942
rect 3656 11931 4032 11940
rect 3528 11716 3740 11744
rect 3436 11614 3556 11642
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 2916 11452 3292 11461
rect 2972 11450 2996 11452
rect 3052 11450 3076 11452
rect 3132 11450 3156 11452
rect 3212 11450 3236 11452
rect 2972 11398 2982 11450
rect 3226 11398 3236 11450
rect 2972 11396 2996 11398
rect 3052 11396 3076 11398
rect 3132 11396 3156 11398
rect 3212 11396 3236 11398
rect 2916 11387 3292 11396
rect 3528 11370 3556 11614
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 3344 11342 3556 11370
rect 3344 10674 3372 11342
rect 3516 11144 3568 11150
rect 3620 11132 3648 11494
rect 3712 11354 3740 11716
rect 3790 11384 3846 11393
rect 3700 11348 3752 11354
rect 3790 11319 3792 11328
rect 3700 11290 3752 11296
rect 3844 11319 3846 11328
rect 3884 11348 3936 11354
rect 3792 11290 3844 11296
rect 3884 11290 3936 11296
rect 3568 11104 3648 11132
rect 3516 11086 3568 11092
rect 3896 11014 3924 11290
rect 4172 11218 4200 12038
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4264 11150 4292 11494
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4356 11150 4384 11222
rect 4448 11150 4476 13262
rect 4540 13190 4568 17546
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5460 15910 5488 17138
rect 5736 17134 5764 17546
rect 5724 17128 5776 17134
rect 5724 17070 5776 17076
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5460 15434 5488 15846
rect 5736 15706 5764 17070
rect 5828 17066 5856 17614
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 6276 17264 6328 17270
rect 6276 17206 6328 17212
rect 5816 17060 5868 17066
rect 5816 17002 5868 17008
rect 6184 16720 6236 16726
rect 6184 16662 6236 16668
rect 5908 16584 5960 16590
rect 5906 16552 5908 16561
rect 5960 16552 5962 16561
rect 5906 16487 5962 16496
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5736 15570 5764 15642
rect 5724 15564 5776 15570
rect 5724 15506 5776 15512
rect 5448 15428 5500 15434
rect 5448 15370 5500 15376
rect 5920 15366 5948 16487
rect 6000 16176 6052 16182
rect 6000 16118 6052 16124
rect 6092 16176 6144 16182
rect 6092 16118 6144 16124
rect 5908 15360 5960 15366
rect 5908 15302 5960 15308
rect 6012 14958 6040 16118
rect 6104 15502 6132 16118
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6000 14952 6052 14958
rect 6000 14894 6052 14900
rect 5724 14884 5776 14890
rect 5724 14826 5776 14832
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 5736 12238 5764 14826
rect 6012 14006 6040 14894
rect 6000 14000 6052 14006
rect 6000 13942 6052 13948
rect 6012 13326 6040 13942
rect 6104 13870 6132 15438
rect 6196 14958 6224 16662
rect 6184 14952 6236 14958
rect 6184 14894 6236 14900
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6104 13530 6132 13806
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6288 13394 6316 17206
rect 6380 17202 6408 17478
rect 6840 17270 6868 17682
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6644 17128 6696 17134
rect 6644 17070 6696 17076
rect 6736 17128 6788 17134
rect 6736 17070 6788 17076
rect 6656 16794 6684 17070
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6748 16726 6776 17070
rect 6840 16998 6868 17206
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6736 16720 6788 16726
rect 6736 16662 6788 16668
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6472 15570 6500 16526
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6564 14226 6592 16526
rect 6644 16516 6696 16522
rect 6644 16458 6696 16464
rect 6656 15502 6684 16458
rect 6748 15910 6776 16662
rect 6932 16590 6960 17614
rect 7116 17338 7144 17614
rect 7748 17604 7800 17610
rect 7748 17546 7800 17552
rect 7760 17338 7788 17546
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 7484 16794 7512 17138
rect 7840 17060 7892 17066
rect 7840 17002 7892 17008
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 7116 16250 7144 16526
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 7196 16176 7248 16182
rect 7196 16118 7248 16124
rect 7288 16176 7340 16182
rect 7288 16118 7340 16124
rect 6736 15904 6788 15910
rect 6736 15846 6788 15852
rect 7208 15706 7236 16118
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7300 15638 7328 16118
rect 7288 15632 7340 15638
rect 7288 15574 7340 15580
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6656 15026 6684 15438
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6472 14198 6592 14226
rect 6472 13938 6500 14198
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 6472 13682 6500 13874
rect 6472 13654 6592 13682
rect 6460 13524 6512 13530
rect 6460 13466 6512 13472
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 6288 12850 6316 13330
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6288 12646 6316 12786
rect 6472 12782 6500 13466
rect 6564 13326 6592 13654
rect 7024 13530 7052 13874
rect 7104 13796 7156 13802
rect 7104 13738 7156 13744
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6564 13190 6592 13262
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6564 12986 6592 13126
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 6276 12640 6328 12646
rect 6276 12582 6328 12588
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3884 11008 3936 11014
rect 3884 10950 3936 10956
rect 3528 10810 3556 10950
rect 3656 10908 4032 10917
rect 3712 10906 3736 10908
rect 3792 10906 3816 10908
rect 3872 10906 3896 10908
rect 3952 10906 3976 10908
rect 3712 10854 3722 10906
rect 3966 10854 3976 10906
rect 3712 10852 3736 10854
rect 3792 10852 3816 10854
rect 3872 10852 3896 10854
rect 3952 10852 3976 10854
rect 3656 10843 4032 10852
rect 3516 10804 3568 10810
rect 3516 10746 3568 10752
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 1584 9716 1636 9722
rect 1584 9658 1636 9664
rect 1308 9580 1360 9586
rect 1308 9522 1360 9528
rect 1320 9353 1348 9522
rect 1306 9344 1362 9353
rect 1306 9279 1362 9288
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1308 8832 1360 8838
rect 1306 8800 1308 8809
rect 1360 8800 1362 8809
rect 1306 8735 1362 8744
rect 1320 8498 1348 8735
rect 1308 8492 1360 8498
rect 1308 8434 1360 8440
rect 1306 8256 1362 8265
rect 1306 8191 1362 8200
rect 1320 7954 1348 8191
rect 1308 7948 1360 7954
rect 1308 7890 1360 7896
rect 1216 7880 1268 7886
rect 1216 7822 1268 7828
rect 1228 7721 1256 7822
rect 1214 7712 1270 7721
rect 1214 7647 1270 7656
rect 1320 7546 1348 7890
rect 1596 7546 1624 8910
rect 2044 8900 2096 8906
rect 2044 8842 2096 8848
rect 2056 8634 2084 8842
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2792 8430 2820 10542
rect 2916 10364 3292 10373
rect 2972 10362 2996 10364
rect 3052 10362 3076 10364
rect 3132 10362 3156 10364
rect 3212 10362 3236 10364
rect 2972 10310 2982 10362
rect 3226 10310 3236 10362
rect 2972 10308 2996 10310
rect 3052 10308 3076 10310
rect 3132 10308 3156 10310
rect 3212 10308 3236 10310
rect 2916 10299 3292 10308
rect 3656 9820 4032 9829
rect 3712 9818 3736 9820
rect 3792 9818 3816 9820
rect 3872 9818 3896 9820
rect 3952 9818 3976 9820
rect 3712 9766 3722 9818
rect 3966 9766 3976 9818
rect 3712 9764 3736 9766
rect 3792 9764 3816 9766
rect 3872 9764 3896 9766
rect 3952 9764 3976 9766
rect 3656 9755 4032 9764
rect 2916 9276 3292 9285
rect 2972 9274 2996 9276
rect 3052 9274 3076 9276
rect 3132 9274 3156 9276
rect 3212 9274 3236 9276
rect 2972 9222 2982 9274
rect 3226 9222 3236 9274
rect 2972 9220 2996 9222
rect 3052 9220 3076 9222
rect 3132 9220 3156 9222
rect 3212 9220 3236 9222
rect 2916 9211 3292 9220
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 3160 8362 3188 8910
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 1308 7540 1360 7546
rect 1308 7482 1360 7488
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1596 7410 1624 7482
rect 2596 7472 2648 7478
rect 2596 7414 2648 7420
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1214 7168 1270 7177
rect 1214 7103 1270 7112
rect 1228 6730 1256 7103
rect 1308 6792 1360 6798
rect 1308 6734 1360 6740
rect 1216 6724 1268 6730
rect 1216 6666 1268 6672
rect 1320 6633 1348 6734
rect 1306 6624 1362 6633
rect 1306 6559 1362 6568
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 1320 6089 1348 6258
rect 1306 6080 1362 6089
rect 1306 6015 1362 6024
rect 1308 5704 1360 5710
rect 1308 5646 1360 5652
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 1320 5545 1348 5646
rect 1306 5536 1362 5545
rect 1306 5471 1362 5480
rect 2516 5370 2544 5646
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 1308 5228 1360 5234
rect 1308 5170 1360 5176
rect 1320 5001 1348 5170
rect 2608 5098 2636 7414
rect 2792 6934 2820 8230
rect 2916 8188 3292 8197
rect 2972 8186 2996 8188
rect 3052 8186 3076 8188
rect 3132 8186 3156 8188
rect 3212 8186 3236 8188
rect 2972 8134 2982 8186
rect 3226 8134 3236 8186
rect 2972 8132 2996 8134
rect 3052 8132 3076 8134
rect 3132 8132 3156 8134
rect 3212 8132 3236 8134
rect 2916 8123 3292 8132
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 2916 7100 3292 7109
rect 2972 7098 2996 7100
rect 3052 7098 3076 7100
rect 3132 7098 3156 7100
rect 3212 7098 3236 7100
rect 2972 7046 2982 7098
rect 3226 7046 3236 7098
rect 2972 7044 2996 7046
rect 3052 7044 3076 7046
rect 3132 7044 3156 7046
rect 3212 7044 3236 7046
rect 2916 7035 3292 7044
rect 2688 6928 2740 6934
rect 2688 6870 2740 6876
rect 2780 6928 2832 6934
rect 2780 6870 2832 6876
rect 2700 5370 2728 6870
rect 2916 6012 3292 6021
rect 2972 6010 2996 6012
rect 3052 6010 3076 6012
rect 3132 6010 3156 6012
rect 3212 6010 3236 6012
rect 2972 5958 2982 6010
rect 3226 5958 3236 6010
rect 2972 5956 2996 5958
rect 3052 5956 3076 5958
rect 3132 5956 3156 5958
rect 3212 5956 3236 5958
rect 2916 5947 3292 5956
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 3068 5234 3096 5850
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3252 5234 3280 5510
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 2596 5092 2648 5098
rect 2596 5034 2648 5040
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 1306 4992 1362 5001
rect 1306 4927 1362 4936
rect 2792 4622 2820 5034
rect 3068 5030 3096 5170
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 2916 4924 3292 4933
rect 2972 4922 2996 4924
rect 3052 4922 3076 4924
rect 3132 4922 3156 4924
rect 3212 4922 3236 4924
rect 2972 4870 2982 4922
rect 3226 4870 3236 4922
rect 2972 4868 2996 4870
rect 3052 4868 3076 4870
rect 3132 4868 3156 4870
rect 3212 4868 3236 4870
rect 2916 4859 3292 4868
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 1030 4448 1086 4457
rect 1030 4383 1086 4392
rect 1688 4282 1716 4490
rect 2976 4282 3004 4762
rect 3344 4690 3372 7482
rect 3436 6866 3464 8910
rect 3528 8634 3556 9046
rect 3656 8732 4032 8741
rect 3712 8730 3736 8732
rect 3792 8730 3816 8732
rect 3872 8730 3896 8732
rect 3952 8730 3976 8732
rect 3712 8678 3722 8730
rect 3966 8678 3976 8730
rect 3712 8676 3736 8678
rect 3792 8676 3816 8678
rect 3872 8676 3896 8678
rect 3952 8676 3976 8678
rect 3656 8667 4032 8676
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 3712 8090 3740 8434
rect 3700 8084 3752 8090
rect 3700 8026 3752 8032
rect 3804 7818 3832 8434
rect 3516 7812 3568 7818
rect 3516 7754 3568 7760
rect 3792 7812 3844 7818
rect 3792 7754 3844 7760
rect 3528 7410 3556 7754
rect 3896 7750 3924 8434
rect 4172 8022 4200 8434
rect 4264 8362 4292 9114
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 4356 7954 4384 8774
rect 4448 8022 4476 11086
rect 4816 10810 4844 11086
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 6932 10742 6960 13330
rect 7116 13258 7144 13738
rect 7852 13394 7880 17002
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8208 16516 8260 16522
rect 8208 16458 8260 16464
rect 8220 16250 8248 16458
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8312 15978 8340 16594
rect 8404 16590 8432 17138
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8300 15972 8352 15978
rect 8300 15914 8352 15920
rect 8392 15632 8444 15638
rect 8392 15574 8444 15580
rect 8024 15088 8076 15094
rect 8024 15030 8076 15036
rect 8036 14006 8064 15030
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 8036 13462 8064 13942
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8128 13530 8156 13874
rect 8404 13734 8432 15574
rect 8496 14074 8524 18090
rect 8588 16794 8616 21830
rect 8956 21078 8984 22918
rect 9048 22030 9076 23530
rect 10916 23420 11292 23429
rect 10972 23418 10996 23420
rect 11052 23418 11076 23420
rect 11132 23418 11156 23420
rect 11212 23418 11236 23420
rect 10972 23366 10982 23418
rect 11226 23366 11236 23418
rect 10972 23364 10996 23366
rect 11052 23364 11076 23366
rect 11132 23364 11156 23366
rect 11212 23364 11236 23366
rect 10916 23355 11292 23364
rect 18916 23420 19292 23429
rect 18972 23418 18996 23420
rect 19052 23418 19076 23420
rect 19132 23418 19156 23420
rect 19212 23418 19236 23420
rect 18972 23366 18982 23418
rect 19226 23366 19236 23418
rect 18972 23364 18996 23366
rect 19052 23364 19076 23366
rect 19132 23364 19156 23366
rect 19212 23364 19236 23366
rect 18916 23355 19292 23364
rect 26916 23420 27292 23429
rect 26972 23418 26996 23420
rect 27052 23418 27076 23420
rect 27132 23418 27156 23420
rect 27212 23418 27236 23420
rect 26972 23366 26982 23418
rect 27226 23366 27236 23418
rect 26972 23364 26996 23366
rect 27052 23364 27076 23366
rect 27132 23364 27156 23366
rect 27212 23364 27236 23366
rect 26916 23355 27292 23364
rect 11656 22876 12032 22885
rect 11712 22874 11736 22876
rect 11792 22874 11816 22876
rect 11872 22874 11896 22876
rect 11952 22874 11976 22876
rect 11712 22822 11722 22874
rect 11966 22822 11976 22874
rect 11712 22820 11736 22822
rect 11792 22820 11816 22822
rect 11872 22820 11896 22822
rect 11952 22820 11976 22822
rect 11656 22811 12032 22820
rect 19656 22876 20032 22885
rect 19712 22874 19736 22876
rect 19792 22874 19816 22876
rect 19872 22874 19896 22876
rect 19952 22874 19976 22876
rect 19712 22822 19722 22874
rect 19966 22822 19976 22874
rect 19712 22820 19736 22822
rect 19792 22820 19816 22822
rect 19872 22820 19896 22822
rect 19952 22820 19976 22822
rect 19656 22811 20032 22820
rect 27656 22876 28032 22885
rect 27712 22874 27736 22876
rect 27792 22874 27816 22876
rect 27872 22874 27896 22876
rect 27952 22874 27976 22876
rect 27712 22822 27722 22874
rect 27966 22822 27976 22874
rect 27712 22820 27736 22822
rect 27792 22820 27816 22822
rect 27872 22820 27896 22822
rect 27952 22820 27976 22822
rect 27656 22811 28032 22820
rect 28080 22636 28132 22642
rect 28080 22578 28132 22584
rect 10916 22332 11292 22341
rect 10972 22330 10996 22332
rect 11052 22330 11076 22332
rect 11132 22330 11156 22332
rect 11212 22330 11236 22332
rect 10972 22278 10982 22330
rect 11226 22278 11236 22330
rect 10972 22276 10996 22278
rect 11052 22276 11076 22278
rect 11132 22276 11156 22278
rect 11212 22276 11236 22278
rect 10916 22267 11292 22276
rect 18916 22332 19292 22341
rect 18972 22330 18996 22332
rect 19052 22330 19076 22332
rect 19132 22330 19156 22332
rect 19212 22330 19236 22332
rect 18972 22278 18982 22330
rect 19226 22278 19236 22330
rect 18972 22276 18996 22278
rect 19052 22276 19076 22278
rect 19132 22276 19156 22278
rect 19212 22276 19236 22278
rect 18916 22267 19292 22276
rect 26916 22332 27292 22341
rect 26972 22330 26996 22332
rect 27052 22330 27076 22332
rect 27132 22330 27156 22332
rect 27212 22330 27236 22332
rect 26972 22278 26982 22330
rect 27226 22278 27236 22330
rect 26972 22276 26996 22278
rect 27052 22276 27076 22278
rect 27132 22276 27156 22278
rect 27212 22276 27236 22278
rect 26916 22267 27292 22276
rect 9036 22024 9088 22030
rect 9036 21966 9088 21972
rect 8944 21072 8996 21078
rect 8944 21014 8996 21020
rect 8956 20466 8984 21014
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 9048 17270 9076 21966
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 9128 21004 9180 21010
rect 9128 20946 9180 20952
rect 9140 20466 9168 20946
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 9404 19780 9456 19786
rect 9404 19722 9456 19728
rect 9416 19514 9444 19722
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9232 18222 9260 19110
rect 9508 18358 9536 21830
rect 11656 21788 12032 21797
rect 11712 21786 11736 21788
rect 11792 21786 11816 21788
rect 11872 21786 11896 21788
rect 11952 21786 11976 21788
rect 11712 21734 11722 21786
rect 11966 21734 11976 21786
rect 11712 21732 11736 21734
rect 11792 21732 11816 21734
rect 11872 21732 11896 21734
rect 11952 21732 11976 21734
rect 11656 21723 12032 21732
rect 19656 21788 20032 21797
rect 19712 21786 19736 21788
rect 19792 21786 19816 21788
rect 19872 21786 19896 21788
rect 19952 21786 19976 21788
rect 19712 21734 19722 21786
rect 19966 21734 19976 21786
rect 19712 21732 19736 21734
rect 19792 21732 19816 21734
rect 19872 21732 19896 21734
rect 19952 21732 19976 21734
rect 19656 21723 20032 21732
rect 27656 21788 28032 21797
rect 27712 21786 27736 21788
rect 27792 21786 27816 21788
rect 27872 21786 27896 21788
rect 27952 21786 27976 21788
rect 27712 21734 27722 21786
rect 27966 21734 27976 21786
rect 27712 21732 27736 21734
rect 27792 21732 27816 21734
rect 27872 21732 27896 21734
rect 27952 21732 27976 21734
rect 27656 21723 28032 21732
rect 10916 21244 11292 21253
rect 10972 21242 10996 21244
rect 11052 21242 11076 21244
rect 11132 21242 11156 21244
rect 11212 21242 11236 21244
rect 10972 21190 10982 21242
rect 11226 21190 11236 21242
rect 10972 21188 10996 21190
rect 11052 21188 11076 21190
rect 11132 21188 11156 21190
rect 11212 21188 11236 21190
rect 10916 21179 11292 21188
rect 18916 21244 19292 21253
rect 18972 21242 18996 21244
rect 19052 21242 19076 21244
rect 19132 21242 19156 21244
rect 19212 21242 19236 21244
rect 18972 21190 18982 21242
rect 19226 21190 19236 21242
rect 18972 21188 18996 21190
rect 19052 21188 19076 21190
rect 19132 21188 19156 21190
rect 19212 21188 19236 21190
rect 18916 21179 19292 21188
rect 26916 21244 27292 21253
rect 26972 21242 26996 21244
rect 27052 21242 27076 21244
rect 27132 21242 27156 21244
rect 27212 21242 27236 21244
rect 26972 21190 26982 21242
rect 27226 21190 27236 21242
rect 26972 21188 26996 21190
rect 27052 21188 27076 21190
rect 27132 21188 27156 21190
rect 27212 21188 27236 21190
rect 26916 21179 27292 21188
rect 12900 20868 12952 20874
rect 12900 20810 12952 20816
rect 9864 20800 9916 20806
rect 9864 20742 9916 20748
rect 9588 20324 9640 20330
rect 9588 20266 9640 20272
rect 9600 19786 9628 20266
rect 9876 19922 9904 20742
rect 11656 20700 12032 20709
rect 11712 20698 11736 20700
rect 11792 20698 11816 20700
rect 11872 20698 11896 20700
rect 11952 20698 11976 20700
rect 11712 20646 11722 20698
rect 11966 20646 11976 20698
rect 11712 20644 11736 20646
rect 11792 20644 11816 20646
rect 11872 20644 11896 20646
rect 11952 20644 11976 20646
rect 11656 20635 12032 20644
rect 10048 20324 10100 20330
rect 10048 20266 10100 20272
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9588 19780 9640 19786
rect 9588 19722 9640 19728
rect 9784 19514 9812 19790
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9876 19446 9904 19858
rect 10060 19854 10088 20266
rect 10232 20256 10284 20262
rect 10232 20198 10284 20204
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 10048 19848 10100 19854
rect 10048 19790 10100 19796
rect 9864 19440 9916 19446
rect 9864 19382 9916 19388
rect 10152 18358 10180 19994
rect 10244 19854 10272 20198
rect 10916 20156 11292 20165
rect 10972 20154 10996 20156
rect 11052 20154 11076 20156
rect 11132 20154 11156 20156
rect 11212 20154 11236 20156
rect 10972 20102 10982 20154
rect 11226 20102 11236 20154
rect 10972 20100 10996 20102
rect 11052 20100 11076 20102
rect 11132 20100 11156 20102
rect 11212 20100 11236 20102
rect 10916 20091 11292 20100
rect 12440 19916 12492 19922
rect 12440 19858 12492 19864
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 10244 19378 10272 19790
rect 11656 19612 12032 19621
rect 11712 19610 11736 19612
rect 11792 19610 11816 19612
rect 11872 19610 11896 19612
rect 11952 19610 11976 19612
rect 11712 19558 11722 19610
rect 11966 19558 11976 19610
rect 11712 19556 11736 19558
rect 11792 19556 11816 19558
rect 11872 19556 11896 19558
rect 11952 19556 11976 19558
rect 11656 19547 12032 19556
rect 10232 19372 10284 19378
rect 10232 19314 10284 19320
rect 10916 19068 11292 19077
rect 10972 19066 10996 19068
rect 11052 19066 11076 19068
rect 11132 19066 11156 19068
rect 11212 19066 11236 19068
rect 10972 19014 10982 19066
rect 11226 19014 11236 19066
rect 10972 19012 10996 19014
rect 11052 19012 11076 19014
rect 11132 19012 11156 19014
rect 11212 19012 11236 19014
rect 10916 19003 11292 19012
rect 11336 18760 11388 18766
rect 11336 18702 11388 18708
rect 9496 18352 9548 18358
rect 9496 18294 9548 18300
rect 10140 18352 10192 18358
rect 10140 18294 10192 18300
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9588 18284 9640 18290
rect 9864 18284 9916 18290
rect 9640 18244 9864 18272
rect 9588 18226 9640 18232
rect 9864 18226 9916 18232
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 9036 17264 9088 17270
rect 9036 17206 9088 17212
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 9140 16658 9168 16934
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 8864 15638 8892 16050
rect 8852 15632 8904 15638
rect 8852 15574 8904 15580
rect 8956 15570 8984 16050
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 9232 15162 9260 18158
rect 9416 17338 9444 18226
rect 9496 18080 9548 18086
rect 9548 18028 9720 18034
rect 9496 18022 9720 18028
rect 9508 18006 9720 18022
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9600 15706 9628 16050
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9692 15162 9720 18006
rect 10916 17980 11292 17989
rect 10972 17978 10996 17980
rect 11052 17978 11076 17980
rect 11132 17978 11156 17980
rect 11212 17978 11236 17980
rect 10972 17926 10982 17978
rect 11226 17926 11236 17978
rect 10972 17924 10996 17926
rect 11052 17924 11076 17926
rect 11132 17924 11156 17926
rect 11212 17924 11236 17926
rect 10916 17915 11292 17924
rect 9864 17264 9916 17270
rect 9864 17206 9916 17212
rect 9876 16250 9904 17206
rect 10916 16892 11292 16901
rect 10972 16890 10996 16892
rect 11052 16890 11076 16892
rect 11132 16890 11156 16892
rect 11212 16890 11236 16892
rect 10972 16838 10982 16890
rect 11226 16838 11236 16890
rect 10972 16836 10996 16838
rect 11052 16836 11076 16838
rect 11132 16836 11156 16838
rect 11212 16836 11236 16838
rect 10916 16827 11292 16836
rect 11348 16658 11376 18702
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 11656 18524 12032 18533
rect 11712 18522 11736 18524
rect 11792 18522 11816 18524
rect 11872 18522 11896 18524
rect 11952 18522 11976 18524
rect 11712 18470 11722 18522
rect 11966 18470 11976 18522
rect 11712 18468 11736 18470
rect 11792 18468 11816 18470
rect 11872 18468 11896 18470
rect 11952 18468 11976 18470
rect 11656 18459 12032 18468
rect 12084 18426 12112 18566
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 12452 18358 12480 19858
rect 12624 19780 12676 19786
rect 12624 19722 12676 19728
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12544 19514 12572 19654
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 12440 18352 12492 18358
rect 12636 18306 12664 19722
rect 12912 19310 12940 20810
rect 19656 20700 20032 20709
rect 19712 20698 19736 20700
rect 19792 20698 19816 20700
rect 19872 20698 19896 20700
rect 19952 20698 19976 20700
rect 19712 20646 19722 20698
rect 19966 20646 19976 20698
rect 19712 20644 19736 20646
rect 19792 20644 19816 20646
rect 19872 20644 19896 20646
rect 19952 20644 19976 20646
rect 19656 20635 20032 20644
rect 27656 20700 28032 20709
rect 27712 20698 27736 20700
rect 27792 20698 27816 20700
rect 27872 20698 27896 20700
rect 27952 20698 27976 20700
rect 27712 20646 27722 20698
rect 27966 20646 27976 20698
rect 27712 20644 27736 20646
rect 27792 20644 27816 20646
rect 27872 20644 27896 20646
rect 27952 20644 27976 20646
rect 27656 20635 28032 20644
rect 21916 20256 21968 20262
rect 21916 20198 21968 20204
rect 24032 20256 24084 20262
rect 24032 20198 24084 20204
rect 18916 20156 19292 20165
rect 18972 20154 18996 20156
rect 19052 20154 19076 20156
rect 19132 20154 19156 20156
rect 19212 20154 19236 20156
rect 18972 20102 18982 20154
rect 19226 20102 19236 20154
rect 18972 20100 18996 20102
rect 19052 20100 19076 20102
rect 19132 20100 19156 20102
rect 19212 20100 19236 20102
rect 18916 20091 19292 20100
rect 21928 19854 21956 20198
rect 23204 20052 23256 20058
rect 23204 19994 23256 20000
rect 23572 20052 23624 20058
rect 23572 19994 23624 20000
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 23020 19916 23072 19922
rect 23020 19858 23072 19864
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 21916 19848 21968 19854
rect 21916 19790 21968 19796
rect 22192 19848 22244 19854
rect 22192 19790 22244 19796
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 12820 18970 12848 19246
rect 14476 18970 14504 19790
rect 22204 19718 22232 19790
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 18156 19446 18184 19654
rect 18144 19440 18196 19446
rect 18144 19382 18196 19388
rect 18788 19440 18840 19446
rect 18788 19382 18840 19388
rect 15108 19372 15160 19378
rect 15108 19314 15160 19320
rect 15292 19372 15344 19378
rect 15292 19314 15344 19320
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 12808 18964 12860 18970
rect 12728 18924 12808 18952
rect 12728 18426 12756 18924
rect 12808 18906 12860 18912
rect 14464 18964 14516 18970
rect 14516 18924 14596 18952
rect 14464 18906 14516 18912
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12440 18294 12492 18300
rect 12544 18278 12664 18306
rect 12164 18148 12216 18154
rect 12164 18090 12216 18096
rect 11656 17436 12032 17445
rect 11712 17434 11736 17436
rect 11792 17434 11816 17436
rect 11872 17434 11896 17436
rect 11952 17434 11976 17436
rect 11712 17382 11722 17434
rect 11966 17382 11976 17434
rect 11712 17380 11736 17382
rect 11792 17380 11816 17382
rect 11872 17380 11896 17382
rect 11952 17380 11976 17382
rect 11656 17371 12032 17380
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 10140 16176 10192 16182
rect 10140 16118 10192 16124
rect 10152 15706 10180 16118
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10612 15706 10640 15846
rect 10916 15804 11292 15813
rect 10972 15802 10996 15804
rect 11052 15802 11076 15804
rect 11132 15802 11156 15804
rect 11212 15802 11236 15804
rect 10972 15750 10982 15802
rect 11226 15750 11236 15802
rect 10972 15748 10996 15750
rect 11052 15748 11076 15750
rect 11132 15748 11156 15750
rect 11212 15748 11236 15750
rect 10916 15739 11292 15748
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9600 14074 9628 14962
rect 9784 14958 9812 15438
rect 10428 15026 10456 15438
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9864 14884 9916 14890
rect 9864 14826 9916 14832
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9220 14000 9272 14006
rect 9220 13942 9272 13948
rect 9496 14000 9548 14006
rect 9496 13942 9548 13948
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8024 13456 8076 13462
rect 8024 13398 8076 13404
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 8404 13326 8432 13670
rect 8956 13530 8984 13806
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7208 12986 7236 13126
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 8404 12918 8432 13262
rect 8392 12912 8444 12918
rect 8392 12854 8444 12860
rect 8864 12850 8892 13262
rect 9232 13190 9260 13942
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 9416 13394 9444 13670
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9508 13326 9536 13942
rect 9876 13326 9904 14826
rect 10060 13870 10088 14962
rect 10916 14716 11292 14725
rect 10972 14714 10996 14716
rect 11052 14714 11076 14716
rect 11132 14714 11156 14716
rect 11212 14714 11236 14716
rect 10972 14662 10982 14714
rect 11226 14662 11236 14714
rect 10972 14660 10996 14662
rect 11052 14660 11076 14662
rect 11132 14660 11156 14662
rect 11212 14660 11236 14662
rect 10916 14651 11292 14660
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 10060 13326 10088 13806
rect 10916 13628 11292 13637
rect 10972 13626 10996 13628
rect 11052 13626 11076 13628
rect 11132 13626 11156 13628
rect 11212 13626 11236 13628
rect 10972 13574 10982 13626
rect 11226 13574 11236 13626
rect 10972 13572 10996 13574
rect 11052 13572 11076 13574
rect 11132 13572 11156 13574
rect 11212 13572 11236 13574
rect 10916 13563 11292 13572
rect 11348 13326 11376 16594
rect 11656 16348 12032 16357
rect 11712 16346 11736 16348
rect 11792 16346 11816 16348
rect 11872 16346 11896 16348
rect 11952 16346 11976 16348
rect 11712 16294 11722 16346
rect 11966 16294 11976 16346
rect 11712 16292 11736 16294
rect 11792 16292 11816 16294
rect 11872 16292 11896 16294
rect 11952 16292 11976 16294
rect 11656 16283 12032 16292
rect 12084 16250 12112 16594
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 11656 15260 12032 15269
rect 11712 15258 11736 15260
rect 11792 15258 11816 15260
rect 11872 15258 11896 15260
rect 11952 15258 11976 15260
rect 11712 15206 11722 15258
rect 11966 15206 11976 15258
rect 11712 15204 11736 15206
rect 11792 15204 11816 15206
rect 11872 15204 11896 15206
rect 11952 15204 11976 15206
rect 11656 15195 12032 15204
rect 11656 14172 12032 14181
rect 11712 14170 11736 14172
rect 11792 14170 11816 14172
rect 11872 14170 11896 14172
rect 11952 14170 11976 14172
rect 11712 14118 11722 14170
rect 11966 14118 11976 14170
rect 11712 14116 11736 14118
rect 11792 14116 11816 14118
rect 11872 14116 11896 14118
rect 11952 14116 11976 14118
rect 11656 14107 12032 14116
rect 12176 14074 12204 18090
rect 12544 16454 12572 18278
rect 12820 18272 12848 18702
rect 14200 18290 14228 18770
rect 12728 18244 12848 18272
rect 14188 18284 14240 18290
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12544 16250 12572 16390
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12544 15706 12572 15982
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12636 15162 12664 18158
rect 12728 16794 12756 18244
rect 14188 18226 14240 18232
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14476 17882 14504 18158
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14568 17678 14596 18924
rect 15120 18426 15148 19314
rect 15108 18420 15160 18426
rect 15108 18362 15160 18368
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12728 16590 12756 16730
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12176 13802 12204 14010
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12164 13796 12216 13802
rect 12164 13738 12216 13744
rect 12072 13728 12124 13734
rect 12072 13670 12124 13676
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9232 12986 9260 13126
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 11348 12850 11376 13262
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 10916 12540 11292 12549
rect 10972 12538 10996 12540
rect 11052 12538 11076 12540
rect 11132 12538 11156 12540
rect 11212 12538 11236 12540
rect 10972 12486 10982 12538
rect 11226 12486 11236 12538
rect 10972 12484 10996 12486
rect 11052 12484 11076 12486
rect 11132 12484 11156 12486
rect 11212 12484 11236 12486
rect 10916 12475 11292 12484
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 7288 10736 7340 10742
rect 7288 10678 7340 10684
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 6380 10130 6408 10542
rect 7116 10266 7144 10542
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5460 9178 5488 9454
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 4436 8016 4488 8022
rect 4436 7958 4488 7964
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3656 7644 4032 7653
rect 3712 7642 3736 7644
rect 3792 7642 3816 7644
rect 3872 7642 3896 7644
rect 3952 7642 3976 7644
rect 3712 7590 3722 7642
rect 3966 7590 3976 7642
rect 3712 7588 3736 7590
rect 3792 7588 3816 7590
rect 3872 7588 3896 7590
rect 3952 7588 3976 7590
rect 3656 7579 4032 7588
rect 4080 7546 4108 7822
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3608 7472 3660 7478
rect 4172 7426 4200 7686
rect 3608 7414 3660 7420
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3620 6882 3648 7414
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3528 6854 3648 6882
rect 4080 7398 4200 7426
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3436 5098 3464 6666
rect 3528 5352 3556 6854
rect 3656 6556 4032 6565
rect 3712 6554 3736 6556
rect 3792 6554 3816 6556
rect 3872 6554 3896 6556
rect 3952 6554 3976 6556
rect 3712 6502 3722 6554
rect 3966 6502 3976 6554
rect 3712 6500 3736 6502
rect 3792 6500 3816 6502
rect 3872 6500 3896 6502
rect 3952 6500 3976 6502
rect 3656 6491 4032 6500
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3620 5914 3648 6190
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3712 5710 3740 6054
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3656 5468 4032 5477
rect 3712 5466 3736 5468
rect 3792 5466 3816 5468
rect 3872 5466 3896 5468
rect 3952 5466 3976 5468
rect 3712 5414 3722 5466
rect 3966 5414 3976 5466
rect 3712 5412 3736 5414
rect 3792 5412 3816 5414
rect 3872 5412 3896 5414
rect 3952 5412 3976 5414
rect 3656 5403 4032 5412
rect 3700 5364 3752 5370
rect 3528 5324 3700 5352
rect 3700 5306 3752 5312
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3424 5092 3476 5098
rect 3424 5034 3476 5040
rect 3528 4758 3556 5102
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3516 4752 3568 4758
rect 3516 4694 3568 4700
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 2916 3836 3292 3845
rect 2972 3834 2996 3836
rect 3052 3834 3076 3836
rect 3132 3834 3156 3836
rect 3212 3834 3236 3836
rect 2972 3782 2982 3834
rect 3226 3782 3236 3834
rect 2972 3780 2996 3782
rect 3052 3780 3076 3782
rect 3132 3780 3156 3782
rect 3212 3780 3236 3782
rect 2916 3771 3292 3780
rect 3344 3602 3372 4626
rect 3620 4622 3648 4966
rect 4080 4826 4108 7398
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4632 7002 4660 7278
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4724 5302 4752 8842
rect 5460 6866 5488 9114
rect 6288 9042 6316 9930
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6748 9654 6776 9862
rect 7024 9722 7052 10202
rect 7300 9994 7328 10678
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5552 5914 5580 6598
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 5000 5234 5028 5510
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 4264 4826 4292 5170
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3656 4380 4032 4389
rect 3712 4378 3736 4380
rect 3792 4378 3816 4380
rect 3872 4378 3896 4380
rect 3952 4378 3976 4380
rect 3712 4326 3722 4378
rect 3966 4326 3976 4378
rect 3712 4324 3736 4326
rect 3792 4324 3816 4326
rect 3872 4324 3896 4326
rect 3952 4324 3976 4326
rect 3656 4315 4032 4324
rect 4632 4146 4660 4966
rect 4724 4690 4752 4966
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 5000 4282 5028 5170
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 5184 4214 5212 5510
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 5184 3738 5212 4150
rect 5368 4010 5396 5102
rect 5644 4486 5672 7414
rect 6104 7206 6132 8774
rect 6656 8634 6684 9454
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6932 8242 6960 8298
rect 6840 8214 6960 8242
rect 6736 7812 6788 7818
rect 6736 7754 6788 7760
rect 6748 7546 6776 7754
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6012 5914 6040 7142
rect 6104 6798 6132 7142
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6182 6216 6238 6225
rect 6182 6151 6184 6160
rect 6236 6151 6238 6160
rect 6184 6122 6236 6128
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 6092 5840 6144 5846
rect 6092 5782 6144 5788
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5736 5574 5764 5714
rect 6104 5642 6132 5782
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5736 5030 5764 5510
rect 6196 5302 6224 6122
rect 6184 5296 6236 5302
rect 6184 5238 6236 5244
rect 6840 5030 6868 8214
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 6866 6960 7686
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6932 6390 6960 6802
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6932 4690 6960 6326
rect 7116 6186 7144 7890
rect 7208 6390 7236 8366
rect 7300 7818 7328 9930
rect 7576 9178 7604 10066
rect 7668 9586 7696 10066
rect 8128 9994 8156 10406
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7668 8922 7696 9522
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7852 9042 7880 9318
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7668 8894 7880 8922
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7668 8566 7696 8774
rect 7760 8634 7788 8774
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7760 8090 7788 8570
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 7104 6180 7156 6186
rect 7104 6122 7156 6128
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5460 4282 5488 4422
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 3656 3292 4032 3301
rect 3712 3290 3736 3292
rect 3792 3290 3816 3292
rect 3872 3290 3896 3292
rect 3952 3290 3976 3292
rect 3712 3238 3722 3290
rect 3966 3238 3976 3290
rect 3712 3236 3736 3238
rect 3792 3236 3816 3238
rect 3872 3236 3896 3238
rect 3952 3236 3976 3238
rect 3656 3227 4032 3236
rect 4080 3194 4108 3402
rect 5184 3194 5212 3674
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5368 2990 5396 3946
rect 5644 3466 5672 4422
rect 6932 4162 6960 4626
rect 7196 4548 7248 4554
rect 7196 4490 7248 4496
rect 7208 4282 7236 4490
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 6840 4134 6960 4162
rect 6840 3602 6868 4134
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 7300 3466 7328 7754
rect 7760 7546 7788 8026
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7852 7342 7880 8894
rect 8864 7546 8892 11834
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9416 11150 9444 11630
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9416 11014 9444 11086
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8956 9926 8984 10542
rect 9416 10062 9444 10950
rect 9692 10810 9720 11630
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 10704 10742 10732 12174
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11164 11558 11192 12038
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 10796 10810 10824 11494
rect 10916 11452 11292 11461
rect 10972 11450 10996 11452
rect 11052 11450 11076 11452
rect 11132 11450 11156 11452
rect 11212 11450 11236 11452
rect 10972 11398 10982 11450
rect 11226 11398 11236 11450
rect 10972 11396 10996 11398
rect 11052 11396 11076 11398
rect 11132 11396 11156 11398
rect 11212 11396 11236 11398
rect 10916 11387 11292 11396
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 9588 10736 9640 10742
rect 9588 10678 9640 10684
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 9416 9042 9444 9998
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7668 6458 7696 7278
rect 8864 6730 8892 7482
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8852 6724 8904 6730
rect 8852 6666 8904 6672
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 8036 6254 8064 6598
rect 8772 6458 8800 6666
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8036 5778 8064 6190
rect 8128 5778 8156 6326
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8220 5710 8248 6258
rect 8864 6118 8892 6666
rect 9600 6390 9628 10678
rect 11348 10674 11376 12786
rect 11440 12646 11468 12922
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11440 11830 11468 12582
rect 11428 11824 11480 11830
rect 11428 11766 11480 11772
rect 11532 11642 11560 13194
rect 11656 13084 12032 13093
rect 11712 13082 11736 13084
rect 11792 13082 11816 13084
rect 11872 13082 11896 13084
rect 11952 13082 11976 13084
rect 11712 13030 11722 13082
rect 11966 13030 11976 13082
rect 11712 13028 11736 13030
rect 11792 13028 11816 13030
rect 11872 13028 11896 13030
rect 11952 13028 11976 13030
rect 11656 13019 12032 13028
rect 12084 12918 12112 13670
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 11656 11996 12032 12005
rect 11712 11994 11736 11996
rect 11792 11994 11816 11996
rect 11872 11994 11896 11996
rect 11952 11994 11976 11996
rect 11712 11942 11722 11994
rect 11966 11942 11976 11994
rect 11712 11940 11736 11942
rect 11792 11940 11816 11942
rect 11872 11940 11896 11942
rect 11952 11940 11976 11942
rect 11656 11931 12032 11940
rect 11440 11614 11560 11642
rect 11440 11558 11468 11614
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 11440 11082 11468 11494
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 10916 10364 11292 10373
rect 10972 10362 10996 10364
rect 11052 10362 11076 10364
rect 11132 10362 11156 10364
rect 11212 10362 11236 10364
rect 10972 10310 10982 10362
rect 11226 10310 11236 10362
rect 10972 10308 10996 10310
rect 11052 10308 11076 10310
rect 11132 10308 11156 10310
rect 11212 10308 11236 10310
rect 10916 10299 11292 10308
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 10244 8634 10272 8842
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10324 6724 10376 6730
rect 10324 6666 10376 6672
rect 9588 6384 9640 6390
rect 9588 6326 9640 6332
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 9784 5914 9812 6190
rect 10336 6186 10364 6666
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10324 6180 10376 6186
rect 10324 6122 10376 6128
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8220 4826 8248 5646
rect 9784 5574 9812 5850
rect 10704 5658 10732 6258
rect 10796 6118 10824 10134
rect 10916 9276 11292 9285
rect 10972 9274 10996 9276
rect 11052 9274 11076 9276
rect 11132 9274 11156 9276
rect 11212 9274 11236 9276
rect 10972 9222 10982 9274
rect 11226 9222 11236 9274
rect 10972 9220 10996 9222
rect 11052 9220 11076 9222
rect 11132 9220 11156 9222
rect 11212 9220 11236 9222
rect 10916 9211 11292 9220
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11072 8430 11100 8774
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 11256 8378 11284 8910
rect 11348 8498 11376 8978
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11256 8350 11376 8378
rect 10916 8188 11292 8197
rect 10972 8186 10996 8188
rect 11052 8186 11076 8188
rect 11132 8186 11156 8188
rect 11212 8186 11236 8188
rect 10972 8134 10982 8186
rect 11226 8134 11236 8186
rect 10972 8132 10996 8134
rect 11052 8132 11076 8134
rect 11132 8132 11156 8134
rect 11212 8132 11236 8134
rect 10916 8123 11292 8132
rect 10916 7100 11292 7109
rect 10972 7098 10996 7100
rect 11052 7098 11076 7100
rect 11132 7098 11156 7100
rect 11212 7098 11236 7100
rect 10972 7046 10982 7098
rect 11226 7046 11236 7098
rect 10972 7044 10996 7046
rect 11052 7044 11076 7046
rect 11132 7044 11156 7046
rect 11212 7044 11236 7046
rect 10916 7035 11292 7044
rect 11348 6798 11376 8350
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11348 6186 11376 6598
rect 11440 6458 11468 11018
rect 11656 10908 12032 10917
rect 11712 10906 11736 10908
rect 11792 10906 11816 10908
rect 11872 10906 11896 10908
rect 11952 10906 11976 10908
rect 11712 10854 11722 10906
rect 11966 10854 11976 10906
rect 11712 10852 11736 10854
rect 11792 10852 11816 10854
rect 11872 10852 11896 10854
rect 11952 10852 11976 10854
rect 11656 10843 12032 10852
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11808 10266 11836 10542
rect 12176 10470 12204 13738
rect 12544 12442 12572 13806
rect 12728 12986 12756 16526
rect 14752 16182 14780 17682
rect 15120 17610 15148 18362
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 14556 16176 14608 16182
rect 14556 16118 14608 16124
rect 14740 16176 14792 16182
rect 14740 16118 14792 16124
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13556 15502 13584 15846
rect 14568 15638 14596 16118
rect 14556 15632 14608 15638
rect 14556 15574 14608 15580
rect 14752 15570 14780 16118
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 15028 15706 15056 15982
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 15212 15570 15240 15846
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 14740 15564 14792 15570
rect 14740 15506 14792 15512
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13096 15162 13124 15438
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 13280 14958 13308 15302
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13280 13938 13308 14894
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13280 12986 13308 13874
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 13372 12306 13400 14894
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 13464 12850 13492 13126
rect 13648 12850 13676 15506
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 13820 13252 13872 13258
rect 13820 13194 13872 13200
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 12544 12170 12572 12242
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 12440 10736 12492 10742
rect 12440 10678 12492 10684
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 11796 10260 11848 10266
rect 12176 10248 12204 10406
rect 12176 10220 12296 10248
rect 11796 10202 11848 10208
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 11656 9820 12032 9829
rect 11712 9818 11736 9820
rect 11792 9818 11816 9820
rect 11872 9818 11896 9820
rect 11952 9818 11976 9820
rect 11712 9766 11722 9818
rect 11966 9766 11976 9818
rect 11712 9764 11736 9766
rect 11792 9764 11816 9766
rect 11872 9764 11896 9766
rect 11952 9764 11976 9766
rect 11656 9755 12032 9764
rect 12084 9722 12112 9862
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11532 8838 11560 9522
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11992 9178 12020 9454
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11992 9042 12020 9114
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 11532 8634 11560 8774
rect 11656 8732 12032 8741
rect 11712 8730 11736 8732
rect 11792 8730 11816 8732
rect 11872 8730 11896 8732
rect 11952 8730 11976 8732
rect 11712 8678 11722 8730
rect 11966 8678 11976 8730
rect 11712 8676 11736 8678
rect 11792 8676 11816 8678
rect 11872 8676 11896 8678
rect 11952 8676 11976 8678
rect 11656 8667 12032 8676
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 12176 8430 12204 10066
rect 12164 8424 12216 8430
rect 12084 8372 12164 8378
rect 12084 8366 12216 8372
rect 12084 8350 12204 8366
rect 11656 7644 12032 7653
rect 11712 7642 11736 7644
rect 11792 7642 11816 7644
rect 11872 7642 11896 7644
rect 11952 7642 11976 7644
rect 11712 7590 11722 7642
rect 11966 7590 11976 7642
rect 11712 7588 11736 7590
rect 11792 7588 11816 7590
rect 11872 7588 11896 7590
rect 11952 7588 11976 7590
rect 11656 7579 12032 7588
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10796 5778 10824 6054
rect 10916 6012 11292 6021
rect 10972 6010 10996 6012
rect 11052 6010 11076 6012
rect 11132 6010 11156 6012
rect 11212 6010 11236 6012
rect 10972 5958 10982 6010
rect 11226 5958 11236 6010
rect 10972 5956 10996 5958
rect 11052 5956 11076 5958
rect 11132 5956 11156 5958
rect 11212 5956 11236 5958
rect 10916 5947 11292 5956
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 11348 5710 11376 6122
rect 11336 5704 11388 5710
rect 10704 5630 11008 5658
rect 11336 5646 11388 5652
rect 10980 5574 11008 5630
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 11336 5568 11388 5574
rect 11336 5510 11388 5516
rect 10888 5370 10916 5510
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8220 4282 8248 4762
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 7288 3460 7340 3466
rect 7288 3402 7340 3408
rect 6840 3194 6868 3402
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 8128 2990 8156 4014
rect 8312 3602 8340 4966
rect 10916 4924 11292 4933
rect 10972 4922 10996 4924
rect 11052 4922 11076 4924
rect 11132 4922 11156 4924
rect 11212 4922 11236 4924
rect 10972 4870 10982 4922
rect 11226 4870 11236 4922
rect 10972 4868 10996 4870
rect 11052 4868 11076 4870
rect 11132 4868 11156 4870
rect 11212 4868 11236 4870
rect 10916 4859 11292 4868
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9312 4208 9364 4214
rect 9312 4150 9364 4156
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8772 3466 8800 4014
rect 8956 3738 8984 4014
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9324 3534 9352 4150
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8312 3194 8340 3334
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8956 3126 8984 3334
rect 9324 3194 9352 3470
rect 9692 3466 9720 4626
rect 11348 4214 11376 5510
rect 11532 4690 11560 6666
rect 11656 6556 12032 6565
rect 11712 6554 11736 6556
rect 11792 6554 11816 6556
rect 11872 6554 11896 6556
rect 11952 6554 11976 6556
rect 11712 6502 11722 6554
rect 11966 6502 11976 6554
rect 11712 6500 11736 6502
rect 11792 6500 11816 6502
rect 11872 6500 11896 6502
rect 11952 6500 11976 6502
rect 11656 6491 12032 6500
rect 11612 5840 11664 5846
rect 11612 5782 11664 5788
rect 11624 5574 11652 5782
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11656 5468 12032 5477
rect 11712 5466 11736 5468
rect 11792 5466 11816 5468
rect 11872 5466 11896 5468
rect 11952 5466 11976 5468
rect 11712 5414 11722 5466
rect 11966 5414 11976 5466
rect 11712 5412 11736 5414
rect 11792 5412 11816 5414
rect 11872 5412 11896 5414
rect 11952 5412 11976 5414
rect 11656 5403 12032 5412
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11656 4380 12032 4389
rect 11712 4378 11736 4380
rect 11792 4378 11816 4380
rect 11872 4378 11896 4380
rect 11952 4378 11976 4380
rect 11712 4326 11722 4378
rect 11966 4326 11976 4378
rect 11712 4324 11736 4326
rect 11792 4324 11816 4326
rect 11872 4324 11896 4326
rect 11952 4324 11976 4326
rect 11656 4315 12032 4324
rect 11336 4208 11388 4214
rect 11336 4150 11388 4156
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9692 3126 9720 3402
rect 10796 3194 10824 4014
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 10916 3836 11292 3845
rect 10972 3834 10996 3836
rect 11052 3834 11076 3836
rect 11132 3834 11156 3836
rect 11212 3834 11236 3836
rect 10972 3782 10982 3834
rect 11226 3782 11236 3834
rect 10972 3780 10996 3782
rect 11052 3780 11076 3782
rect 11132 3780 11156 3782
rect 11212 3780 11236 3782
rect 10916 3771 11292 3780
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 11440 3126 11468 3878
rect 11808 3738 11836 4150
rect 12084 4078 12112 8350
rect 12164 5908 12216 5914
rect 12268 5896 12296 10220
rect 12452 8974 12480 10678
rect 13280 10470 13308 12038
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13280 10062 13308 10406
rect 13464 10198 13492 12786
rect 13648 12442 13676 12786
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13648 12170 13676 12378
rect 13832 12374 13860 13194
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13636 12164 13688 12170
rect 13636 12106 13688 12112
rect 13740 11286 13768 12242
rect 14384 11354 14412 15302
rect 14752 14090 14780 15506
rect 15212 15178 15240 15506
rect 15120 15150 15240 15178
rect 14752 14062 14872 14090
rect 15120 14074 15148 15150
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15212 14278 15240 14418
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 14740 14000 14792 14006
rect 14740 13942 14792 13948
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14476 13530 14504 13806
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14752 12306 14780 13942
rect 14844 13462 14872 14062
rect 15108 14068 15160 14074
rect 15108 14010 15160 14016
rect 14832 13456 14884 13462
rect 14832 13398 14884 13404
rect 14844 12986 14872 13398
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 15028 11218 15056 11698
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 15212 11150 15240 14214
rect 15304 12918 15332 19314
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15488 17746 15516 19110
rect 16868 18766 16896 19314
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 15936 18692 15988 18698
rect 15936 18634 15988 18640
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15580 18290 15608 18566
rect 15568 18284 15620 18290
rect 15568 18226 15620 18232
rect 15948 17882 15976 18634
rect 16488 18284 16540 18290
rect 16488 18226 16540 18232
rect 16500 17882 16528 18226
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 16212 17604 16264 17610
rect 16212 17546 16264 17552
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15580 13938 15608 15574
rect 15856 14618 15884 17478
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 15304 11898 15332 12106
rect 15580 11898 15608 13874
rect 15948 13870 15976 14282
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 15948 13326 15976 13806
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15856 11694 15884 12922
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 15764 11354 15792 11630
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 16040 11150 16068 16186
rect 16224 14618 16252 17546
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 16132 13870 16160 14418
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 16132 11762 16160 13806
rect 16500 12170 16528 17818
rect 16868 17134 16896 18702
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16868 16658 16896 17070
rect 17696 16794 17724 17478
rect 18248 17202 18276 18022
rect 18696 17604 18748 17610
rect 18696 17546 18748 17552
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18616 17338 18644 17478
rect 18604 17332 18656 17338
rect 18604 17274 18656 17280
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 17684 16788 17736 16794
rect 17684 16730 17736 16736
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17328 15570 17356 16594
rect 18248 16522 18276 17138
rect 18708 16794 18736 17546
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18236 16516 18288 16522
rect 18236 16458 18288 16464
rect 18708 16114 18736 16730
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18800 15994 18828 19382
rect 19352 19174 19380 19654
rect 19656 19612 20032 19621
rect 19712 19610 19736 19612
rect 19792 19610 19816 19612
rect 19872 19610 19896 19612
rect 19952 19610 19976 19612
rect 19712 19558 19722 19610
rect 19966 19558 19976 19610
rect 19712 19556 19736 19558
rect 19792 19556 19816 19558
rect 19872 19556 19896 19558
rect 19952 19556 19976 19558
rect 19656 19547 20032 19556
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 18916 19068 19292 19077
rect 18972 19066 18996 19068
rect 19052 19066 19076 19068
rect 19132 19066 19156 19068
rect 19212 19066 19236 19068
rect 18972 19014 18982 19066
rect 19226 19014 19236 19066
rect 18972 19012 18996 19014
rect 19052 19012 19076 19014
rect 19132 19012 19156 19014
rect 19212 19012 19236 19014
rect 18916 19003 19292 19012
rect 19656 18524 20032 18533
rect 19712 18522 19736 18524
rect 19792 18522 19816 18524
rect 19872 18522 19896 18524
rect 19952 18522 19976 18524
rect 19712 18470 19722 18522
rect 19966 18470 19976 18522
rect 19712 18468 19736 18470
rect 19792 18468 19816 18470
rect 19872 18468 19896 18470
rect 19952 18468 19976 18470
rect 19656 18459 20032 18468
rect 18916 17980 19292 17989
rect 18972 17978 18996 17980
rect 19052 17978 19076 17980
rect 19132 17978 19156 17980
rect 19212 17978 19236 17980
rect 18972 17926 18982 17978
rect 19226 17926 19236 17978
rect 18972 17924 18996 17926
rect 19052 17924 19076 17926
rect 19132 17924 19156 17926
rect 19212 17924 19236 17926
rect 18916 17915 19292 17924
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 18892 17270 18920 17682
rect 19656 17436 20032 17445
rect 19712 17434 19736 17436
rect 19792 17434 19816 17436
rect 19872 17434 19896 17436
rect 19952 17434 19976 17436
rect 19712 17382 19722 17434
rect 19966 17382 19976 17434
rect 19712 17380 19736 17382
rect 19792 17380 19816 17382
rect 19872 17380 19896 17382
rect 19952 17380 19976 17382
rect 19656 17371 20032 17380
rect 18880 17264 18932 17270
rect 18880 17206 18932 17212
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 18916 16892 19292 16901
rect 18972 16890 18996 16892
rect 19052 16890 19076 16892
rect 19132 16890 19156 16892
rect 19212 16890 19236 16892
rect 18972 16838 18982 16890
rect 19226 16838 19236 16890
rect 18972 16836 18996 16838
rect 19052 16836 19076 16838
rect 19132 16836 19156 16838
rect 19212 16836 19236 16838
rect 18916 16827 19292 16836
rect 19904 16590 19932 17070
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 19656 16348 20032 16357
rect 19712 16346 19736 16348
rect 19792 16346 19816 16348
rect 19872 16346 19896 16348
rect 19952 16346 19976 16348
rect 19712 16294 19722 16346
rect 19966 16294 19976 16346
rect 19712 16292 19736 16294
rect 19792 16292 19816 16294
rect 19872 16292 19896 16294
rect 19952 16292 19976 16294
rect 19656 16283 20032 16292
rect 18708 15966 18828 15994
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 17328 14482 17356 15506
rect 18420 15088 18472 15094
rect 18420 15030 18472 15036
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16592 12434 16620 14214
rect 17328 13938 17356 14418
rect 17972 14006 18000 14758
rect 17960 14000 18012 14006
rect 17960 13942 18012 13948
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 16948 12912 17000 12918
rect 16948 12854 17000 12860
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16592 12406 16712 12434
rect 16212 12164 16264 12170
rect 16212 12106 16264 12112
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16224 11898 16252 12106
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16500 11762 16528 12106
rect 16684 12102 16712 12406
rect 16776 12238 16804 12582
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16684 11830 16712 12038
rect 16672 11824 16724 11830
rect 16672 11766 16724 11772
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16672 11688 16724 11694
rect 16500 11636 16672 11642
rect 16500 11630 16724 11636
rect 16500 11614 16712 11630
rect 16500 11150 16528 11614
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 14004 11076 14056 11082
rect 14004 11018 14056 11024
rect 14280 11076 14332 11082
rect 14280 11018 14332 11024
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 13452 10192 13504 10198
rect 13452 10134 13504 10140
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12216 5868 12296 5896
rect 12164 5850 12216 5856
rect 12544 4826 12572 9386
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 12808 6724 12860 6730
rect 12808 6666 12860 6672
rect 13728 6724 13780 6730
rect 13728 6666 13780 6672
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12728 5710 12756 6054
rect 12820 5914 12848 6666
rect 13740 6254 13768 6666
rect 13832 6322 13860 6802
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12164 4208 12216 4214
rect 12164 4150 12216 4156
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11900 3602 11928 3878
rect 12176 3738 12204 4150
rect 12544 4146 12572 4762
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 12820 3602 12848 3878
rect 13832 3602 13860 6258
rect 13924 5710 13952 6258
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13924 4554 13952 5646
rect 14016 5302 14044 11018
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14108 10266 14136 10542
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14200 9178 14228 9454
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 14108 6866 14136 8910
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 6322 14136 6598
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 14096 5840 14148 5846
rect 14096 5782 14148 5788
rect 14004 5296 14056 5302
rect 14004 5238 14056 5244
rect 13912 4548 13964 4554
rect 13912 4490 13964 4496
rect 13924 4078 13952 4490
rect 13912 4072 13964 4078
rect 13912 4014 13964 4020
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 11428 3120 11480 3126
rect 11428 3062 11480 3068
rect 11532 2990 11560 3538
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 11656 3292 12032 3301
rect 11712 3290 11736 3292
rect 11792 3290 11816 3292
rect 11872 3290 11896 3292
rect 11952 3290 11976 3292
rect 11712 3238 11722 3290
rect 11966 3238 11976 3290
rect 11712 3236 11736 3238
rect 11792 3236 11816 3238
rect 11872 3236 11896 3238
rect 11952 3236 11976 3238
rect 11656 3227 12032 3236
rect 12176 3058 12204 3470
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12636 3194 12664 3334
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12728 3126 12756 3538
rect 12716 3120 12768 3126
rect 12716 3062 12768 3068
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 5356 2984 5408 2990
rect 5356 2926 5408 2932
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 14108 2922 14136 5782
rect 14200 5642 14228 7142
rect 14292 6225 14320 11018
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15304 10606 15332 10950
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15304 10062 15332 10542
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15396 9586 15424 11018
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14384 9042 14412 9318
rect 14372 9036 14424 9042
rect 14372 8978 14424 8984
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14568 7410 14596 8230
rect 14844 7478 14872 9386
rect 15384 8900 15436 8906
rect 15384 8842 15436 8848
rect 15396 7546 15424 8842
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 14832 7472 14884 7478
rect 14832 7414 14884 7420
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14372 6724 14424 6730
rect 14372 6666 14424 6672
rect 14384 6458 14412 6666
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14752 6458 14780 6598
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14278 6216 14334 6225
rect 14278 6151 14334 6160
rect 14752 5846 14780 6394
rect 14844 6254 14872 7414
rect 15396 6730 15424 7482
rect 15580 7410 15608 11086
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 15856 9178 15884 9522
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 16776 8294 16804 12174
rect 16960 12170 16988 12854
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16960 11762 16988 12106
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 17604 11218 17632 11494
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17328 9586 17356 11086
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 18064 10742 18092 11018
rect 18052 10736 18104 10742
rect 18052 10678 18104 10684
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17328 8634 17356 9522
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 17328 7954 17356 8570
rect 17880 8022 17908 10066
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17040 7812 17092 7818
rect 17040 7754 17092 7760
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16960 7410 16988 7686
rect 17052 7546 17080 7754
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 14844 5846 14872 6190
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 14832 5840 14884 5846
rect 14832 5782 14884 5788
rect 14188 5636 14240 5642
rect 14188 5578 14240 5584
rect 14844 4690 14872 5782
rect 15396 5370 15424 6666
rect 15580 5574 15608 7346
rect 16960 6458 16988 7346
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16684 5778 16712 6054
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 16960 5710 16988 6394
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 17052 5642 17080 6258
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17040 5636 17092 5642
rect 17040 5578 17092 5584
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 16028 5568 16080 5574
rect 16028 5510 16080 5516
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 14832 4684 14884 4690
rect 14832 4626 14884 4632
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 14384 3602 14412 4422
rect 14752 3738 14780 4422
rect 15396 4214 15424 5306
rect 16040 4622 16068 5510
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 15660 4480 15712 4486
rect 15660 4422 15712 4428
rect 15672 4214 15700 4422
rect 15384 4208 15436 4214
rect 15384 4150 15436 4156
rect 15660 4208 15712 4214
rect 15660 4150 15712 4156
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 15396 3516 15424 4150
rect 15476 3528 15528 3534
rect 15396 3488 15476 3516
rect 15476 3470 15528 3476
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 16316 3194 16344 3334
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 17144 2990 17172 3334
rect 17236 2990 17264 5782
rect 17328 5234 17356 7890
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 17512 7478 17540 7754
rect 17500 7472 17552 7478
rect 17500 7414 17552 7420
rect 17880 7342 17908 7958
rect 17972 7886 18000 10610
rect 18064 9722 18092 10678
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 18064 8498 18092 9658
rect 18156 9654 18184 9862
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 18064 8090 18092 8434
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17972 7274 18000 7822
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17972 5914 18000 7210
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 18432 5658 18460 15030
rect 18708 14414 18736 15966
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 18800 15162 18828 15846
rect 18916 15804 19292 15813
rect 18972 15802 18996 15804
rect 19052 15802 19076 15804
rect 19132 15802 19156 15804
rect 19212 15802 19236 15804
rect 18972 15750 18982 15802
rect 19226 15750 19236 15802
rect 18972 15748 18996 15750
rect 19052 15748 19076 15750
rect 19132 15748 19156 15750
rect 19212 15748 19236 15750
rect 18916 15739 19292 15748
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18696 14408 18748 14414
rect 18524 14356 18696 14362
rect 18524 14350 18748 14356
rect 18524 14334 18736 14350
rect 18524 14006 18552 14334
rect 18800 14074 18828 14962
rect 18916 14716 19292 14725
rect 18972 14714 18996 14716
rect 19052 14714 19076 14716
rect 19132 14714 19156 14716
rect 19212 14714 19236 14716
rect 18972 14662 18982 14714
rect 19226 14662 19236 14714
rect 18972 14660 18996 14662
rect 19052 14660 19076 14662
rect 19132 14660 19156 14662
rect 19212 14660 19236 14662
rect 18916 14651 19292 14660
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 18788 14068 18840 14074
rect 18708 14028 18788 14056
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18524 13870 18552 13942
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18708 12918 18736 14028
rect 18788 14010 18840 14016
rect 18892 13716 18920 14214
rect 18800 13688 18920 13716
rect 18800 12986 18828 13688
rect 18916 13628 19292 13637
rect 18972 13626 18996 13628
rect 19052 13626 19076 13628
rect 19132 13626 19156 13628
rect 19212 13626 19236 13628
rect 18972 13574 18982 13626
rect 19226 13574 19236 13626
rect 18972 13572 18996 13574
rect 19052 13572 19076 13574
rect 19132 13572 19156 13574
rect 19212 13572 19236 13574
rect 18916 13563 19292 13572
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18696 12912 18748 12918
rect 18696 12854 18748 12860
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18708 11898 18736 12582
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18800 8514 18828 12718
rect 18916 12540 19292 12549
rect 18972 12538 18996 12540
rect 19052 12538 19076 12540
rect 19132 12538 19156 12540
rect 19212 12538 19236 12540
rect 18972 12486 18982 12538
rect 19226 12486 19236 12538
rect 18972 12484 18996 12486
rect 19052 12484 19076 12486
rect 19132 12484 19156 12486
rect 19212 12484 19236 12486
rect 18916 12475 19292 12484
rect 19352 11626 19380 15438
rect 19656 15260 20032 15269
rect 19712 15258 19736 15260
rect 19792 15258 19816 15260
rect 19872 15258 19896 15260
rect 19952 15258 19976 15260
rect 19712 15206 19722 15258
rect 19966 15206 19976 15258
rect 19712 15204 19736 15206
rect 19792 15204 19816 15206
rect 19872 15204 19896 15206
rect 19952 15204 19976 15206
rect 19656 15195 20032 15204
rect 19616 15020 19668 15026
rect 19616 14962 19668 14968
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 19536 12782 19564 14418
rect 19628 14414 19656 14962
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19656 14172 20032 14181
rect 19712 14170 19736 14172
rect 19792 14170 19816 14172
rect 19872 14170 19896 14172
rect 19952 14170 19976 14172
rect 19712 14118 19722 14170
rect 19966 14118 19976 14170
rect 19712 14116 19736 14118
rect 19792 14116 19816 14118
rect 19872 14116 19896 14118
rect 19952 14116 19976 14118
rect 19656 14107 20032 14116
rect 19656 13084 20032 13093
rect 19712 13082 19736 13084
rect 19792 13082 19816 13084
rect 19872 13082 19896 13084
rect 19952 13082 19976 13084
rect 19712 13030 19722 13082
rect 19966 13030 19976 13082
rect 19712 13028 19736 13030
rect 19792 13028 19816 13030
rect 19872 13028 19896 13030
rect 19952 13028 19976 13030
rect 19656 13019 20032 13028
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19656 11996 20032 12005
rect 19712 11994 19736 11996
rect 19792 11994 19816 11996
rect 19872 11994 19896 11996
rect 19952 11994 19976 11996
rect 19712 11942 19722 11994
rect 19966 11942 19976 11994
rect 19712 11940 19736 11942
rect 19792 11940 19816 11942
rect 19872 11940 19896 11942
rect 19952 11940 19976 11942
rect 19656 11931 20032 11940
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 18916 11452 19292 11461
rect 18972 11450 18996 11452
rect 19052 11450 19076 11452
rect 19132 11450 19156 11452
rect 19212 11450 19236 11452
rect 18972 11398 18982 11450
rect 19226 11398 19236 11450
rect 18972 11396 18996 11398
rect 19052 11396 19076 11398
rect 19132 11396 19156 11398
rect 19212 11396 19236 11398
rect 18916 11387 19292 11396
rect 18916 10364 19292 10373
rect 18972 10362 18996 10364
rect 19052 10362 19076 10364
rect 19132 10362 19156 10364
rect 19212 10362 19236 10364
rect 18972 10310 18982 10362
rect 19226 10310 19236 10362
rect 18972 10308 18996 10310
rect 19052 10308 19076 10310
rect 19132 10308 19156 10310
rect 19212 10308 19236 10310
rect 18916 10299 19292 10308
rect 18916 9276 19292 9285
rect 18972 9274 18996 9276
rect 19052 9274 19076 9276
rect 19132 9274 19156 9276
rect 19212 9274 19236 9276
rect 18972 9222 18982 9274
rect 19226 9222 19236 9274
rect 18972 9220 18996 9222
rect 19052 9220 19076 9222
rect 19132 9220 19156 9222
rect 19212 9220 19236 9222
rect 18916 9211 19292 9220
rect 19352 9178 19380 11562
rect 19444 11354 19472 11698
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19524 11008 19576 11014
rect 19524 10950 19576 10956
rect 19536 10130 19564 10950
rect 19656 10908 20032 10917
rect 19712 10906 19736 10908
rect 19792 10906 19816 10908
rect 19872 10906 19896 10908
rect 19952 10906 19976 10908
rect 19712 10854 19722 10906
rect 19966 10854 19976 10906
rect 19712 10852 19736 10854
rect 19792 10852 19816 10854
rect 19872 10852 19896 10854
rect 19952 10852 19976 10854
rect 19656 10843 20032 10852
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19904 10130 19932 10406
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19892 10124 19944 10130
rect 19892 10066 19944 10072
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19536 9722 19564 9862
rect 19656 9820 20032 9829
rect 19712 9818 19736 9820
rect 19792 9818 19816 9820
rect 19872 9818 19896 9820
rect 19952 9818 19976 9820
rect 19712 9766 19722 9818
rect 19966 9766 19976 9818
rect 19712 9764 19736 9766
rect 19792 9764 19816 9766
rect 19872 9764 19896 9766
rect 19952 9764 19976 9766
rect 19656 9755 20032 9764
rect 19524 9716 19576 9722
rect 19524 9658 19576 9664
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 18708 8486 18828 8514
rect 19352 8548 19380 9114
rect 19432 8560 19484 8566
rect 19352 8520 19432 8548
rect 18708 7954 18736 8486
rect 18788 8424 18840 8430
rect 18788 8366 18840 8372
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18708 7342 18736 7890
rect 18800 7750 18828 8366
rect 18916 8188 19292 8197
rect 18972 8186 18996 8188
rect 19052 8186 19076 8188
rect 19132 8186 19156 8188
rect 19212 8186 19236 8188
rect 18972 8134 18982 8186
rect 19226 8134 19236 8186
rect 18972 8132 18996 8134
rect 19052 8132 19076 8134
rect 19132 8132 19156 8134
rect 19212 8132 19236 8134
rect 18916 8123 19292 8132
rect 19352 8090 19380 8520
rect 19432 8502 19484 8508
rect 19536 8514 19564 9658
rect 19656 8732 20032 8741
rect 19712 8730 19736 8732
rect 19792 8730 19816 8732
rect 19872 8730 19896 8732
rect 19952 8730 19976 8732
rect 19712 8678 19722 8730
rect 19966 8678 19976 8730
rect 19712 8676 19736 8678
rect 19792 8676 19816 8678
rect 19872 8676 19896 8678
rect 19952 8676 19976 8678
rect 19656 8667 20032 8676
rect 19536 8486 19656 8514
rect 19524 8356 19576 8362
rect 19524 8298 19576 8304
rect 19536 8090 19564 8298
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19628 7886 19656 8486
rect 20456 8090 20484 19110
rect 22204 18970 22232 19654
rect 22848 19394 22876 19858
rect 22756 19378 22876 19394
rect 23032 19378 23060 19858
rect 22744 19372 22876 19378
rect 22796 19366 22876 19372
rect 23020 19372 23072 19378
rect 22744 19314 22796 19320
rect 23020 19314 23072 19320
rect 22756 18970 22784 19314
rect 22192 18964 22244 18970
rect 22192 18906 22244 18912
rect 22744 18964 22796 18970
rect 22744 18906 22796 18912
rect 21824 18760 21876 18766
rect 21824 18702 21876 18708
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20812 18080 20864 18086
rect 20812 18022 20864 18028
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 20628 17128 20680 17134
rect 20628 17070 20680 17076
rect 20640 14958 20668 17070
rect 20732 16726 20760 17682
rect 20824 17542 20852 18022
rect 20812 17536 20864 17542
rect 20812 17478 20864 17484
rect 20916 17338 20944 18226
rect 21836 17882 21864 18702
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22112 18442 22140 18566
rect 22020 18426 22140 18442
rect 22020 18420 22152 18426
rect 22020 18414 22100 18420
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 21824 17876 21876 17882
rect 21824 17818 21876 17824
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 21192 17202 21220 17818
rect 21824 17264 21876 17270
rect 21824 17206 21876 17212
rect 21180 17196 21232 17202
rect 21180 17138 21232 17144
rect 21192 16998 21220 17138
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 20720 16720 20772 16726
rect 20720 16662 20772 16668
rect 20732 15366 20760 16662
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 20732 15094 20760 15302
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20640 14278 20668 14894
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 21100 13938 21128 14350
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 21192 12782 21220 14962
rect 21376 14482 21404 15302
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21376 14006 21404 14418
rect 21364 14000 21416 14006
rect 21364 13942 21416 13948
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 20444 8084 20496 8090
rect 20444 8026 20496 8032
rect 20548 8022 20576 12718
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20640 10810 20668 11222
rect 20732 11014 20760 11698
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20732 10742 20760 10950
rect 20720 10736 20772 10742
rect 20720 10678 20772 10684
rect 20824 10606 20852 12378
rect 21836 12170 21864 17206
rect 22020 16658 22048 18414
rect 22100 18362 22152 18368
rect 22388 18290 22416 18566
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 23032 17270 23060 19314
rect 23216 18698 23244 19994
rect 23296 19984 23348 19990
rect 23296 19926 23348 19932
rect 23308 19446 23336 19926
rect 23584 19854 23612 19994
rect 23572 19848 23624 19854
rect 23572 19790 23624 19796
rect 23388 19780 23440 19786
rect 23388 19722 23440 19728
rect 23400 19514 23428 19722
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23388 19508 23440 19514
rect 23388 19450 23440 19456
rect 23296 19440 23348 19446
rect 23296 19382 23348 19388
rect 23400 18970 23428 19450
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 23204 18692 23256 18698
rect 23204 18634 23256 18640
rect 23216 18154 23244 18634
rect 23400 18358 23428 18906
rect 23492 18698 23520 19654
rect 24044 19446 24072 20198
rect 26916 20156 27292 20165
rect 26972 20154 26996 20156
rect 27052 20154 27076 20156
rect 27132 20154 27156 20156
rect 27212 20154 27236 20156
rect 26972 20102 26982 20154
rect 27226 20102 27236 20154
rect 26972 20100 26996 20102
rect 27052 20100 27076 20102
rect 27132 20100 27156 20102
rect 27212 20100 27236 20102
rect 26916 20091 27292 20100
rect 28092 20058 28120 22578
rect 28356 22568 28408 22574
rect 28356 22510 28408 22516
rect 28368 22409 28396 22510
rect 28354 22400 28410 22409
rect 28354 22335 28410 22344
rect 28080 20052 28132 20058
rect 28080 19994 28132 20000
rect 24308 19780 24360 19786
rect 24308 19722 24360 19728
rect 24216 19712 24268 19718
rect 24216 19654 24268 19660
rect 24032 19440 24084 19446
rect 24084 19388 24164 19394
rect 24032 19382 24164 19388
rect 24044 19366 24164 19382
rect 23480 18692 23532 18698
rect 23480 18634 23532 18640
rect 23388 18352 23440 18358
rect 23388 18294 23440 18300
rect 23388 18216 23440 18222
rect 23492 18170 23520 18634
rect 23440 18164 23520 18170
rect 23388 18158 23520 18164
rect 23204 18148 23256 18154
rect 23400 18142 23520 18158
rect 23204 18090 23256 18096
rect 23112 18080 23164 18086
rect 23112 18022 23164 18028
rect 23124 17270 23152 18022
rect 23020 17264 23072 17270
rect 23020 17206 23072 17212
rect 23112 17264 23164 17270
rect 23112 17206 23164 17212
rect 23032 16726 23060 17206
rect 23216 16998 23244 18090
rect 23204 16992 23256 16998
rect 23204 16934 23256 16940
rect 23020 16720 23072 16726
rect 23020 16662 23072 16668
rect 23216 16658 23244 16934
rect 22008 16652 22060 16658
rect 22008 16594 22060 16600
rect 23204 16652 23256 16658
rect 23204 16594 23256 16600
rect 23492 16590 23520 18142
rect 24136 17746 24164 19366
rect 24124 17740 24176 17746
rect 24124 17682 24176 17688
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 24136 16522 24164 17682
rect 24228 17202 24256 19654
rect 24320 18970 24348 19722
rect 27656 19612 28032 19621
rect 27712 19610 27736 19612
rect 27792 19610 27816 19612
rect 27872 19610 27896 19612
rect 27952 19610 27976 19612
rect 27712 19558 27722 19610
rect 27966 19558 27976 19610
rect 27712 19556 27736 19558
rect 27792 19556 27816 19558
rect 27872 19556 27896 19558
rect 27952 19556 27976 19558
rect 27656 19547 28032 19556
rect 26916 19068 27292 19077
rect 26972 19066 26996 19068
rect 27052 19066 27076 19068
rect 27132 19066 27156 19068
rect 27212 19066 27236 19068
rect 26972 19014 26982 19066
rect 27226 19014 27236 19066
rect 26972 19012 26996 19014
rect 27052 19012 27076 19014
rect 27132 19012 27156 19014
rect 27212 19012 27236 19014
rect 26916 19003 27292 19012
rect 24308 18964 24360 18970
rect 24308 18906 24360 18912
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 24492 18692 24544 18698
rect 24492 18634 24544 18640
rect 24504 18426 24532 18634
rect 24492 18420 24544 18426
rect 24492 18362 24544 18368
rect 24216 17196 24268 17202
rect 24216 17138 24268 17144
rect 24124 16516 24176 16522
rect 24124 16458 24176 16464
rect 24228 15094 24256 17138
rect 23480 15088 23532 15094
rect 23480 15030 23532 15036
rect 24216 15088 24268 15094
rect 24216 15030 24268 15036
rect 21916 14816 21968 14822
rect 21916 14758 21968 14764
rect 21928 13870 21956 14758
rect 23204 14476 23256 14482
rect 23204 14418 23256 14424
rect 23112 14272 23164 14278
rect 23112 14214 23164 14220
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 21916 13864 21968 13870
rect 21916 13806 21968 13812
rect 22008 12640 22060 12646
rect 22008 12582 22060 12588
rect 21916 12368 21968 12374
rect 21916 12310 21968 12316
rect 21824 12164 21876 12170
rect 21824 12106 21876 12112
rect 21928 11694 21956 12310
rect 22020 12306 22048 12582
rect 22008 12300 22060 12306
rect 22008 12242 22060 12248
rect 22296 11898 22324 14010
rect 22388 13870 22416 14010
rect 23124 13938 23152 14214
rect 23112 13932 23164 13938
rect 23112 13874 23164 13880
rect 23216 13870 23244 14418
rect 23492 14346 23520 15030
rect 23480 14340 23532 14346
rect 23480 14282 23532 14288
rect 24228 14006 24256 15030
rect 24216 14000 24268 14006
rect 24216 13942 24268 13948
rect 22376 13864 22428 13870
rect 22376 13806 22428 13812
rect 23204 13864 23256 13870
rect 24216 13864 24268 13870
rect 23256 13812 23520 13818
rect 23204 13806 23520 13812
rect 24216 13806 24268 13812
rect 23216 13790 23520 13806
rect 23296 12096 23348 12102
rect 23296 12038 23348 12044
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 23308 11830 23336 12038
rect 23296 11824 23348 11830
rect 23296 11766 23348 11772
rect 21916 11688 21968 11694
rect 21916 11630 21968 11636
rect 22008 11620 22060 11626
rect 22008 11562 22060 11568
rect 22020 11218 22048 11562
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 22008 11212 22060 11218
rect 22008 11154 22060 11160
rect 21640 11076 21692 11082
rect 21640 11018 21692 11024
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 19892 8016 19944 8022
rect 20536 8016 20588 8022
rect 19944 7964 20116 7970
rect 19892 7958 20116 7964
rect 20536 7958 20588 7964
rect 19904 7954 20116 7958
rect 19904 7948 20128 7954
rect 19904 7942 20076 7948
rect 20076 7890 20128 7896
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 19524 7744 19576 7750
rect 19524 7686 19576 7692
rect 18800 7546 18828 7686
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18696 7336 18748 7342
rect 18696 7278 18748 7284
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18524 5778 18552 6598
rect 18708 6254 18736 7278
rect 18916 7100 19292 7109
rect 18972 7098 18996 7100
rect 19052 7098 19076 7100
rect 19132 7098 19156 7100
rect 19212 7098 19236 7100
rect 18972 7046 18982 7098
rect 19226 7046 19236 7098
rect 18972 7044 18996 7046
rect 19052 7044 19076 7046
rect 19132 7044 19156 7046
rect 19212 7044 19236 7046
rect 18916 7035 19292 7044
rect 19536 6866 19564 7686
rect 19656 7644 20032 7653
rect 19712 7642 19736 7644
rect 19792 7642 19816 7644
rect 19872 7642 19896 7644
rect 19952 7642 19976 7644
rect 19712 7590 19722 7642
rect 19966 7590 19976 7642
rect 19712 7588 19736 7590
rect 19792 7588 19816 7590
rect 19872 7588 19896 7590
rect 19952 7588 19976 7590
rect 19656 7579 20032 7588
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18916 6012 19292 6021
rect 18972 6010 18996 6012
rect 19052 6010 19076 6012
rect 19132 6010 19156 6012
rect 19212 6010 19236 6012
rect 18972 5958 18982 6010
rect 19226 5958 19236 6010
rect 18972 5956 18996 5958
rect 19052 5956 19076 5958
rect 19132 5956 19156 5958
rect 19212 5956 19236 5958
rect 18916 5947 19292 5956
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 19352 5710 19380 6734
rect 19628 6730 19656 7346
rect 20548 6866 20576 7958
rect 21284 7750 21312 8910
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19656 6556 20032 6565
rect 19712 6554 19736 6556
rect 19792 6554 19816 6556
rect 19872 6554 19896 6556
rect 19952 6554 19976 6556
rect 19712 6502 19722 6554
rect 19966 6502 19976 6554
rect 19712 6500 19736 6502
rect 19792 6500 19816 6502
rect 19872 6500 19896 6502
rect 19952 6500 19976 6502
rect 19656 6491 20032 6500
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 19340 5704 19392 5710
rect 18432 5630 18552 5658
rect 19340 5646 19392 5652
rect 20916 5642 20944 6394
rect 21284 6390 21312 7686
rect 21652 7478 21680 11018
rect 22020 9518 22048 11154
rect 22112 11082 22140 11494
rect 23492 11286 23520 13790
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 23848 13728 23900 13734
rect 23848 13670 23900 13676
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23584 11898 23612 12038
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 22100 11076 22152 11082
rect 22100 11018 22152 11024
rect 23676 10606 23704 13670
rect 23860 13394 23888 13670
rect 24228 13530 24256 13806
rect 24216 13524 24268 13530
rect 24216 13466 24268 13472
rect 24504 13462 24532 18362
rect 24596 18222 24624 18702
rect 27656 18524 28032 18533
rect 27712 18522 27736 18524
rect 27792 18522 27816 18524
rect 27872 18522 27896 18524
rect 27952 18522 27976 18524
rect 27712 18470 27722 18522
rect 27966 18470 27976 18522
rect 27712 18468 27736 18470
rect 27792 18468 27816 18470
rect 27872 18468 27896 18470
rect 27952 18468 27976 18470
rect 27656 18459 28032 18468
rect 24584 18216 24636 18222
rect 24584 18158 24636 18164
rect 24596 17338 24624 18158
rect 26916 17980 27292 17989
rect 26972 17978 26996 17980
rect 27052 17978 27076 17980
rect 27132 17978 27156 17980
rect 27212 17978 27236 17980
rect 26972 17926 26982 17978
rect 27226 17926 27236 17978
rect 26972 17924 26996 17926
rect 27052 17924 27076 17926
rect 27132 17924 27156 17926
rect 27212 17924 27236 17926
rect 26916 17915 27292 17924
rect 27656 17436 28032 17445
rect 27712 17434 27736 17436
rect 27792 17434 27816 17436
rect 27872 17434 27896 17436
rect 27952 17434 27976 17436
rect 27712 17382 27722 17434
rect 27966 17382 27976 17434
rect 27712 17380 27736 17382
rect 27792 17380 27816 17382
rect 27872 17380 27896 17382
rect 27952 17380 27976 17382
rect 27656 17371 28032 17380
rect 24584 17332 24636 17338
rect 24584 17274 24636 17280
rect 26916 16892 27292 16901
rect 26972 16890 26996 16892
rect 27052 16890 27076 16892
rect 27132 16890 27156 16892
rect 27212 16890 27236 16892
rect 26972 16838 26982 16890
rect 27226 16838 27236 16890
rect 26972 16836 26996 16838
rect 27052 16836 27076 16838
rect 27132 16836 27156 16838
rect 27212 16836 27236 16838
rect 26916 16827 27292 16836
rect 27656 16348 28032 16357
rect 27712 16346 27736 16348
rect 27792 16346 27816 16348
rect 27872 16346 27896 16348
rect 27952 16346 27976 16348
rect 27712 16294 27722 16346
rect 27966 16294 27976 16346
rect 27712 16292 27736 16294
rect 27792 16292 27816 16294
rect 27872 16292 27896 16294
rect 27952 16292 27976 16294
rect 27656 16283 28032 16292
rect 26916 15804 27292 15813
rect 26972 15802 26996 15804
rect 27052 15802 27076 15804
rect 27132 15802 27156 15804
rect 27212 15802 27236 15804
rect 26972 15750 26982 15802
rect 27226 15750 27236 15802
rect 26972 15748 26996 15750
rect 27052 15748 27076 15750
rect 27132 15748 27156 15750
rect 27212 15748 27236 15750
rect 26916 15739 27292 15748
rect 27656 15260 28032 15269
rect 27712 15258 27736 15260
rect 27792 15258 27816 15260
rect 27872 15258 27896 15260
rect 27952 15258 27976 15260
rect 27712 15206 27722 15258
rect 27966 15206 27976 15258
rect 27712 15204 27736 15206
rect 27792 15204 27816 15206
rect 27872 15204 27896 15206
rect 27952 15204 27976 15206
rect 27656 15195 28032 15204
rect 26916 14716 27292 14725
rect 26972 14714 26996 14716
rect 27052 14714 27076 14716
rect 27132 14714 27156 14716
rect 27212 14714 27236 14716
rect 26972 14662 26982 14714
rect 27226 14662 27236 14714
rect 26972 14660 26996 14662
rect 27052 14660 27076 14662
rect 27132 14660 27156 14662
rect 27212 14660 27236 14662
rect 26916 14651 27292 14660
rect 27656 14172 28032 14181
rect 27712 14170 27736 14172
rect 27792 14170 27816 14172
rect 27872 14170 27896 14172
rect 27952 14170 27976 14172
rect 27712 14118 27722 14170
rect 27966 14118 27976 14170
rect 27712 14116 27736 14118
rect 27792 14116 27816 14118
rect 27872 14116 27896 14118
rect 27952 14116 27976 14118
rect 27656 14107 28032 14116
rect 24676 14000 24728 14006
rect 24676 13942 24728 13948
rect 24492 13456 24544 13462
rect 24492 13398 24544 13404
rect 23848 13388 23900 13394
rect 23848 13330 23900 13336
rect 24504 12374 24532 13398
rect 24688 12374 24716 13942
rect 24768 13864 24820 13870
rect 24768 13806 24820 13812
rect 24780 13326 24808 13806
rect 26916 13628 27292 13637
rect 26972 13626 26996 13628
rect 27052 13626 27076 13628
rect 27132 13626 27156 13628
rect 27212 13626 27236 13628
rect 26972 13574 26982 13626
rect 27226 13574 27236 13626
rect 26972 13572 26996 13574
rect 27052 13572 27076 13574
rect 27132 13572 27156 13574
rect 27212 13572 27236 13574
rect 26916 13563 27292 13572
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24492 12368 24544 12374
rect 24676 12368 24728 12374
rect 24492 12310 24544 12316
rect 24596 12316 24676 12322
rect 24596 12310 24728 12316
rect 24596 12294 24716 12310
rect 24596 11830 24624 12294
rect 24780 12186 24808 13262
rect 27656 13084 28032 13093
rect 27712 13082 27736 13084
rect 27792 13082 27816 13084
rect 27872 13082 27896 13084
rect 27952 13082 27976 13084
rect 27712 13030 27722 13082
rect 27966 13030 27976 13082
rect 27712 13028 27736 13030
rect 27792 13028 27816 13030
rect 27872 13028 27896 13030
rect 27952 13028 27976 13030
rect 27656 13019 28032 13028
rect 26916 12540 27292 12549
rect 26972 12538 26996 12540
rect 27052 12538 27076 12540
rect 27132 12538 27156 12540
rect 27212 12538 27236 12540
rect 26972 12486 26982 12538
rect 27226 12486 27236 12538
rect 26972 12484 26996 12486
rect 27052 12484 27076 12486
rect 27132 12484 27156 12486
rect 27212 12484 27236 12486
rect 26916 12475 27292 12484
rect 24688 12158 24808 12186
rect 24584 11824 24636 11830
rect 24584 11766 24636 11772
rect 24584 11280 24636 11286
rect 24584 11222 24636 11228
rect 24400 11008 24452 11014
rect 24400 10950 24452 10956
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 24216 10600 24268 10606
rect 24216 10542 24268 10548
rect 23388 10464 23440 10470
rect 23388 10406 23440 10412
rect 23664 10464 23716 10470
rect 23664 10406 23716 10412
rect 23400 9722 23428 10406
rect 23388 9716 23440 9722
rect 23388 9658 23440 9664
rect 23676 9654 23704 10406
rect 23664 9648 23716 9654
rect 23664 9590 23716 9596
rect 22376 9580 22428 9586
rect 22376 9522 22428 9528
rect 22008 9512 22060 9518
rect 22008 9454 22060 9460
rect 21824 9444 21876 9450
rect 21824 9386 21876 9392
rect 21836 8838 21864 9386
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 21824 8832 21876 8838
rect 21824 8774 21876 8780
rect 21836 8430 21864 8774
rect 22112 8566 22140 9318
rect 22100 8560 22152 8566
rect 22100 8502 22152 8508
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 21836 7886 21864 8366
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 21640 7472 21692 7478
rect 21640 7414 21692 7420
rect 21364 7336 21416 7342
rect 21364 7278 21416 7284
rect 21272 6384 21324 6390
rect 21272 6326 21324 6332
rect 21376 5778 21404 7278
rect 21652 6458 21680 7414
rect 21836 7342 21864 7822
rect 22388 7818 22416 9522
rect 22744 9512 22796 9518
rect 22744 9454 22796 9460
rect 22376 7812 22428 7818
rect 22376 7754 22428 7760
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 21824 7336 21876 7342
rect 21824 7278 21876 7284
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 22112 7002 22140 7278
rect 22100 6996 22152 7002
rect 22100 6938 22152 6944
rect 22008 6860 22060 6866
rect 22008 6802 22060 6808
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 21364 5772 21416 5778
rect 21364 5714 21416 5720
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 18420 5568 18472 5574
rect 18420 5510 18472 5516
rect 17972 5302 18000 5510
rect 18432 5370 18460 5510
rect 18420 5364 18472 5370
rect 18420 5306 18472 5312
rect 17960 5296 18012 5302
rect 17960 5238 18012 5244
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17328 4146 17356 5170
rect 17868 4548 17920 4554
rect 17868 4490 17920 4496
rect 17880 4282 17908 4490
rect 18432 4282 18460 5306
rect 18524 4826 18552 5630
rect 20904 5636 20956 5642
rect 20904 5578 20956 5584
rect 19656 5468 20032 5477
rect 19712 5466 19736 5468
rect 19792 5466 19816 5468
rect 19872 5466 19896 5468
rect 19952 5466 19976 5468
rect 19712 5414 19722 5466
rect 19966 5414 19976 5466
rect 19712 5412 19736 5414
rect 19792 5412 19816 5414
rect 19872 5412 19896 5414
rect 19952 5412 19976 5414
rect 19656 5403 20032 5412
rect 20916 5302 20944 5578
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 21192 5370 21220 5510
rect 21180 5364 21232 5370
rect 21180 5306 21232 5312
rect 20904 5296 20956 5302
rect 20904 5238 20956 5244
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 18916 4924 19292 4933
rect 18972 4922 18996 4924
rect 19052 4922 19076 4924
rect 19132 4922 19156 4924
rect 19212 4922 19236 4924
rect 18972 4870 18982 4922
rect 19226 4870 19236 4922
rect 18972 4868 18996 4870
rect 19052 4868 19076 4870
rect 19132 4868 19156 4870
rect 19212 4868 19236 4870
rect 18916 4859 19292 4868
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 18524 4690 18552 4762
rect 18512 4684 18564 4690
rect 18512 4626 18564 4632
rect 17868 4276 17920 4282
rect 17868 4218 17920 4224
rect 18420 4276 18472 4282
rect 18420 4218 18472 4224
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17328 3602 17356 4082
rect 18524 4078 18552 4626
rect 19656 4380 20032 4389
rect 19712 4378 19736 4380
rect 19792 4378 19816 4380
rect 19872 4378 19896 4380
rect 19952 4378 19976 4380
rect 19712 4326 19722 4378
rect 19966 4326 19976 4378
rect 19712 4324 19736 4326
rect 19792 4324 19816 4326
rect 19872 4324 19896 4326
rect 19952 4324 19976 4326
rect 19656 4315 20032 4324
rect 20444 4208 20496 4214
rect 20444 4150 20496 4156
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17420 3126 17448 3878
rect 18616 3738 18644 3946
rect 18916 3836 19292 3845
rect 18972 3834 18996 3836
rect 19052 3834 19076 3836
rect 19132 3834 19156 3836
rect 19212 3834 19236 3836
rect 18972 3782 18982 3834
rect 19226 3782 19236 3834
rect 18972 3780 18996 3782
rect 19052 3780 19076 3782
rect 19132 3780 19156 3782
rect 19212 3780 19236 3782
rect 18916 3771 19292 3780
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 17880 3194 17908 3402
rect 19536 3194 19564 3402
rect 20456 3398 20484 4150
rect 20732 4078 20760 5102
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 19656 3292 20032 3301
rect 19712 3290 19736 3292
rect 19792 3290 19816 3292
rect 19872 3290 19896 3292
rect 19952 3290 19976 3292
rect 19712 3238 19722 3290
rect 19966 3238 19976 3290
rect 19712 3236 19736 3238
rect 19792 3236 19816 3238
rect 19872 3236 19896 3238
rect 19952 3236 19976 3238
rect 19656 3227 20032 3236
rect 20456 3194 20484 3334
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 17408 3120 17460 3126
rect 17408 3062 17460 3068
rect 20732 2990 20760 4014
rect 21376 3602 21404 5714
rect 22020 5642 22048 6802
rect 21456 5636 21508 5642
rect 21456 5578 21508 5584
rect 22008 5636 22060 5642
rect 22008 5578 22060 5584
rect 21468 5370 21496 5578
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 21824 5296 21876 5302
rect 21824 5238 21876 5244
rect 21456 3936 21508 3942
rect 21456 3878 21508 3884
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21468 3466 21496 3878
rect 21836 3466 21864 5238
rect 21916 5160 21968 5166
rect 21916 5102 21968 5108
rect 21928 4826 21956 5102
rect 21916 4820 21968 4826
rect 21916 4762 21968 4768
rect 22020 4758 22048 5578
rect 22008 4752 22060 4758
rect 22008 4694 22060 4700
rect 22020 4078 22048 4694
rect 22296 4146 22324 7686
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 22572 6798 22600 7142
rect 22756 6866 22784 9454
rect 23388 8832 23440 8838
rect 23388 8774 23440 8780
rect 23400 8566 23428 8774
rect 23388 8560 23440 8566
rect 23388 8502 23440 8508
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 23400 7818 23428 8298
rect 23388 7812 23440 7818
rect 23388 7754 23440 7760
rect 24228 7342 24256 10542
rect 24412 8634 24440 10950
rect 24492 10532 24544 10538
rect 24492 10474 24544 10480
rect 24504 10130 24532 10474
rect 24492 10124 24544 10130
rect 24492 10066 24544 10072
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 24504 8430 24532 10066
rect 24492 8424 24544 8430
rect 24492 8366 24544 8372
rect 24400 7880 24452 7886
rect 24400 7822 24452 7828
rect 24216 7336 24268 7342
rect 24216 7278 24268 7284
rect 23664 7200 23716 7206
rect 23664 7142 23716 7148
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 23676 6798 23704 7142
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 23664 6792 23716 6798
rect 23664 6734 23716 6740
rect 23296 5024 23348 5030
rect 23296 4966 23348 4972
rect 23308 4622 23336 4966
rect 24228 4690 24256 7278
rect 24412 5370 24440 7822
rect 24596 7342 24624 11222
rect 24688 11082 24716 12158
rect 27656 11996 28032 12005
rect 27712 11994 27736 11996
rect 27792 11994 27816 11996
rect 27872 11994 27896 11996
rect 27952 11994 27976 11996
rect 27712 11942 27722 11994
rect 27966 11942 27976 11994
rect 27712 11940 27736 11942
rect 27792 11940 27816 11942
rect 27872 11940 27896 11942
rect 27952 11940 27976 11942
rect 27656 11931 28032 11940
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24780 11218 24808 11834
rect 26916 11452 27292 11461
rect 26972 11450 26996 11452
rect 27052 11450 27076 11452
rect 27132 11450 27156 11452
rect 27212 11450 27236 11452
rect 26972 11398 26982 11450
rect 27226 11398 27236 11450
rect 26972 11396 26996 11398
rect 27052 11396 27076 11398
rect 27132 11396 27156 11398
rect 27212 11396 27236 11398
rect 26916 11387 27292 11396
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 24676 11076 24728 11082
rect 24676 11018 24728 11024
rect 24688 10606 24716 11018
rect 24780 10742 24808 11154
rect 27656 10908 28032 10917
rect 27712 10906 27736 10908
rect 27792 10906 27816 10908
rect 27872 10906 27896 10908
rect 27952 10906 27976 10908
rect 27712 10854 27722 10906
rect 27966 10854 27976 10906
rect 27712 10852 27736 10854
rect 27792 10852 27816 10854
rect 27872 10852 27896 10854
rect 27952 10852 27976 10854
rect 27656 10843 28032 10852
rect 24768 10736 24820 10742
rect 24768 10678 24820 10684
rect 25044 10668 25096 10674
rect 25044 10610 25096 10616
rect 24676 10600 24728 10606
rect 24676 10542 24728 10548
rect 25056 9518 25084 10610
rect 26916 10364 27292 10373
rect 26972 10362 26996 10364
rect 27052 10362 27076 10364
rect 27132 10362 27156 10364
rect 27212 10362 27236 10364
rect 26972 10310 26982 10362
rect 27226 10310 27236 10362
rect 26972 10308 26996 10310
rect 27052 10308 27076 10310
rect 27132 10308 27156 10310
rect 27212 10308 27236 10310
rect 26916 10299 27292 10308
rect 27656 9820 28032 9829
rect 27712 9818 27736 9820
rect 27792 9818 27816 9820
rect 27872 9818 27896 9820
rect 27952 9818 27976 9820
rect 27712 9766 27722 9818
rect 27966 9766 27976 9818
rect 27712 9764 27736 9766
rect 27792 9764 27816 9766
rect 27872 9764 27896 9766
rect 27952 9764 27976 9766
rect 27656 9755 28032 9764
rect 25136 9648 25188 9654
rect 25136 9590 25188 9596
rect 25044 9512 25096 9518
rect 25044 9454 25096 9460
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 24688 7954 24716 8230
rect 24676 7948 24728 7954
rect 24676 7890 24728 7896
rect 24780 7750 24808 8434
rect 24768 7744 24820 7750
rect 24768 7686 24820 7692
rect 24780 7546 24808 7686
rect 25056 7546 25084 9454
rect 25148 8566 25176 9590
rect 26916 9276 27292 9285
rect 26972 9274 26996 9276
rect 27052 9274 27076 9276
rect 27132 9274 27156 9276
rect 27212 9274 27236 9276
rect 26972 9222 26982 9274
rect 27226 9222 27236 9274
rect 26972 9220 26996 9222
rect 27052 9220 27076 9222
rect 27132 9220 27156 9222
rect 27212 9220 27236 9222
rect 26916 9211 27292 9220
rect 27656 8732 28032 8741
rect 27712 8730 27736 8732
rect 27792 8730 27816 8732
rect 27872 8730 27896 8732
rect 27952 8730 27976 8732
rect 27712 8678 27722 8730
rect 27966 8678 27976 8730
rect 27712 8676 27736 8678
rect 27792 8676 27816 8678
rect 27872 8676 27896 8678
rect 27952 8676 27976 8678
rect 27656 8667 28032 8676
rect 25136 8560 25188 8566
rect 25136 8502 25188 8508
rect 25148 7818 25176 8502
rect 26916 8188 27292 8197
rect 26972 8186 26996 8188
rect 27052 8186 27076 8188
rect 27132 8186 27156 8188
rect 27212 8186 27236 8188
rect 26972 8134 26982 8186
rect 27226 8134 27236 8186
rect 26972 8132 26996 8134
rect 27052 8132 27076 8134
rect 27132 8132 27156 8134
rect 27212 8132 27236 8134
rect 26916 8123 27292 8132
rect 25136 7812 25188 7818
rect 25136 7754 25188 7760
rect 28356 7812 28408 7818
rect 28356 7754 28408 7760
rect 27656 7644 28032 7653
rect 27712 7642 27736 7644
rect 27792 7642 27816 7644
rect 27872 7642 27896 7644
rect 27952 7642 27976 7644
rect 27712 7590 27722 7642
rect 27966 7590 27976 7642
rect 27712 7588 27736 7590
rect 27792 7588 27816 7590
rect 27872 7588 27896 7590
rect 27952 7588 27976 7590
rect 27656 7579 28032 7588
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 25044 7540 25096 7546
rect 25044 7482 25096 7488
rect 28368 7449 28396 7754
rect 28354 7440 28410 7449
rect 28354 7375 28410 7384
rect 24584 7336 24636 7342
rect 24584 7278 24636 7284
rect 24768 7336 24820 7342
rect 24768 7278 24820 7284
rect 24676 7200 24728 7206
rect 24676 7142 24728 7148
rect 24400 5364 24452 5370
rect 24400 5306 24452 5312
rect 24688 4690 24716 7142
rect 24216 4684 24268 4690
rect 24216 4626 24268 4632
rect 24676 4684 24728 4690
rect 24676 4626 24728 4632
rect 23296 4616 23348 4622
rect 23296 4558 23348 4564
rect 22376 4480 22428 4486
rect 22376 4422 22428 4428
rect 22388 4282 22416 4422
rect 23308 4282 23336 4558
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 23296 4276 23348 4282
rect 23296 4218 23348 4224
rect 22836 4208 22888 4214
rect 22836 4150 22888 4156
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22008 4072 22060 4078
rect 22008 4014 22060 4020
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 21456 3460 21508 3466
rect 21456 3402 21508 3408
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 22664 3194 22692 3878
rect 22848 3738 22876 4150
rect 24780 4078 24808 7278
rect 26916 7100 27292 7109
rect 26972 7098 26996 7100
rect 27052 7098 27076 7100
rect 27132 7098 27156 7100
rect 27212 7098 27236 7100
rect 26972 7046 26982 7098
rect 27226 7046 27236 7098
rect 26972 7044 26996 7046
rect 27052 7044 27076 7046
rect 27132 7044 27156 7046
rect 27212 7044 27236 7046
rect 26916 7035 27292 7044
rect 27656 6556 28032 6565
rect 27712 6554 27736 6556
rect 27792 6554 27816 6556
rect 27872 6554 27896 6556
rect 27952 6554 27976 6556
rect 27712 6502 27722 6554
rect 27966 6502 27976 6554
rect 27712 6500 27736 6502
rect 27792 6500 27816 6502
rect 27872 6500 27896 6502
rect 27952 6500 27976 6502
rect 27656 6491 28032 6500
rect 26916 6012 27292 6021
rect 26972 6010 26996 6012
rect 27052 6010 27076 6012
rect 27132 6010 27156 6012
rect 27212 6010 27236 6012
rect 26972 5958 26982 6010
rect 27226 5958 27236 6010
rect 26972 5956 26996 5958
rect 27052 5956 27076 5958
rect 27132 5956 27156 5958
rect 27212 5956 27236 5958
rect 26916 5947 27292 5956
rect 27656 5468 28032 5477
rect 27712 5466 27736 5468
rect 27792 5466 27816 5468
rect 27872 5466 27896 5468
rect 27952 5466 27976 5468
rect 27712 5414 27722 5466
rect 27966 5414 27976 5466
rect 27712 5412 27736 5414
rect 27792 5412 27816 5414
rect 27872 5412 27896 5414
rect 27952 5412 27976 5414
rect 27656 5403 28032 5412
rect 25136 5160 25188 5166
rect 25136 5102 25188 5108
rect 25148 4826 25176 5102
rect 26916 4924 27292 4933
rect 26972 4922 26996 4924
rect 27052 4922 27076 4924
rect 27132 4922 27156 4924
rect 27212 4922 27236 4924
rect 26972 4870 26982 4922
rect 27226 4870 27236 4922
rect 26972 4868 26996 4870
rect 27052 4868 27076 4870
rect 27132 4868 27156 4870
rect 27212 4868 27236 4870
rect 26916 4859 27292 4868
rect 25136 4820 25188 4826
rect 25136 4762 25188 4768
rect 27656 4380 28032 4389
rect 27712 4378 27736 4380
rect 27792 4378 27816 4380
rect 27872 4378 27896 4380
rect 27952 4378 27976 4380
rect 27712 4326 27722 4378
rect 27966 4326 27976 4378
rect 27712 4324 27736 4326
rect 27792 4324 27816 4326
rect 27872 4324 27896 4326
rect 27952 4324 27976 4326
rect 27656 4315 28032 4324
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 26916 3836 27292 3845
rect 26972 3834 26996 3836
rect 27052 3834 27076 3836
rect 27132 3834 27156 3836
rect 27212 3834 27236 3836
rect 26972 3782 26982 3834
rect 27226 3782 27236 3834
rect 26972 3780 26996 3782
rect 27052 3780 27076 3782
rect 27132 3780 27156 3782
rect 27212 3780 27236 3782
rect 26916 3771 27292 3780
rect 22836 3732 22888 3738
rect 22836 3674 22888 3680
rect 27656 3292 28032 3301
rect 27712 3290 27736 3292
rect 27792 3290 27816 3292
rect 27872 3290 27896 3292
rect 27952 3290 27976 3292
rect 27712 3238 27722 3290
rect 27966 3238 27976 3290
rect 27712 3236 27736 3238
rect 27792 3236 27816 3238
rect 27872 3236 27896 3238
rect 27952 3236 27976 3238
rect 27656 3227 28032 3236
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 17132 2984 17184 2990
rect 17132 2926 17184 2932
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 14096 2916 14148 2922
rect 14096 2858 14148 2864
rect 2916 2748 3292 2757
rect 2972 2746 2996 2748
rect 3052 2746 3076 2748
rect 3132 2746 3156 2748
rect 3212 2746 3236 2748
rect 2972 2694 2982 2746
rect 3226 2694 3236 2746
rect 2972 2692 2996 2694
rect 3052 2692 3076 2694
rect 3132 2692 3156 2694
rect 3212 2692 3236 2694
rect 2916 2683 3292 2692
rect 10916 2748 11292 2757
rect 10972 2746 10996 2748
rect 11052 2746 11076 2748
rect 11132 2746 11156 2748
rect 11212 2746 11236 2748
rect 10972 2694 10982 2746
rect 11226 2694 11236 2746
rect 10972 2692 10996 2694
rect 11052 2692 11076 2694
rect 11132 2692 11156 2694
rect 11212 2692 11236 2694
rect 10916 2683 11292 2692
rect 18916 2748 19292 2757
rect 18972 2746 18996 2748
rect 19052 2746 19076 2748
rect 19132 2746 19156 2748
rect 19212 2746 19236 2748
rect 18972 2694 18982 2746
rect 19226 2694 19236 2746
rect 18972 2692 18996 2694
rect 19052 2692 19076 2694
rect 19132 2692 19156 2694
rect 19212 2692 19236 2694
rect 18916 2683 19292 2692
rect 26916 2748 27292 2757
rect 26972 2746 26996 2748
rect 27052 2746 27076 2748
rect 27132 2746 27156 2748
rect 27212 2746 27236 2748
rect 26972 2694 26982 2746
rect 27226 2694 27236 2746
rect 26972 2692 26996 2694
rect 27052 2692 27076 2694
rect 27132 2692 27156 2694
rect 27212 2692 27236 2694
rect 26916 2683 27292 2692
rect 3656 2204 4032 2213
rect 3712 2202 3736 2204
rect 3792 2202 3816 2204
rect 3872 2202 3896 2204
rect 3952 2202 3976 2204
rect 3712 2150 3722 2202
rect 3966 2150 3976 2202
rect 3712 2148 3736 2150
rect 3792 2148 3816 2150
rect 3872 2148 3896 2150
rect 3952 2148 3976 2150
rect 3656 2139 4032 2148
rect 11656 2204 12032 2213
rect 11712 2202 11736 2204
rect 11792 2202 11816 2204
rect 11872 2202 11896 2204
rect 11952 2202 11976 2204
rect 11712 2150 11722 2202
rect 11966 2150 11976 2202
rect 11712 2148 11736 2150
rect 11792 2148 11816 2150
rect 11872 2148 11896 2150
rect 11952 2148 11976 2150
rect 11656 2139 12032 2148
rect 19656 2204 20032 2213
rect 19712 2202 19736 2204
rect 19792 2202 19816 2204
rect 19872 2202 19896 2204
rect 19952 2202 19976 2204
rect 19712 2150 19722 2202
rect 19966 2150 19976 2202
rect 19712 2148 19736 2150
rect 19792 2148 19816 2150
rect 19872 2148 19896 2150
rect 19952 2148 19976 2150
rect 19656 2139 20032 2148
rect 27656 2204 28032 2213
rect 27712 2202 27736 2204
rect 27792 2202 27816 2204
rect 27872 2202 27896 2204
rect 27952 2202 27976 2204
rect 27712 2150 27722 2202
rect 27966 2150 27976 2202
rect 27712 2148 27736 2150
rect 27792 2148 27816 2150
rect 27872 2148 27896 2150
rect 27952 2148 27976 2150
rect 27656 2139 28032 2148
<< via2 >>
rect 2916 27770 2972 27772
rect 2996 27770 3052 27772
rect 3076 27770 3132 27772
rect 3156 27770 3212 27772
rect 3236 27770 3292 27772
rect 2916 27718 2918 27770
rect 2918 27718 2970 27770
rect 2970 27718 2972 27770
rect 2996 27718 3034 27770
rect 3034 27718 3046 27770
rect 3046 27718 3052 27770
rect 3076 27718 3098 27770
rect 3098 27718 3110 27770
rect 3110 27718 3132 27770
rect 3156 27718 3162 27770
rect 3162 27718 3174 27770
rect 3174 27718 3212 27770
rect 3236 27718 3238 27770
rect 3238 27718 3290 27770
rect 3290 27718 3292 27770
rect 2916 27716 2972 27718
rect 2996 27716 3052 27718
rect 3076 27716 3132 27718
rect 3156 27716 3212 27718
rect 3236 27716 3292 27718
rect 10916 27770 10972 27772
rect 10996 27770 11052 27772
rect 11076 27770 11132 27772
rect 11156 27770 11212 27772
rect 11236 27770 11292 27772
rect 10916 27718 10918 27770
rect 10918 27718 10970 27770
rect 10970 27718 10972 27770
rect 10996 27718 11034 27770
rect 11034 27718 11046 27770
rect 11046 27718 11052 27770
rect 11076 27718 11098 27770
rect 11098 27718 11110 27770
rect 11110 27718 11132 27770
rect 11156 27718 11162 27770
rect 11162 27718 11174 27770
rect 11174 27718 11212 27770
rect 11236 27718 11238 27770
rect 11238 27718 11290 27770
rect 11290 27718 11292 27770
rect 10916 27716 10972 27718
rect 10996 27716 11052 27718
rect 11076 27716 11132 27718
rect 11156 27716 11212 27718
rect 11236 27716 11292 27718
rect 18916 27770 18972 27772
rect 18996 27770 19052 27772
rect 19076 27770 19132 27772
rect 19156 27770 19212 27772
rect 19236 27770 19292 27772
rect 18916 27718 18918 27770
rect 18918 27718 18970 27770
rect 18970 27718 18972 27770
rect 18996 27718 19034 27770
rect 19034 27718 19046 27770
rect 19046 27718 19052 27770
rect 19076 27718 19098 27770
rect 19098 27718 19110 27770
rect 19110 27718 19132 27770
rect 19156 27718 19162 27770
rect 19162 27718 19174 27770
rect 19174 27718 19212 27770
rect 19236 27718 19238 27770
rect 19238 27718 19290 27770
rect 19290 27718 19292 27770
rect 18916 27716 18972 27718
rect 18996 27716 19052 27718
rect 19076 27716 19132 27718
rect 19156 27716 19212 27718
rect 19236 27716 19292 27718
rect 26916 27770 26972 27772
rect 26996 27770 27052 27772
rect 27076 27770 27132 27772
rect 27156 27770 27212 27772
rect 27236 27770 27292 27772
rect 26916 27718 26918 27770
rect 26918 27718 26970 27770
rect 26970 27718 26972 27770
rect 26996 27718 27034 27770
rect 27034 27718 27046 27770
rect 27046 27718 27052 27770
rect 27076 27718 27098 27770
rect 27098 27718 27110 27770
rect 27110 27718 27132 27770
rect 27156 27718 27162 27770
rect 27162 27718 27174 27770
rect 27174 27718 27212 27770
rect 27236 27718 27238 27770
rect 27238 27718 27290 27770
rect 27290 27718 27292 27770
rect 26916 27716 26972 27718
rect 26996 27716 27052 27718
rect 27076 27716 27132 27718
rect 27156 27716 27212 27718
rect 27236 27716 27292 27718
rect 3656 27226 3712 27228
rect 3736 27226 3792 27228
rect 3816 27226 3872 27228
rect 3896 27226 3952 27228
rect 3976 27226 4032 27228
rect 3656 27174 3658 27226
rect 3658 27174 3710 27226
rect 3710 27174 3712 27226
rect 3736 27174 3774 27226
rect 3774 27174 3786 27226
rect 3786 27174 3792 27226
rect 3816 27174 3838 27226
rect 3838 27174 3850 27226
rect 3850 27174 3872 27226
rect 3896 27174 3902 27226
rect 3902 27174 3914 27226
rect 3914 27174 3952 27226
rect 3976 27174 3978 27226
rect 3978 27174 4030 27226
rect 4030 27174 4032 27226
rect 3656 27172 3712 27174
rect 3736 27172 3792 27174
rect 3816 27172 3872 27174
rect 3896 27172 3952 27174
rect 3976 27172 4032 27174
rect 11656 27226 11712 27228
rect 11736 27226 11792 27228
rect 11816 27226 11872 27228
rect 11896 27226 11952 27228
rect 11976 27226 12032 27228
rect 11656 27174 11658 27226
rect 11658 27174 11710 27226
rect 11710 27174 11712 27226
rect 11736 27174 11774 27226
rect 11774 27174 11786 27226
rect 11786 27174 11792 27226
rect 11816 27174 11838 27226
rect 11838 27174 11850 27226
rect 11850 27174 11872 27226
rect 11896 27174 11902 27226
rect 11902 27174 11914 27226
rect 11914 27174 11952 27226
rect 11976 27174 11978 27226
rect 11978 27174 12030 27226
rect 12030 27174 12032 27226
rect 11656 27172 11712 27174
rect 11736 27172 11792 27174
rect 11816 27172 11872 27174
rect 11896 27172 11952 27174
rect 11976 27172 12032 27174
rect 19656 27226 19712 27228
rect 19736 27226 19792 27228
rect 19816 27226 19872 27228
rect 19896 27226 19952 27228
rect 19976 27226 20032 27228
rect 19656 27174 19658 27226
rect 19658 27174 19710 27226
rect 19710 27174 19712 27226
rect 19736 27174 19774 27226
rect 19774 27174 19786 27226
rect 19786 27174 19792 27226
rect 19816 27174 19838 27226
rect 19838 27174 19850 27226
rect 19850 27174 19872 27226
rect 19896 27174 19902 27226
rect 19902 27174 19914 27226
rect 19914 27174 19952 27226
rect 19976 27174 19978 27226
rect 19978 27174 20030 27226
rect 20030 27174 20032 27226
rect 19656 27172 19712 27174
rect 19736 27172 19792 27174
rect 19816 27172 19872 27174
rect 19896 27172 19952 27174
rect 19976 27172 20032 27174
rect 27656 27226 27712 27228
rect 27736 27226 27792 27228
rect 27816 27226 27872 27228
rect 27896 27226 27952 27228
rect 27976 27226 28032 27228
rect 27656 27174 27658 27226
rect 27658 27174 27710 27226
rect 27710 27174 27712 27226
rect 27736 27174 27774 27226
rect 27774 27174 27786 27226
rect 27786 27174 27792 27226
rect 27816 27174 27838 27226
rect 27838 27174 27850 27226
rect 27850 27174 27872 27226
rect 27896 27174 27902 27226
rect 27902 27174 27914 27226
rect 27914 27174 27952 27226
rect 27976 27174 27978 27226
rect 27978 27174 28030 27226
rect 28030 27174 28032 27226
rect 27656 27172 27712 27174
rect 27736 27172 27792 27174
rect 27816 27172 27872 27174
rect 27896 27172 27952 27174
rect 27976 27172 28032 27174
rect 2916 26682 2972 26684
rect 2996 26682 3052 26684
rect 3076 26682 3132 26684
rect 3156 26682 3212 26684
rect 3236 26682 3292 26684
rect 2916 26630 2918 26682
rect 2918 26630 2970 26682
rect 2970 26630 2972 26682
rect 2996 26630 3034 26682
rect 3034 26630 3046 26682
rect 3046 26630 3052 26682
rect 3076 26630 3098 26682
rect 3098 26630 3110 26682
rect 3110 26630 3132 26682
rect 3156 26630 3162 26682
rect 3162 26630 3174 26682
rect 3174 26630 3212 26682
rect 3236 26630 3238 26682
rect 3238 26630 3290 26682
rect 3290 26630 3292 26682
rect 2916 26628 2972 26630
rect 2996 26628 3052 26630
rect 3076 26628 3132 26630
rect 3156 26628 3212 26630
rect 3236 26628 3292 26630
rect 10916 26682 10972 26684
rect 10996 26682 11052 26684
rect 11076 26682 11132 26684
rect 11156 26682 11212 26684
rect 11236 26682 11292 26684
rect 10916 26630 10918 26682
rect 10918 26630 10970 26682
rect 10970 26630 10972 26682
rect 10996 26630 11034 26682
rect 11034 26630 11046 26682
rect 11046 26630 11052 26682
rect 11076 26630 11098 26682
rect 11098 26630 11110 26682
rect 11110 26630 11132 26682
rect 11156 26630 11162 26682
rect 11162 26630 11174 26682
rect 11174 26630 11212 26682
rect 11236 26630 11238 26682
rect 11238 26630 11290 26682
rect 11290 26630 11292 26682
rect 10916 26628 10972 26630
rect 10996 26628 11052 26630
rect 11076 26628 11132 26630
rect 11156 26628 11212 26630
rect 11236 26628 11292 26630
rect 18916 26682 18972 26684
rect 18996 26682 19052 26684
rect 19076 26682 19132 26684
rect 19156 26682 19212 26684
rect 19236 26682 19292 26684
rect 18916 26630 18918 26682
rect 18918 26630 18970 26682
rect 18970 26630 18972 26682
rect 18996 26630 19034 26682
rect 19034 26630 19046 26682
rect 19046 26630 19052 26682
rect 19076 26630 19098 26682
rect 19098 26630 19110 26682
rect 19110 26630 19132 26682
rect 19156 26630 19162 26682
rect 19162 26630 19174 26682
rect 19174 26630 19212 26682
rect 19236 26630 19238 26682
rect 19238 26630 19290 26682
rect 19290 26630 19292 26682
rect 18916 26628 18972 26630
rect 18996 26628 19052 26630
rect 19076 26628 19132 26630
rect 19156 26628 19212 26630
rect 19236 26628 19292 26630
rect 26916 26682 26972 26684
rect 26996 26682 27052 26684
rect 27076 26682 27132 26684
rect 27156 26682 27212 26684
rect 27236 26682 27292 26684
rect 26916 26630 26918 26682
rect 26918 26630 26970 26682
rect 26970 26630 26972 26682
rect 26996 26630 27034 26682
rect 27034 26630 27046 26682
rect 27046 26630 27052 26682
rect 27076 26630 27098 26682
rect 27098 26630 27110 26682
rect 27110 26630 27132 26682
rect 27156 26630 27162 26682
rect 27162 26630 27174 26682
rect 27174 26630 27212 26682
rect 27236 26630 27238 26682
rect 27238 26630 27290 26682
rect 27290 26630 27292 26682
rect 26916 26628 26972 26630
rect 26996 26628 27052 26630
rect 27076 26628 27132 26630
rect 27156 26628 27212 26630
rect 27236 26628 27292 26630
rect 3656 26138 3712 26140
rect 3736 26138 3792 26140
rect 3816 26138 3872 26140
rect 3896 26138 3952 26140
rect 3976 26138 4032 26140
rect 3656 26086 3658 26138
rect 3658 26086 3710 26138
rect 3710 26086 3712 26138
rect 3736 26086 3774 26138
rect 3774 26086 3786 26138
rect 3786 26086 3792 26138
rect 3816 26086 3838 26138
rect 3838 26086 3850 26138
rect 3850 26086 3872 26138
rect 3896 26086 3902 26138
rect 3902 26086 3914 26138
rect 3914 26086 3952 26138
rect 3976 26086 3978 26138
rect 3978 26086 4030 26138
rect 4030 26086 4032 26138
rect 3656 26084 3712 26086
rect 3736 26084 3792 26086
rect 3816 26084 3872 26086
rect 3896 26084 3952 26086
rect 3976 26084 4032 26086
rect 11656 26138 11712 26140
rect 11736 26138 11792 26140
rect 11816 26138 11872 26140
rect 11896 26138 11952 26140
rect 11976 26138 12032 26140
rect 11656 26086 11658 26138
rect 11658 26086 11710 26138
rect 11710 26086 11712 26138
rect 11736 26086 11774 26138
rect 11774 26086 11786 26138
rect 11786 26086 11792 26138
rect 11816 26086 11838 26138
rect 11838 26086 11850 26138
rect 11850 26086 11872 26138
rect 11896 26086 11902 26138
rect 11902 26086 11914 26138
rect 11914 26086 11952 26138
rect 11976 26086 11978 26138
rect 11978 26086 12030 26138
rect 12030 26086 12032 26138
rect 11656 26084 11712 26086
rect 11736 26084 11792 26086
rect 11816 26084 11872 26086
rect 11896 26084 11952 26086
rect 11976 26084 12032 26086
rect 19656 26138 19712 26140
rect 19736 26138 19792 26140
rect 19816 26138 19872 26140
rect 19896 26138 19952 26140
rect 19976 26138 20032 26140
rect 19656 26086 19658 26138
rect 19658 26086 19710 26138
rect 19710 26086 19712 26138
rect 19736 26086 19774 26138
rect 19774 26086 19786 26138
rect 19786 26086 19792 26138
rect 19816 26086 19838 26138
rect 19838 26086 19850 26138
rect 19850 26086 19872 26138
rect 19896 26086 19902 26138
rect 19902 26086 19914 26138
rect 19914 26086 19952 26138
rect 19976 26086 19978 26138
rect 19978 26086 20030 26138
rect 20030 26086 20032 26138
rect 19656 26084 19712 26086
rect 19736 26084 19792 26086
rect 19816 26084 19872 26086
rect 19896 26084 19952 26086
rect 19976 26084 20032 26086
rect 27656 26138 27712 26140
rect 27736 26138 27792 26140
rect 27816 26138 27872 26140
rect 27896 26138 27952 26140
rect 27976 26138 28032 26140
rect 27656 26086 27658 26138
rect 27658 26086 27710 26138
rect 27710 26086 27712 26138
rect 27736 26086 27774 26138
rect 27774 26086 27786 26138
rect 27786 26086 27792 26138
rect 27816 26086 27838 26138
rect 27838 26086 27850 26138
rect 27850 26086 27872 26138
rect 27896 26086 27902 26138
rect 27902 26086 27914 26138
rect 27914 26086 27952 26138
rect 27976 26086 27978 26138
rect 27978 26086 28030 26138
rect 28030 26086 28032 26138
rect 27656 26084 27712 26086
rect 27736 26084 27792 26086
rect 27816 26084 27872 26086
rect 27896 26084 27952 26086
rect 27976 26084 28032 26086
rect 2916 25594 2972 25596
rect 2996 25594 3052 25596
rect 3076 25594 3132 25596
rect 3156 25594 3212 25596
rect 3236 25594 3292 25596
rect 2916 25542 2918 25594
rect 2918 25542 2970 25594
rect 2970 25542 2972 25594
rect 2996 25542 3034 25594
rect 3034 25542 3046 25594
rect 3046 25542 3052 25594
rect 3076 25542 3098 25594
rect 3098 25542 3110 25594
rect 3110 25542 3132 25594
rect 3156 25542 3162 25594
rect 3162 25542 3174 25594
rect 3174 25542 3212 25594
rect 3236 25542 3238 25594
rect 3238 25542 3290 25594
rect 3290 25542 3292 25594
rect 2916 25540 2972 25542
rect 2996 25540 3052 25542
rect 3076 25540 3132 25542
rect 3156 25540 3212 25542
rect 3236 25540 3292 25542
rect 10916 25594 10972 25596
rect 10996 25594 11052 25596
rect 11076 25594 11132 25596
rect 11156 25594 11212 25596
rect 11236 25594 11292 25596
rect 10916 25542 10918 25594
rect 10918 25542 10970 25594
rect 10970 25542 10972 25594
rect 10996 25542 11034 25594
rect 11034 25542 11046 25594
rect 11046 25542 11052 25594
rect 11076 25542 11098 25594
rect 11098 25542 11110 25594
rect 11110 25542 11132 25594
rect 11156 25542 11162 25594
rect 11162 25542 11174 25594
rect 11174 25542 11212 25594
rect 11236 25542 11238 25594
rect 11238 25542 11290 25594
rect 11290 25542 11292 25594
rect 10916 25540 10972 25542
rect 10996 25540 11052 25542
rect 11076 25540 11132 25542
rect 11156 25540 11212 25542
rect 11236 25540 11292 25542
rect 18916 25594 18972 25596
rect 18996 25594 19052 25596
rect 19076 25594 19132 25596
rect 19156 25594 19212 25596
rect 19236 25594 19292 25596
rect 18916 25542 18918 25594
rect 18918 25542 18970 25594
rect 18970 25542 18972 25594
rect 18996 25542 19034 25594
rect 19034 25542 19046 25594
rect 19046 25542 19052 25594
rect 19076 25542 19098 25594
rect 19098 25542 19110 25594
rect 19110 25542 19132 25594
rect 19156 25542 19162 25594
rect 19162 25542 19174 25594
rect 19174 25542 19212 25594
rect 19236 25542 19238 25594
rect 19238 25542 19290 25594
rect 19290 25542 19292 25594
rect 18916 25540 18972 25542
rect 18996 25540 19052 25542
rect 19076 25540 19132 25542
rect 19156 25540 19212 25542
rect 19236 25540 19292 25542
rect 26916 25594 26972 25596
rect 26996 25594 27052 25596
rect 27076 25594 27132 25596
rect 27156 25594 27212 25596
rect 27236 25594 27292 25596
rect 26916 25542 26918 25594
rect 26918 25542 26970 25594
rect 26970 25542 26972 25594
rect 26996 25542 27034 25594
rect 27034 25542 27046 25594
rect 27046 25542 27052 25594
rect 27076 25542 27098 25594
rect 27098 25542 27110 25594
rect 27110 25542 27132 25594
rect 27156 25542 27162 25594
rect 27162 25542 27174 25594
rect 27174 25542 27212 25594
rect 27236 25542 27238 25594
rect 27238 25542 27290 25594
rect 27290 25542 27292 25594
rect 26916 25540 26972 25542
rect 26996 25540 27052 25542
rect 27076 25540 27132 25542
rect 27156 25540 27212 25542
rect 27236 25540 27292 25542
rect 1214 25064 1270 25120
rect 1306 24520 1362 24576
rect 1306 23976 1362 24032
rect 1306 23432 1362 23488
rect 1398 22888 1454 22944
rect 1214 22344 1270 22400
rect 1214 21800 1270 21856
rect 1306 21256 1362 21312
rect 1306 20712 1362 20768
rect 1582 20712 1638 20768
rect 1306 20168 1362 20224
rect 1306 19624 1362 19680
rect 1398 19080 1454 19136
rect 1306 18536 1362 18592
rect 1306 17992 1362 18048
rect 1214 17448 1270 17504
rect 1306 16904 1362 16960
rect 1490 16360 1546 16416
rect 1582 16244 1638 16280
rect 1582 16224 1584 16244
rect 1584 16224 1636 16244
rect 1636 16224 1638 16244
rect 1306 15816 1362 15872
rect 3656 25050 3712 25052
rect 3736 25050 3792 25052
rect 3816 25050 3872 25052
rect 3896 25050 3952 25052
rect 3976 25050 4032 25052
rect 3656 24998 3658 25050
rect 3658 24998 3710 25050
rect 3710 24998 3712 25050
rect 3736 24998 3774 25050
rect 3774 24998 3786 25050
rect 3786 24998 3792 25050
rect 3816 24998 3838 25050
rect 3838 24998 3850 25050
rect 3850 24998 3872 25050
rect 3896 24998 3902 25050
rect 3902 24998 3914 25050
rect 3914 24998 3952 25050
rect 3976 24998 3978 25050
rect 3978 24998 4030 25050
rect 4030 24998 4032 25050
rect 3656 24996 3712 24998
rect 3736 24996 3792 24998
rect 3816 24996 3872 24998
rect 3896 24996 3952 24998
rect 3976 24996 4032 24998
rect 11656 25050 11712 25052
rect 11736 25050 11792 25052
rect 11816 25050 11872 25052
rect 11896 25050 11952 25052
rect 11976 25050 12032 25052
rect 11656 24998 11658 25050
rect 11658 24998 11710 25050
rect 11710 24998 11712 25050
rect 11736 24998 11774 25050
rect 11774 24998 11786 25050
rect 11786 24998 11792 25050
rect 11816 24998 11838 25050
rect 11838 24998 11850 25050
rect 11850 24998 11872 25050
rect 11896 24998 11902 25050
rect 11902 24998 11914 25050
rect 11914 24998 11952 25050
rect 11976 24998 11978 25050
rect 11978 24998 12030 25050
rect 12030 24998 12032 25050
rect 11656 24996 11712 24998
rect 11736 24996 11792 24998
rect 11816 24996 11872 24998
rect 11896 24996 11952 24998
rect 11976 24996 12032 24998
rect 19656 25050 19712 25052
rect 19736 25050 19792 25052
rect 19816 25050 19872 25052
rect 19896 25050 19952 25052
rect 19976 25050 20032 25052
rect 19656 24998 19658 25050
rect 19658 24998 19710 25050
rect 19710 24998 19712 25050
rect 19736 24998 19774 25050
rect 19774 24998 19786 25050
rect 19786 24998 19792 25050
rect 19816 24998 19838 25050
rect 19838 24998 19850 25050
rect 19850 24998 19872 25050
rect 19896 24998 19902 25050
rect 19902 24998 19914 25050
rect 19914 24998 19952 25050
rect 19976 24998 19978 25050
rect 19978 24998 20030 25050
rect 20030 24998 20032 25050
rect 19656 24996 19712 24998
rect 19736 24996 19792 24998
rect 19816 24996 19872 24998
rect 19896 24996 19952 24998
rect 19976 24996 20032 24998
rect 27656 25050 27712 25052
rect 27736 25050 27792 25052
rect 27816 25050 27872 25052
rect 27896 25050 27952 25052
rect 27976 25050 28032 25052
rect 27656 24998 27658 25050
rect 27658 24998 27710 25050
rect 27710 24998 27712 25050
rect 27736 24998 27774 25050
rect 27774 24998 27786 25050
rect 27786 24998 27792 25050
rect 27816 24998 27838 25050
rect 27838 24998 27850 25050
rect 27850 24998 27872 25050
rect 27896 24998 27902 25050
rect 27902 24998 27914 25050
rect 27914 24998 27952 25050
rect 27976 24998 27978 25050
rect 27978 24998 28030 25050
rect 28030 24998 28032 25050
rect 27656 24996 27712 24998
rect 27736 24996 27792 24998
rect 27816 24996 27872 24998
rect 27896 24996 27952 24998
rect 27976 24996 28032 24998
rect 2916 24506 2972 24508
rect 2996 24506 3052 24508
rect 3076 24506 3132 24508
rect 3156 24506 3212 24508
rect 3236 24506 3292 24508
rect 2916 24454 2918 24506
rect 2918 24454 2970 24506
rect 2970 24454 2972 24506
rect 2996 24454 3034 24506
rect 3034 24454 3046 24506
rect 3046 24454 3052 24506
rect 3076 24454 3098 24506
rect 3098 24454 3110 24506
rect 3110 24454 3132 24506
rect 3156 24454 3162 24506
rect 3162 24454 3174 24506
rect 3174 24454 3212 24506
rect 3236 24454 3238 24506
rect 3238 24454 3290 24506
rect 3290 24454 3292 24506
rect 2916 24452 2972 24454
rect 2996 24452 3052 24454
rect 3076 24452 3132 24454
rect 3156 24452 3212 24454
rect 3236 24452 3292 24454
rect 10916 24506 10972 24508
rect 10996 24506 11052 24508
rect 11076 24506 11132 24508
rect 11156 24506 11212 24508
rect 11236 24506 11292 24508
rect 10916 24454 10918 24506
rect 10918 24454 10970 24506
rect 10970 24454 10972 24506
rect 10996 24454 11034 24506
rect 11034 24454 11046 24506
rect 11046 24454 11052 24506
rect 11076 24454 11098 24506
rect 11098 24454 11110 24506
rect 11110 24454 11132 24506
rect 11156 24454 11162 24506
rect 11162 24454 11174 24506
rect 11174 24454 11212 24506
rect 11236 24454 11238 24506
rect 11238 24454 11290 24506
rect 11290 24454 11292 24506
rect 10916 24452 10972 24454
rect 10996 24452 11052 24454
rect 11076 24452 11132 24454
rect 11156 24452 11212 24454
rect 11236 24452 11292 24454
rect 18916 24506 18972 24508
rect 18996 24506 19052 24508
rect 19076 24506 19132 24508
rect 19156 24506 19212 24508
rect 19236 24506 19292 24508
rect 18916 24454 18918 24506
rect 18918 24454 18970 24506
rect 18970 24454 18972 24506
rect 18996 24454 19034 24506
rect 19034 24454 19046 24506
rect 19046 24454 19052 24506
rect 19076 24454 19098 24506
rect 19098 24454 19110 24506
rect 19110 24454 19132 24506
rect 19156 24454 19162 24506
rect 19162 24454 19174 24506
rect 19174 24454 19212 24506
rect 19236 24454 19238 24506
rect 19238 24454 19290 24506
rect 19290 24454 19292 24506
rect 18916 24452 18972 24454
rect 18996 24452 19052 24454
rect 19076 24452 19132 24454
rect 19156 24452 19212 24454
rect 19236 24452 19292 24454
rect 26916 24506 26972 24508
rect 26996 24506 27052 24508
rect 27076 24506 27132 24508
rect 27156 24506 27212 24508
rect 27236 24506 27292 24508
rect 26916 24454 26918 24506
rect 26918 24454 26970 24506
rect 26970 24454 26972 24506
rect 26996 24454 27034 24506
rect 27034 24454 27046 24506
rect 27046 24454 27052 24506
rect 27076 24454 27098 24506
rect 27098 24454 27110 24506
rect 27110 24454 27132 24506
rect 27156 24454 27162 24506
rect 27162 24454 27174 24506
rect 27174 24454 27212 24506
rect 27236 24454 27238 24506
rect 27238 24454 27290 24506
rect 27290 24454 27292 24506
rect 26916 24452 26972 24454
rect 26996 24452 27052 24454
rect 27076 24452 27132 24454
rect 27156 24452 27212 24454
rect 27236 24452 27292 24454
rect 3656 23962 3712 23964
rect 3736 23962 3792 23964
rect 3816 23962 3872 23964
rect 3896 23962 3952 23964
rect 3976 23962 4032 23964
rect 3656 23910 3658 23962
rect 3658 23910 3710 23962
rect 3710 23910 3712 23962
rect 3736 23910 3774 23962
rect 3774 23910 3786 23962
rect 3786 23910 3792 23962
rect 3816 23910 3838 23962
rect 3838 23910 3850 23962
rect 3850 23910 3872 23962
rect 3896 23910 3902 23962
rect 3902 23910 3914 23962
rect 3914 23910 3952 23962
rect 3976 23910 3978 23962
rect 3978 23910 4030 23962
rect 4030 23910 4032 23962
rect 3656 23908 3712 23910
rect 3736 23908 3792 23910
rect 3816 23908 3872 23910
rect 3896 23908 3952 23910
rect 3976 23908 4032 23910
rect 2916 23418 2972 23420
rect 2996 23418 3052 23420
rect 3076 23418 3132 23420
rect 3156 23418 3212 23420
rect 3236 23418 3292 23420
rect 2916 23366 2918 23418
rect 2918 23366 2970 23418
rect 2970 23366 2972 23418
rect 2996 23366 3034 23418
rect 3034 23366 3046 23418
rect 3046 23366 3052 23418
rect 3076 23366 3098 23418
rect 3098 23366 3110 23418
rect 3110 23366 3132 23418
rect 3156 23366 3162 23418
rect 3162 23366 3174 23418
rect 3174 23366 3212 23418
rect 3236 23366 3238 23418
rect 3238 23366 3290 23418
rect 3290 23366 3292 23418
rect 2916 23364 2972 23366
rect 2996 23364 3052 23366
rect 3076 23364 3132 23366
rect 3156 23364 3212 23366
rect 3236 23364 3292 23366
rect 1398 15272 1454 15328
rect 1306 14728 1362 14784
rect 1306 14184 1362 14240
rect 1306 13640 1362 13696
rect 1214 13096 1270 13152
rect 1306 12552 1362 12608
rect 2916 22330 2972 22332
rect 2996 22330 3052 22332
rect 3076 22330 3132 22332
rect 3156 22330 3212 22332
rect 3236 22330 3292 22332
rect 2916 22278 2918 22330
rect 2918 22278 2970 22330
rect 2970 22278 2972 22330
rect 2996 22278 3034 22330
rect 3034 22278 3046 22330
rect 3046 22278 3052 22330
rect 3076 22278 3098 22330
rect 3098 22278 3110 22330
rect 3110 22278 3132 22330
rect 3156 22278 3162 22330
rect 3162 22278 3174 22330
rect 3174 22278 3212 22330
rect 3236 22278 3238 22330
rect 3238 22278 3290 22330
rect 3290 22278 3292 22330
rect 2916 22276 2972 22278
rect 2996 22276 3052 22278
rect 3076 22276 3132 22278
rect 3156 22276 3212 22278
rect 3236 22276 3292 22278
rect 2410 21292 2412 21312
rect 2412 21292 2464 21312
rect 2464 21292 2466 21312
rect 2410 21256 2466 21292
rect 1306 12008 1362 12064
rect 1950 12008 2006 12064
rect 1306 11464 1362 11520
rect 1398 10920 1454 10976
rect 1306 10376 1362 10432
rect 1306 9832 1362 9888
rect 2916 21242 2972 21244
rect 2996 21242 3052 21244
rect 3076 21242 3132 21244
rect 3156 21242 3212 21244
rect 3236 21242 3292 21244
rect 2916 21190 2918 21242
rect 2918 21190 2970 21242
rect 2970 21190 2972 21242
rect 2996 21190 3034 21242
rect 3034 21190 3046 21242
rect 3046 21190 3052 21242
rect 3076 21190 3098 21242
rect 3098 21190 3110 21242
rect 3110 21190 3132 21242
rect 3156 21190 3162 21242
rect 3162 21190 3174 21242
rect 3174 21190 3212 21242
rect 3236 21190 3238 21242
rect 3238 21190 3290 21242
rect 3290 21190 3292 21242
rect 2916 21188 2972 21190
rect 2996 21188 3052 21190
rect 3076 21188 3132 21190
rect 3156 21188 3212 21190
rect 3236 21188 3292 21190
rect 2594 19216 2650 19272
rect 3790 23060 3792 23080
rect 3792 23060 3844 23080
rect 3844 23060 3846 23080
rect 3790 23024 3846 23060
rect 2962 20304 3018 20360
rect 2916 20154 2972 20156
rect 2996 20154 3052 20156
rect 3076 20154 3132 20156
rect 3156 20154 3212 20156
rect 3236 20154 3292 20156
rect 2916 20102 2918 20154
rect 2918 20102 2970 20154
rect 2970 20102 2972 20154
rect 2996 20102 3034 20154
rect 3034 20102 3046 20154
rect 3046 20102 3052 20154
rect 3076 20102 3098 20154
rect 3098 20102 3110 20154
rect 3110 20102 3132 20154
rect 3156 20102 3162 20154
rect 3162 20102 3174 20154
rect 3174 20102 3212 20154
rect 3236 20102 3238 20154
rect 3238 20102 3290 20154
rect 3290 20102 3292 20154
rect 2916 20100 2972 20102
rect 2996 20100 3052 20102
rect 3076 20100 3132 20102
rect 3156 20100 3212 20102
rect 3236 20100 3292 20102
rect 2962 19896 3018 19952
rect 2870 19372 2926 19408
rect 2870 19352 2872 19372
rect 2872 19352 2924 19372
rect 2924 19352 2926 19372
rect 3656 22874 3712 22876
rect 3736 22874 3792 22876
rect 3816 22874 3872 22876
rect 3896 22874 3952 22876
rect 3976 22874 4032 22876
rect 3656 22822 3658 22874
rect 3658 22822 3710 22874
rect 3710 22822 3712 22874
rect 3736 22822 3774 22874
rect 3774 22822 3786 22874
rect 3786 22822 3792 22874
rect 3816 22822 3838 22874
rect 3838 22822 3850 22874
rect 3850 22822 3872 22874
rect 3896 22822 3902 22874
rect 3902 22822 3914 22874
rect 3914 22822 3952 22874
rect 3976 22822 3978 22874
rect 3978 22822 4030 22874
rect 4030 22822 4032 22874
rect 3656 22820 3712 22822
rect 3736 22820 3792 22822
rect 3816 22820 3872 22822
rect 3896 22820 3952 22822
rect 3976 22820 4032 22822
rect 4066 22480 4122 22536
rect 3974 21936 4030 21992
rect 3656 21786 3712 21788
rect 3736 21786 3792 21788
rect 3816 21786 3872 21788
rect 3896 21786 3952 21788
rect 3976 21786 4032 21788
rect 3656 21734 3658 21786
rect 3658 21734 3710 21786
rect 3710 21734 3712 21786
rect 3736 21734 3774 21786
rect 3774 21734 3786 21786
rect 3786 21734 3792 21786
rect 3816 21734 3838 21786
rect 3838 21734 3850 21786
rect 3850 21734 3872 21786
rect 3896 21734 3902 21786
rect 3902 21734 3914 21786
rect 3914 21734 3952 21786
rect 3976 21734 3978 21786
rect 3978 21734 4030 21786
rect 4030 21734 4032 21786
rect 3656 21732 3712 21734
rect 3736 21732 3792 21734
rect 3816 21732 3872 21734
rect 3896 21732 3952 21734
rect 3976 21732 4032 21734
rect 3656 20698 3712 20700
rect 3736 20698 3792 20700
rect 3816 20698 3872 20700
rect 3896 20698 3952 20700
rect 3976 20698 4032 20700
rect 3656 20646 3658 20698
rect 3658 20646 3710 20698
rect 3710 20646 3712 20698
rect 3736 20646 3774 20698
rect 3774 20646 3786 20698
rect 3786 20646 3792 20698
rect 3816 20646 3838 20698
rect 3838 20646 3850 20698
rect 3850 20646 3872 20698
rect 3896 20646 3902 20698
rect 3902 20646 3914 20698
rect 3914 20646 3952 20698
rect 3976 20646 3978 20698
rect 3978 20646 4030 20698
rect 4030 20646 4032 20698
rect 3656 20644 3712 20646
rect 3736 20644 3792 20646
rect 3816 20644 3872 20646
rect 3896 20644 3952 20646
rect 3976 20644 4032 20646
rect 2916 19066 2972 19068
rect 2996 19066 3052 19068
rect 3076 19066 3132 19068
rect 3156 19066 3212 19068
rect 3236 19066 3292 19068
rect 2916 19014 2918 19066
rect 2918 19014 2970 19066
rect 2970 19014 2972 19066
rect 2996 19014 3034 19066
rect 3034 19014 3046 19066
rect 3046 19014 3052 19066
rect 3076 19014 3098 19066
rect 3098 19014 3110 19066
rect 3110 19014 3132 19066
rect 3156 19014 3162 19066
rect 3162 19014 3174 19066
rect 3174 19014 3212 19066
rect 3236 19014 3238 19066
rect 3238 19014 3290 19066
rect 3290 19014 3292 19066
rect 2916 19012 2972 19014
rect 2996 19012 3052 19014
rect 3076 19012 3132 19014
rect 3156 19012 3212 19014
rect 3236 19012 3292 19014
rect 3054 18808 3110 18864
rect 3656 19610 3712 19612
rect 3736 19610 3792 19612
rect 3816 19610 3872 19612
rect 3896 19610 3952 19612
rect 3976 19610 4032 19612
rect 3656 19558 3658 19610
rect 3658 19558 3710 19610
rect 3710 19558 3712 19610
rect 3736 19558 3774 19610
rect 3774 19558 3786 19610
rect 3786 19558 3792 19610
rect 3816 19558 3838 19610
rect 3838 19558 3850 19610
rect 3850 19558 3872 19610
rect 3896 19558 3902 19610
rect 3902 19558 3914 19610
rect 3914 19558 3952 19610
rect 3976 19558 3978 19610
rect 3978 19558 4030 19610
rect 4030 19558 4032 19610
rect 3656 19556 3712 19558
rect 3736 19556 3792 19558
rect 3816 19556 3872 19558
rect 3896 19556 3952 19558
rect 3976 19556 4032 19558
rect 3882 19352 3938 19408
rect 3698 18808 3754 18864
rect 3330 18672 3386 18728
rect 3882 18672 3938 18728
rect 3656 18522 3712 18524
rect 3736 18522 3792 18524
rect 3816 18522 3872 18524
rect 3896 18522 3952 18524
rect 3976 18522 4032 18524
rect 3656 18470 3658 18522
rect 3658 18470 3710 18522
rect 3710 18470 3712 18522
rect 3736 18470 3774 18522
rect 3774 18470 3786 18522
rect 3786 18470 3792 18522
rect 3816 18470 3838 18522
rect 3838 18470 3850 18522
rect 3850 18470 3872 18522
rect 3896 18470 3902 18522
rect 3902 18470 3914 18522
rect 3914 18470 3952 18522
rect 3976 18470 3978 18522
rect 3978 18470 4030 18522
rect 4030 18470 4032 18522
rect 3656 18468 3712 18470
rect 3736 18468 3792 18470
rect 3816 18468 3872 18470
rect 3896 18468 3952 18470
rect 3976 18468 4032 18470
rect 2916 17978 2972 17980
rect 2996 17978 3052 17980
rect 3076 17978 3132 17980
rect 3156 17978 3212 17980
rect 3236 17978 3292 17980
rect 2916 17926 2918 17978
rect 2918 17926 2970 17978
rect 2970 17926 2972 17978
rect 2996 17926 3034 17978
rect 3034 17926 3046 17978
rect 3046 17926 3052 17978
rect 3076 17926 3098 17978
rect 3098 17926 3110 17978
rect 3110 17926 3132 17978
rect 3156 17926 3162 17978
rect 3162 17926 3174 17978
rect 3174 17926 3212 17978
rect 3236 17926 3238 17978
rect 3238 17926 3290 17978
rect 3290 17926 3292 17978
rect 2916 17924 2972 17926
rect 2996 17924 3052 17926
rect 3076 17924 3132 17926
rect 3156 17924 3212 17926
rect 3236 17924 3292 17926
rect 3054 17040 3110 17096
rect 2916 16890 2972 16892
rect 2996 16890 3052 16892
rect 3076 16890 3132 16892
rect 3156 16890 3212 16892
rect 3236 16890 3292 16892
rect 2916 16838 2918 16890
rect 2918 16838 2970 16890
rect 2970 16838 2972 16890
rect 2996 16838 3034 16890
rect 3034 16838 3046 16890
rect 3046 16838 3052 16890
rect 3076 16838 3098 16890
rect 3098 16838 3110 16890
rect 3110 16838 3132 16890
rect 3156 16838 3162 16890
rect 3162 16838 3174 16890
rect 3174 16838 3212 16890
rect 3236 16838 3238 16890
rect 3238 16838 3290 16890
rect 3290 16838 3292 16890
rect 2916 16836 2972 16838
rect 2996 16836 3052 16838
rect 3076 16836 3132 16838
rect 3156 16836 3212 16838
rect 3236 16836 3292 16838
rect 2916 15802 2972 15804
rect 2996 15802 3052 15804
rect 3076 15802 3132 15804
rect 3156 15802 3212 15804
rect 3236 15802 3292 15804
rect 2916 15750 2918 15802
rect 2918 15750 2970 15802
rect 2970 15750 2972 15802
rect 2996 15750 3034 15802
rect 3034 15750 3046 15802
rect 3046 15750 3052 15802
rect 3076 15750 3098 15802
rect 3098 15750 3110 15802
rect 3110 15750 3132 15802
rect 3156 15750 3162 15802
rect 3162 15750 3174 15802
rect 3174 15750 3212 15802
rect 3236 15750 3238 15802
rect 3238 15750 3290 15802
rect 3290 15750 3292 15802
rect 2916 15748 2972 15750
rect 2996 15748 3052 15750
rect 3076 15748 3132 15750
rect 3156 15748 3212 15750
rect 3236 15748 3292 15750
rect 4250 19352 4306 19408
rect 5814 19372 5870 19408
rect 11656 23962 11712 23964
rect 11736 23962 11792 23964
rect 11816 23962 11872 23964
rect 11896 23962 11952 23964
rect 11976 23962 12032 23964
rect 11656 23910 11658 23962
rect 11658 23910 11710 23962
rect 11710 23910 11712 23962
rect 11736 23910 11774 23962
rect 11774 23910 11786 23962
rect 11786 23910 11792 23962
rect 11816 23910 11838 23962
rect 11838 23910 11850 23962
rect 11850 23910 11872 23962
rect 11896 23910 11902 23962
rect 11902 23910 11914 23962
rect 11914 23910 11952 23962
rect 11976 23910 11978 23962
rect 11978 23910 12030 23962
rect 12030 23910 12032 23962
rect 11656 23908 11712 23910
rect 11736 23908 11792 23910
rect 11816 23908 11872 23910
rect 11896 23908 11952 23910
rect 11976 23908 12032 23910
rect 19656 23962 19712 23964
rect 19736 23962 19792 23964
rect 19816 23962 19872 23964
rect 19896 23962 19952 23964
rect 19976 23962 20032 23964
rect 19656 23910 19658 23962
rect 19658 23910 19710 23962
rect 19710 23910 19712 23962
rect 19736 23910 19774 23962
rect 19774 23910 19786 23962
rect 19786 23910 19792 23962
rect 19816 23910 19838 23962
rect 19838 23910 19850 23962
rect 19850 23910 19872 23962
rect 19896 23910 19902 23962
rect 19902 23910 19914 23962
rect 19914 23910 19952 23962
rect 19976 23910 19978 23962
rect 19978 23910 20030 23962
rect 20030 23910 20032 23962
rect 19656 23908 19712 23910
rect 19736 23908 19792 23910
rect 19816 23908 19872 23910
rect 19896 23908 19952 23910
rect 19976 23908 20032 23910
rect 27656 23962 27712 23964
rect 27736 23962 27792 23964
rect 27816 23962 27872 23964
rect 27896 23962 27952 23964
rect 27976 23962 28032 23964
rect 27656 23910 27658 23962
rect 27658 23910 27710 23962
rect 27710 23910 27712 23962
rect 27736 23910 27774 23962
rect 27774 23910 27786 23962
rect 27786 23910 27792 23962
rect 27816 23910 27838 23962
rect 27838 23910 27850 23962
rect 27850 23910 27872 23962
rect 27896 23910 27902 23962
rect 27902 23910 27914 23962
rect 27914 23910 27952 23962
rect 27976 23910 27978 23962
rect 27978 23910 28030 23962
rect 28030 23910 28032 23962
rect 27656 23908 27712 23910
rect 27736 23908 27792 23910
rect 27816 23908 27872 23910
rect 27896 23908 27952 23910
rect 27976 23908 28032 23910
rect 5814 19352 5816 19372
rect 5816 19352 5868 19372
rect 5868 19352 5870 19372
rect 5630 19236 5686 19272
rect 5630 19216 5632 19236
rect 5632 19216 5684 19236
rect 5684 19216 5686 19236
rect 3656 17434 3712 17436
rect 3736 17434 3792 17436
rect 3816 17434 3872 17436
rect 3896 17434 3952 17436
rect 3976 17434 4032 17436
rect 3656 17382 3658 17434
rect 3658 17382 3710 17434
rect 3710 17382 3712 17434
rect 3736 17382 3774 17434
rect 3774 17382 3786 17434
rect 3786 17382 3792 17434
rect 3816 17382 3838 17434
rect 3838 17382 3850 17434
rect 3850 17382 3872 17434
rect 3896 17382 3902 17434
rect 3902 17382 3914 17434
rect 3914 17382 3952 17434
rect 3976 17382 3978 17434
rect 3978 17382 4030 17434
rect 4030 17382 4032 17434
rect 3656 17380 3712 17382
rect 3736 17380 3792 17382
rect 3816 17380 3872 17382
rect 3896 17380 3952 17382
rect 3976 17380 4032 17382
rect 3656 16346 3712 16348
rect 3736 16346 3792 16348
rect 3816 16346 3872 16348
rect 3896 16346 3952 16348
rect 3976 16346 4032 16348
rect 3656 16294 3658 16346
rect 3658 16294 3710 16346
rect 3710 16294 3712 16346
rect 3736 16294 3774 16346
rect 3774 16294 3786 16346
rect 3786 16294 3792 16346
rect 3816 16294 3838 16346
rect 3838 16294 3850 16346
rect 3850 16294 3872 16346
rect 3896 16294 3902 16346
rect 3902 16294 3914 16346
rect 3914 16294 3952 16346
rect 3976 16294 3978 16346
rect 3978 16294 4030 16346
rect 4030 16294 4032 16346
rect 3656 16292 3712 16294
rect 3736 16292 3792 16294
rect 3816 16292 3872 16294
rect 3896 16292 3952 16294
rect 3976 16292 4032 16294
rect 2962 15020 3018 15056
rect 2962 15000 2964 15020
rect 2964 15000 3016 15020
rect 3016 15000 3018 15020
rect 2916 14714 2972 14716
rect 2996 14714 3052 14716
rect 3076 14714 3132 14716
rect 3156 14714 3212 14716
rect 3236 14714 3292 14716
rect 2916 14662 2918 14714
rect 2918 14662 2970 14714
rect 2970 14662 2972 14714
rect 2996 14662 3034 14714
rect 3034 14662 3046 14714
rect 3046 14662 3052 14714
rect 3076 14662 3098 14714
rect 3098 14662 3110 14714
rect 3110 14662 3132 14714
rect 3156 14662 3162 14714
rect 3162 14662 3174 14714
rect 3174 14662 3212 14714
rect 3236 14662 3238 14714
rect 3238 14662 3290 14714
rect 3290 14662 3292 14714
rect 2916 14660 2972 14662
rect 2996 14660 3052 14662
rect 3076 14660 3132 14662
rect 3156 14660 3212 14662
rect 3236 14660 3292 14662
rect 2962 13932 3018 13968
rect 2962 13912 2964 13932
rect 2964 13912 3016 13932
rect 3016 13912 3018 13932
rect 3656 15258 3712 15260
rect 3736 15258 3792 15260
rect 3816 15258 3872 15260
rect 3896 15258 3952 15260
rect 3976 15258 4032 15260
rect 3656 15206 3658 15258
rect 3658 15206 3710 15258
rect 3710 15206 3712 15258
rect 3736 15206 3774 15258
rect 3774 15206 3786 15258
rect 3786 15206 3792 15258
rect 3816 15206 3838 15258
rect 3838 15206 3850 15258
rect 3850 15206 3872 15258
rect 3896 15206 3902 15258
rect 3902 15206 3914 15258
rect 3914 15206 3952 15258
rect 3976 15206 3978 15258
rect 3978 15206 4030 15258
rect 4030 15206 4032 15258
rect 3656 15204 3712 15206
rect 3736 15204 3792 15206
rect 3816 15204 3872 15206
rect 3896 15204 3952 15206
rect 3976 15204 4032 15206
rect 3656 14170 3712 14172
rect 3736 14170 3792 14172
rect 3816 14170 3872 14172
rect 3896 14170 3952 14172
rect 3976 14170 4032 14172
rect 3656 14118 3658 14170
rect 3658 14118 3710 14170
rect 3710 14118 3712 14170
rect 3736 14118 3774 14170
rect 3774 14118 3786 14170
rect 3786 14118 3792 14170
rect 3816 14118 3838 14170
rect 3838 14118 3850 14170
rect 3850 14118 3872 14170
rect 3896 14118 3902 14170
rect 3902 14118 3914 14170
rect 3914 14118 3952 14170
rect 3976 14118 3978 14170
rect 3978 14118 4030 14170
rect 4030 14118 4032 14170
rect 3656 14116 3712 14118
rect 3736 14116 3792 14118
rect 3816 14116 3872 14118
rect 3896 14116 3952 14118
rect 3976 14116 4032 14118
rect 3514 13912 3570 13968
rect 2916 13626 2972 13628
rect 2996 13626 3052 13628
rect 3076 13626 3132 13628
rect 3156 13626 3212 13628
rect 3236 13626 3292 13628
rect 2916 13574 2918 13626
rect 2918 13574 2970 13626
rect 2970 13574 2972 13626
rect 2996 13574 3034 13626
rect 3034 13574 3046 13626
rect 3046 13574 3052 13626
rect 3076 13574 3098 13626
rect 3098 13574 3110 13626
rect 3110 13574 3132 13626
rect 3156 13574 3162 13626
rect 3162 13574 3174 13626
rect 3174 13574 3212 13626
rect 3236 13574 3238 13626
rect 3238 13574 3290 13626
rect 3290 13574 3292 13626
rect 2916 13572 2972 13574
rect 2996 13572 3052 13574
rect 3076 13572 3132 13574
rect 3156 13572 3212 13574
rect 3236 13572 3292 13574
rect 3882 13932 3938 13968
rect 3882 13912 3884 13932
rect 3884 13912 3936 13932
rect 3936 13912 3938 13932
rect 2916 12538 2972 12540
rect 2996 12538 3052 12540
rect 3076 12538 3132 12540
rect 3156 12538 3212 12540
rect 3236 12538 3292 12540
rect 2916 12486 2918 12538
rect 2918 12486 2970 12538
rect 2970 12486 2972 12538
rect 2996 12486 3034 12538
rect 3034 12486 3046 12538
rect 3046 12486 3052 12538
rect 3076 12486 3098 12538
rect 3098 12486 3110 12538
rect 3110 12486 3132 12538
rect 3156 12486 3162 12538
rect 3162 12486 3174 12538
rect 3174 12486 3212 12538
rect 3236 12486 3238 12538
rect 3238 12486 3290 12538
rect 3290 12486 3292 12538
rect 2916 12484 2972 12486
rect 2996 12484 3052 12486
rect 3076 12484 3132 12486
rect 3156 12484 3212 12486
rect 3236 12484 3292 12486
rect 3656 13082 3712 13084
rect 3736 13082 3792 13084
rect 3816 13082 3872 13084
rect 3896 13082 3952 13084
rect 3976 13082 4032 13084
rect 3656 13030 3658 13082
rect 3658 13030 3710 13082
rect 3710 13030 3712 13082
rect 3736 13030 3774 13082
rect 3774 13030 3786 13082
rect 3786 13030 3792 13082
rect 3816 13030 3838 13082
rect 3838 13030 3850 13082
rect 3850 13030 3872 13082
rect 3896 13030 3902 13082
rect 3902 13030 3914 13082
rect 3914 13030 3952 13082
rect 3976 13030 3978 13082
rect 3978 13030 4030 13082
rect 4030 13030 4032 13082
rect 3656 13028 3712 13030
rect 3736 13028 3792 13030
rect 3816 13028 3872 13030
rect 3896 13028 3952 13030
rect 3976 13028 4032 13030
rect 3656 11994 3712 11996
rect 3736 11994 3792 11996
rect 3816 11994 3872 11996
rect 3896 11994 3952 11996
rect 3976 11994 4032 11996
rect 3656 11942 3658 11994
rect 3658 11942 3710 11994
rect 3710 11942 3712 11994
rect 3736 11942 3774 11994
rect 3774 11942 3786 11994
rect 3786 11942 3792 11994
rect 3816 11942 3838 11994
rect 3838 11942 3850 11994
rect 3850 11942 3872 11994
rect 3896 11942 3902 11994
rect 3902 11942 3914 11994
rect 3914 11942 3952 11994
rect 3976 11942 3978 11994
rect 3978 11942 4030 11994
rect 4030 11942 4032 11994
rect 3656 11940 3712 11942
rect 3736 11940 3792 11942
rect 3816 11940 3872 11942
rect 3896 11940 3952 11942
rect 3976 11940 4032 11942
rect 2916 11450 2972 11452
rect 2996 11450 3052 11452
rect 3076 11450 3132 11452
rect 3156 11450 3212 11452
rect 3236 11450 3292 11452
rect 2916 11398 2918 11450
rect 2918 11398 2970 11450
rect 2970 11398 2972 11450
rect 2996 11398 3034 11450
rect 3034 11398 3046 11450
rect 3046 11398 3052 11450
rect 3076 11398 3098 11450
rect 3098 11398 3110 11450
rect 3110 11398 3132 11450
rect 3156 11398 3162 11450
rect 3162 11398 3174 11450
rect 3174 11398 3212 11450
rect 3236 11398 3238 11450
rect 3238 11398 3290 11450
rect 3290 11398 3292 11450
rect 2916 11396 2972 11398
rect 2996 11396 3052 11398
rect 3076 11396 3132 11398
rect 3156 11396 3212 11398
rect 3236 11396 3292 11398
rect 3790 11348 3846 11384
rect 3790 11328 3792 11348
rect 3792 11328 3844 11348
rect 3844 11328 3846 11348
rect 5906 16532 5908 16552
rect 5908 16532 5960 16552
rect 5960 16532 5962 16552
rect 5906 16496 5962 16532
rect 3656 10906 3712 10908
rect 3736 10906 3792 10908
rect 3816 10906 3872 10908
rect 3896 10906 3952 10908
rect 3976 10906 4032 10908
rect 3656 10854 3658 10906
rect 3658 10854 3710 10906
rect 3710 10854 3712 10906
rect 3736 10854 3774 10906
rect 3774 10854 3786 10906
rect 3786 10854 3792 10906
rect 3816 10854 3838 10906
rect 3838 10854 3850 10906
rect 3850 10854 3872 10906
rect 3896 10854 3902 10906
rect 3902 10854 3914 10906
rect 3914 10854 3952 10906
rect 3976 10854 3978 10906
rect 3978 10854 4030 10906
rect 4030 10854 4032 10906
rect 3656 10852 3712 10854
rect 3736 10852 3792 10854
rect 3816 10852 3872 10854
rect 3896 10852 3952 10854
rect 3976 10852 4032 10854
rect 1306 9288 1362 9344
rect 1306 8780 1308 8800
rect 1308 8780 1360 8800
rect 1360 8780 1362 8800
rect 1306 8744 1362 8780
rect 1306 8200 1362 8256
rect 1214 7656 1270 7712
rect 2916 10362 2972 10364
rect 2996 10362 3052 10364
rect 3076 10362 3132 10364
rect 3156 10362 3212 10364
rect 3236 10362 3292 10364
rect 2916 10310 2918 10362
rect 2918 10310 2970 10362
rect 2970 10310 2972 10362
rect 2996 10310 3034 10362
rect 3034 10310 3046 10362
rect 3046 10310 3052 10362
rect 3076 10310 3098 10362
rect 3098 10310 3110 10362
rect 3110 10310 3132 10362
rect 3156 10310 3162 10362
rect 3162 10310 3174 10362
rect 3174 10310 3212 10362
rect 3236 10310 3238 10362
rect 3238 10310 3290 10362
rect 3290 10310 3292 10362
rect 2916 10308 2972 10310
rect 2996 10308 3052 10310
rect 3076 10308 3132 10310
rect 3156 10308 3212 10310
rect 3236 10308 3292 10310
rect 3656 9818 3712 9820
rect 3736 9818 3792 9820
rect 3816 9818 3872 9820
rect 3896 9818 3952 9820
rect 3976 9818 4032 9820
rect 3656 9766 3658 9818
rect 3658 9766 3710 9818
rect 3710 9766 3712 9818
rect 3736 9766 3774 9818
rect 3774 9766 3786 9818
rect 3786 9766 3792 9818
rect 3816 9766 3838 9818
rect 3838 9766 3850 9818
rect 3850 9766 3872 9818
rect 3896 9766 3902 9818
rect 3902 9766 3914 9818
rect 3914 9766 3952 9818
rect 3976 9766 3978 9818
rect 3978 9766 4030 9818
rect 4030 9766 4032 9818
rect 3656 9764 3712 9766
rect 3736 9764 3792 9766
rect 3816 9764 3872 9766
rect 3896 9764 3952 9766
rect 3976 9764 4032 9766
rect 2916 9274 2972 9276
rect 2996 9274 3052 9276
rect 3076 9274 3132 9276
rect 3156 9274 3212 9276
rect 3236 9274 3292 9276
rect 2916 9222 2918 9274
rect 2918 9222 2970 9274
rect 2970 9222 2972 9274
rect 2996 9222 3034 9274
rect 3034 9222 3046 9274
rect 3046 9222 3052 9274
rect 3076 9222 3098 9274
rect 3098 9222 3110 9274
rect 3110 9222 3132 9274
rect 3156 9222 3162 9274
rect 3162 9222 3174 9274
rect 3174 9222 3212 9274
rect 3236 9222 3238 9274
rect 3238 9222 3290 9274
rect 3290 9222 3292 9274
rect 2916 9220 2972 9222
rect 2996 9220 3052 9222
rect 3076 9220 3132 9222
rect 3156 9220 3212 9222
rect 3236 9220 3292 9222
rect 1214 7112 1270 7168
rect 1306 6568 1362 6624
rect 1306 6024 1362 6080
rect 1306 5480 1362 5536
rect 2916 8186 2972 8188
rect 2996 8186 3052 8188
rect 3076 8186 3132 8188
rect 3156 8186 3212 8188
rect 3236 8186 3292 8188
rect 2916 8134 2918 8186
rect 2918 8134 2970 8186
rect 2970 8134 2972 8186
rect 2996 8134 3034 8186
rect 3034 8134 3046 8186
rect 3046 8134 3052 8186
rect 3076 8134 3098 8186
rect 3098 8134 3110 8186
rect 3110 8134 3132 8186
rect 3156 8134 3162 8186
rect 3162 8134 3174 8186
rect 3174 8134 3212 8186
rect 3236 8134 3238 8186
rect 3238 8134 3290 8186
rect 3290 8134 3292 8186
rect 2916 8132 2972 8134
rect 2996 8132 3052 8134
rect 3076 8132 3132 8134
rect 3156 8132 3212 8134
rect 3236 8132 3292 8134
rect 2916 7098 2972 7100
rect 2996 7098 3052 7100
rect 3076 7098 3132 7100
rect 3156 7098 3212 7100
rect 3236 7098 3292 7100
rect 2916 7046 2918 7098
rect 2918 7046 2970 7098
rect 2970 7046 2972 7098
rect 2996 7046 3034 7098
rect 3034 7046 3046 7098
rect 3046 7046 3052 7098
rect 3076 7046 3098 7098
rect 3098 7046 3110 7098
rect 3110 7046 3132 7098
rect 3156 7046 3162 7098
rect 3162 7046 3174 7098
rect 3174 7046 3212 7098
rect 3236 7046 3238 7098
rect 3238 7046 3290 7098
rect 3290 7046 3292 7098
rect 2916 7044 2972 7046
rect 2996 7044 3052 7046
rect 3076 7044 3132 7046
rect 3156 7044 3212 7046
rect 3236 7044 3292 7046
rect 2916 6010 2972 6012
rect 2996 6010 3052 6012
rect 3076 6010 3132 6012
rect 3156 6010 3212 6012
rect 3236 6010 3292 6012
rect 2916 5958 2918 6010
rect 2918 5958 2970 6010
rect 2970 5958 2972 6010
rect 2996 5958 3034 6010
rect 3034 5958 3046 6010
rect 3046 5958 3052 6010
rect 3076 5958 3098 6010
rect 3098 5958 3110 6010
rect 3110 5958 3132 6010
rect 3156 5958 3162 6010
rect 3162 5958 3174 6010
rect 3174 5958 3212 6010
rect 3236 5958 3238 6010
rect 3238 5958 3290 6010
rect 3290 5958 3292 6010
rect 2916 5956 2972 5958
rect 2996 5956 3052 5958
rect 3076 5956 3132 5958
rect 3156 5956 3212 5958
rect 3236 5956 3292 5958
rect 1306 4936 1362 4992
rect 2916 4922 2972 4924
rect 2996 4922 3052 4924
rect 3076 4922 3132 4924
rect 3156 4922 3212 4924
rect 3236 4922 3292 4924
rect 2916 4870 2918 4922
rect 2918 4870 2970 4922
rect 2970 4870 2972 4922
rect 2996 4870 3034 4922
rect 3034 4870 3046 4922
rect 3046 4870 3052 4922
rect 3076 4870 3098 4922
rect 3098 4870 3110 4922
rect 3110 4870 3132 4922
rect 3156 4870 3162 4922
rect 3162 4870 3174 4922
rect 3174 4870 3212 4922
rect 3236 4870 3238 4922
rect 3238 4870 3290 4922
rect 3290 4870 3292 4922
rect 2916 4868 2972 4870
rect 2996 4868 3052 4870
rect 3076 4868 3132 4870
rect 3156 4868 3212 4870
rect 3236 4868 3292 4870
rect 1030 4392 1086 4448
rect 3656 8730 3712 8732
rect 3736 8730 3792 8732
rect 3816 8730 3872 8732
rect 3896 8730 3952 8732
rect 3976 8730 4032 8732
rect 3656 8678 3658 8730
rect 3658 8678 3710 8730
rect 3710 8678 3712 8730
rect 3736 8678 3774 8730
rect 3774 8678 3786 8730
rect 3786 8678 3792 8730
rect 3816 8678 3838 8730
rect 3838 8678 3850 8730
rect 3850 8678 3872 8730
rect 3896 8678 3902 8730
rect 3902 8678 3914 8730
rect 3914 8678 3952 8730
rect 3976 8678 3978 8730
rect 3978 8678 4030 8730
rect 4030 8678 4032 8730
rect 3656 8676 3712 8678
rect 3736 8676 3792 8678
rect 3816 8676 3872 8678
rect 3896 8676 3952 8678
rect 3976 8676 4032 8678
rect 10916 23418 10972 23420
rect 10996 23418 11052 23420
rect 11076 23418 11132 23420
rect 11156 23418 11212 23420
rect 11236 23418 11292 23420
rect 10916 23366 10918 23418
rect 10918 23366 10970 23418
rect 10970 23366 10972 23418
rect 10996 23366 11034 23418
rect 11034 23366 11046 23418
rect 11046 23366 11052 23418
rect 11076 23366 11098 23418
rect 11098 23366 11110 23418
rect 11110 23366 11132 23418
rect 11156 23366 11162 23418
rect 11162 23366 11174 23418
rect 11174 23366 11212 23418
rect 11236 23366 11238 23418
rect 11238 23366 11290 23418
rect 11290 23366 11292 23418
rect 10916 23364 10972 23366
rect 10996 23364 11052 23366
rect 11076 23364 11132 23366
rect 11156 23364 11212 23366
rect 11236 23364 11292 23366
rect 18916 23418 18972 23420
rect 18996 23418 19052 23420
rect 19076 23418 19132 23420
rect 19156 23418 19212 23420
rect 19236 23418 19292 23420
rect 18916 23366 18918 23418
rect 18918 23366 18970 23418
rect 18970 23366 18972 23418
rect 18996 23366 19034 23418
rect 19034 23366 19046 23418
rect 19046 23366 19052 23418
rect 19076 23366 19098 23418
rect 19098 23366 19110 23418
rect 19110 23366 19132 23418
rect 19156 23366 19162 23418
rect 19162 23366 19174 23418
rect 19174 23366 19212 23418
rect 19236 23366 19238 23418
rect 19238 23366 19290 23418
rect 19290 23366 19292 23418
rect 18916 23364 18972 23366
rect 18996 23364 19052 23366
rect 19076 23364 19132 23366
rect 19156 23364 19212 23366
rect 19236 23364 19292 23366
rect 26916 23418 26972 23420
rect 26996 23418 27052 23420
rect 27076 23418 27132 23420
rect 27156 23418 27212 23420
rect 27236 23418 27292 23420
rect 26916 23366 26918 23418
rect 26918 23366 26970 23418
rect 26970 23366 26972 23418
rect 26996 23366 27034 23418
rect 27034 23366 27046 23418
rect 27046 23366 27052 23418
rect 27076 23366 27098 23418
rect 27098 23366 27110 23418
rect 27110 23366 27132 23418
rect 27156 23366 27162 23418
rect 27162 23366 27174 23418
rect 27174 23366 27212 23418
rect 27236 23366 27238 23418
rect 27238 23366 27290 23418
rect 27290 23366 27292 23418
rect 26916 23364 26972 23366
rect 26996 23364 27052 23366
rect 27076 23364 27132 23366
rect 27156 23364 27212 23366
rect 27236 23364 27292 23366
rect 11656 22874 11712 22876
rect 11736 22874 11792 22876
rect 11816 22874 11872 22876
rect 11896 22874 11952 22876
rect 11976 22874 12032 22876
rect 11656 22822 11658 22874
rect 11658 22822 11710 22874
rect 11710 22822 11712 22874
rect 11736 22822 11774 22874
rect 11774 22822 11786 22874
rect 11786 22822 11792 22874
rect 11816 22822 11838 22874
rect 11838 22822 11850 22874
rect 11850 22822 11872 22874
rect 11896 22822 11902 22874
rect 11902 22822 11914 22874
rect 11914 22822 11952 22874
rect 11976 22822 11978 22874
rect 11978 22822 12030 22874
rect 12030 22822 12032 22874
rect 11656 22820 11712 22822
rect 11736 22820 11792 22822
rect 11816 22820 11872 22822
rect 11896 22820 11952 22822
rect 11976 22820 12032 22822
rect 19656 22874 19712 22876
rect 19736 22874 19792 22876
rect 19816 22874 19872 22876
rect 19896 22874 19952 22876
rect 19976 22874 20032 22876
rect 19656 22822 19658 22874
rect 19658 22822 19710 22874
rect 19710 22822 19712 22874
rect 19736 22822 19774 22874
rect 19774 22822 19786 22874
rect 19786 22822 19792 22874
rect 19816 22822 19838 22874
rect 19838 22822 19850 22874
rect 19850 22822 19872 22874
rect 19896 22822 19902 22874
rect 19902 22822 19914 22874
rect 19914 22822 19952 22874
rect 19976 22822 19978 22874
rect 19978 22822 20030 22874
rect 20030 22822 20032 22874
rect 19656 22820 19712 22822
rect 19736 22820 19792 22822
rect 19816 22820 19872 22822
rect 19896 22820 19952 22822
rect 19976 22820 20032 22822
rect 27656 22874 27712 22876
rect 27736 22874 27792 22876
rect 27816 22874 27872 22876
rect 27896 22874 27952 22876
rect 27976 22874 28032 22876
rect 27656 22822 27658 22874
rect 27658 22822 27710 22874
rect 27710 22822 27712 22874
rect 27736 22822 27774 22874
rect 27774 22822 27786 22874
rect 27786 22822 27792 22874
rect 27816 22822 27838 22874
rect 27838 22822 27850 22874
rect 27850 22822 27872 22874
rect 27896 22822 27902 22874
rect 27902 22822 27914 22874
rect 27914 22822 27952 22874
rect 27976 22822 27978 22874
rect 27978 22822 28030 22874
rect 28030 22822 28032 22874
rect 27656 22820 27712 22822
rect 27736 22820 27792 22822
rect 27816 22820 27872 22822
rect 27896 22820 27952 22822
rect 27976 22820 28032 22822
rect 10916 22330 10972 22332
rect 10996 22330 11052 22332
rect 11076 22330 11132 22332
rect 11156 22330 11212 22332
rect 11236 22330 11292 22332
rect 10916 22278 10918 22330
rect 10918 22278 10970 22330
rect 10970 22278 10972 22330
rect 10996 22278 11034 22330
rect 11034 22278 11046 22330
rect 11046 22278 11052 22330
rect 11076 22278 11098 22330
rect 11098 22278 11110 22330
rect 11110 22278 11132 22330
rect 11156 22278 11162 22330
rect 11162 22278 11174 22330
rect 11174 22278 11212 22330
rect 11236 22278 11238 22330
rect 11238 22278 11290 22330
rect 11290 22278 11292 22330
rect 10916 22276 10972 22278
rect 10996 22276 11052 22278
rect 11076 22276 11132 22278
rect 11156 22276 11212 22278
rect 11236 22276 11292 22278
rect 18916 22330 18972 22332
rect 18996 22330 19052 22332
rect 19076 22330 19132 22332
rect 19156 22330 19212 22332
rect 19236 22330 19292 22332
rect 18916 22278 18918 22330
rect 18918 22278 18970 22330
rect 18970 22278 18972 22330
rect 18996 22278 19034 22330
rect 19034 22278 19046 22330
rect 19046 22278 19052 22330
rect 19076 22278 19098 22330
rect 19098 22278 19110 22330
rect 19110 22278 19132 22330
rect 19156 22278 19162 22330
rect 19162 22278 19174 22330
rect 19174 22278 19212 22330
rect 19236 22278 19238 22330
rect 19238 22278 19290 22330
rect 19290 22278 19292 22330
rect 18916 22276 18972 22278
rect 18996 22276 19052 22278
rect 19076 22276 19132 22278
rect 19156 22276 19212 22278
rect 19236 22276 19292 22278
rect 26916 22330 26972 22332
rect 26996 22330 27052 22332
rect 27076 22330 27132 22332
rect 27156 22330 27212 22332
rect 27236 22330 27292 22332
rect 26916 22278 26918 22330
rect 26918 22278 26970 22330
rect 26970 22278 26972 22330
rect 26996 22278 27034 22330
rect 27034 22278 27046 22330
rect 27046 22278 27052 22330
rect 27076 22278 27098 22330
rect 27098 22278 27110 22330
rect 27110 22278 27132 22330
rect 27156 22278 27162 22330
rect 27162 22278 27174 22330
rect 27174 22278 27212 22330
rect 27236 22278 27238 22330
rect 27238 22278 27290 22330
rect 27290 22278 27292 22330
rect 26916 22276 26972 22278
rect 26996 22276 27052 22278
rect 27076 22276 27132 22278
rect 27156 22276 27212 22278
rect 27236 22276 27292 22278
rect 11656 21786 11712 21788
rect 11736 21786 11792 21788
rect 11816 21786 11872 21788
rect 11896 21786 11952 21788
rect 11976 21786 12032 21788
rect 11656 21734 11658 21786
rect 11658 21734 11710 21786
rect 11710 21734 11712 21786
rect 11736 21734 11774 21786
rect 11774 21734 11786 21786
rect 11786 21734 11792 21786
rect 11816 21734 11838 21786
rect 11838 21734 11850 21786
rect 11850 21734 11872 21786
rect 11896 21734 11902 21786
rect 11902 21734 11914 21786
rect 11914 21734 11952 21786
rect 11976 21734 11978 21786
rect 11978 21734 12030 21786
rect 12030 21734 12032 21786
rect 11656 21732 11712 21734
rect 11736 21732 11792 21734
rect 11816 21732 11872 21734
rect 11896 21732 11952 21734
rect 11976 21732 12032 21734
rect 19656 21786 19712 21788
rect 19736 21786 19792 21788
rect 19816 21786 19872 21788
rect 19896 21786 19952 21788
rect 19976 21786 20032 21788
rect 19656 21734 19658 21786
rect 19658 21734 19710 21786
rect 19710 21734 19712 21786
rect 19736 21734 19774 21786
rect 19774 21734 19786 21786
rect 19786 21734 19792 21786
rect 19816 21734 19838 21786
rect 19838 21734 19850 21786
rect 19850 21734 19872 21786
rect 19896 21734 19902 21786
rect 19902 21734 19914 21786
rect 19914 21734 19952 21786
rect 19976 21734 19978 21786
rect 19978 21734 20030 21786
rect 20030 21734 20032 21786
rect 19656 21732 19712 21734
rect 19736 21732 19792 21734
rect 19816 21732 19872 21734
rect 19896 21732 19952 21734
rect 19976 21732 20032 21734
rect 27656 21786 27712 21788
rect 27736 21786 27792 21788
rect 27816 21786 27872 21788
rect 27896 21786 27952 21788
rect 27976 21786 28032 21788
rect 27656 21734 27658 21786
rect 27658 21734 27710 21786
rect 27710 21734 27712 21786
rect 27736 21734 27774 21786
rect 27774 21734 27786 21786
rect 27786 21734 27792 21786
rect 27816 21734 27838 21786
rect 27838 21734 27850 21786
rect 27850 21734 27872 21786
rect 27896 21734 27902 21786
rect 27902 21734 27914 21786
rect 27914 21734 27952 21786
rect 27976 21734 27978 21786
rect 27978 21734 28030 21786
rect 28030 21734 28032 21786
rect 27656 21732 27712 21734
rect 27736 21732 27792 21734
rect 27816 21732 27872 21734
rect 27896 21732 27952 21734
rect 27976 21732 28032 21734
rect 10916 21242 10972 21244
rect 10996 21242 11052 21244
rect 11076 21242 11132 21244
rect 11156 21242 11212 21244
rect 11236 21242 11292 21244
rect 10916 21190 10918 21242
rect 10918 21190 10970 21242
rect 10970 21190 10972 21242
rect 10996 21190 11034 21242
rect 11034 21190 11046 21242
rect 11046 21190 11052 21242
rect 11076 21190 11098 21242
rect 11098 21190 11110 21242
rect 11110 21190 11132 21242
rect 11156 21190 11162 21242
rect 11162 21190 11174 21242
rect 11174 21190 11212 21242
rect 11236 21190 11238 21242
rect 11238 21190 11290 21242
rect 11290 21190 11292 21242
rect 10916 21188 10972 21190
rect 10996 21188 11052 21190
rect 11076 21188 11132 21190
rect 11156 21188 11212 21190
rect 11236 21188 11292 21190
rect 18916 21242 18972 21244
rect 18996 21242 19052 21244
rect 19076 21242 19132 21244
rect 19156 21242 19212 21244
rect 19236 21242 19292 21244
rect 18916 21190 18918 21242
rect 18918 21190 18970 21242
rect 18970 21190 18972 21242
rect 18996 21190 19034 21242
rect 19034 21190 19046 21242
rect 19046 21190 19052 21242
rect 19076 21190 19098 21242
rect 19098 21190 19110 21242
rect 19110 21190 19132 21242
rect 19156 21190 19162 21242
rect 19162 21190 19174 21242
rect 19174 21190 19212 21242
rect 19236 21190 19238 21242
rect 19238 21190 19290 21242
rect 19290 21190 19292 21242
rect 18916 21188 18972 21190
rect 18996 21188 19052 21190
rect 19076 21188 19132 21190
rect 19156 21188 19212 21190
rect 19236 21188 19292 21190
rect 26916 21242 26972 21244
rect 26996 21242 27052 21244
rect 27076 21242 27132 21244
rect 27156 21242 27212 21244
rect 27236 21242 27292 21244
rect 26916 21190 26918 21242
rect 26918 21190 26970 21242
rect 26970 21190 26972 21242
rect 26996 21190 27034 21242
rect 27034 21190 27046 21242
rect 27046 21190 27052 21242
rect 27076 21190 27098 21242
rect 27098 21190 27110 21242
rect 27110 21190 27132 21242
rect 27156 21190 27162 21242
rect 27162 21190 27174 21242
rect 27174 21190 27212 21242
rect 27236 21190 27238 21242
rect 27238 21190 27290 21242
rect 27290 21190 27292 21242
rect 26916 21188 26972 21190
rect 26996 21188 27052 21190
rect 27076 21188 27132 21190
rect 27156 21188 27212 21190
rect 27236 21188 27292 21190
rect 11656 20698 11712 20700
rect 11736 20698 11792 20700
rect 11816 20698 11872 20700
rect 11896 20698 11952 20700
rect 11976 20698 12032 20700
rect 11656 20646 11658 20698
rect 11658 20646 11710 20698
rect 11710 20646 11712 20698
rect 11736 20646 11774 20698
rect 11774 20646 11786 20698
rect 11786 20646 11792 20698
rect 11816 20646 11838 20698
rect 11838 20646 11850 20698
rect 11850 20646 11872 20698
rect 11896 20646 11902 20698
rect 11902 20646 11914 20698
rect 11914 20646 11952 20698
rect 11976 20646 11978 20698
rect 11978 20646 12030 20698
rect 12030 20646 12032 20698
rect 11656 20644 11712 20646
rect 11736 20644 11792 20646
rect 11816 20644 11872 20646
rect 11896 20644 11952 20646
rect 11976 20644 12032 20646
rect 10916 20154 10972 20156
rect 10996 20154 11052 20156
rect 11076 20154 11132 20156
rect 11156 20154 11212 20156
rect 11236 20154 11292 20156
rect 10916 20102 10918 20154
rect 10918 20102 10970 20154
rect 10970 20102 10972 20154
rect 10996 20102 11034 20154
rect 11034 20102 11046 20154
rect 11046 20102 11052 20154
rect 11076 20102 11098 20154
rect 11098 20102 11110 20154
rect 11110 20102 11132 20154
rect 11156 20102 11162 20154
rect 11162 20102 11174 20154
rect 11174 20102 11212 20154
rect 11236 20102 11238 20154
rect 11238 20102 11290 20154
rect 11290 20102 11292 20154
rect 10916 20100 10972 20102
rect 10996 20100 11052 20102
rect 11076 20100 11132 20102
rect 11156 20100 11212 20102
rect 11236 20100 11292 20102
rect 11656 19610 11712 19612
rect 11736 19610 11792 19612
rect 11816 19610 11872 19612
rect 11896 19610 11952 19612
rect 11976 19610 12032 19612
rect 11656 19558 11658 19610
rect 11658 19558 11710 19610
rect 11710 19558 11712 19610
rect 11736 19558 11774 19610
rect 11774 19558 11786 19610
rect 11786 19558 11792 19610
rect 11816 19558 11838 19610
rect 11838 19558 11850 19610
rect 11850 19558 11872 19610
rect 11896 19558 11902 19610
rect 11902 19558 11914 19610
rect 11914 19558 11952 19610
rect 11976 19558 11978 19610
rect 11978 19558 12030 19610
rect 12030 19558 12032 19610
rect 11656 19556 11712 19558
rect 11736 19556 11792 19558
rect 11816 19556 11872 19558
rect 11896 19556 11952 19558
rect 11976 19556 12032 19558
rect 10916 19066 10972 19068
rect 10996 19066 11052 19068
rect 11076 19066 11132 19068
rect 11156 19066 11212 19068
rect 11236 19066 11292 19068
rect 10916 19014 10918 19066
rect 10918 19014 10970 19066
rect 10970 19014 10972 19066
rect 10996 19014 11034 19066
rect 11034 19014 11046 19066
rect 11046 19014 11052 19066
rect 11076 19014 11098 19066
rect 11098 19014 11110 19066
rect 11110 19014 11132 19066
rect 11156 19014 11162 19066
rect 11162 19014 11174 19066
rect 11174 19014 11212 19066
rect 11236 19014 11238 19066
rect 11238 19014 11290 19066
rect 11290 19014 11292 19066
rect 10916 19012 10972 19014
rect 10996 19012 11052 19014
rect 11076 19012 11132 19014
rect 11156 19012 11212 19014
rect 11236 19012 11292 19014
rect 10916 17978 10972 17980
rect 10996 17978 11052 17980
rect 11076 17978 11132 17980
rect 11156 17978 11212 17980
rect 11236 17978 11292 17980
rect 10916 17926 10918 17978
rect 10918 17926 10970 17978
rect 10970 17926 10972 17978
rect 10996 17926 11034 17978
rect 11034 17926 11046 17978
rect 11046 17926 11052 17978
rect 11076 17926 11098 17978
rect 11098 17926 11110 17978
rect 11110 17926 11132 17978
rect 11156 17926 11162 17978
rect 11162 17926 11174 17978
rect 11174 17926 11212 17978
rect 11236 17926 11238 17978
rect 11238 17926 11290 17978
rect 11290 17926 11292 17978
rect 10916 17924 10972 17926
rect 10996 17924 11052 17926
rect 11076 17924 11132 17926
rect 11156 17924 11212 17926
rect 11236 17924 11292 17926
rect 10916 16890 10972 16892
rect 10996 16890 11052 16892
rect 11076 16890 11132 16892
rect 11156 16890 11212 16892
rect 11236 16890 11292 16892
rect 10916 16838 10918 16890
rect 10918 16838 10970 16890
rect 10970 16838 10972 16890
rect 10996 16838 11034 16890
rect 11034 16838 11046 16890
rect 11046 16838 11052 16890
rect 11076 16838 11098 16890
rect 11098 16838 11110 16890
rect 11110 16838 11132 16890
rect 11156 16838 11162 16890
rect 11162 16838 11174 16890
rect 11174 16838 11212 16890
rect 11236 16838 11238 16890
rect 11238 16838 11290 16890
rect 11290 16838 11292 16890
rect 10916 16836 10972 16838
rect 10996 16836 11052 16838
rect 11076 16836 11132 16838
rect 11156 16836 11212 16838
rect 11236 16836 11292 16838
rect 11656 18522 11712 18524
rect 11736 18522 11792 18524
rect 11816 18522 11872 18524
rect 11896 18522 11952 18524
rect 11976 18522 12032 18524
rect 11656 18470 11658 18522
rect 11658 18470 11710 18522
rect 11710 18470 11712 18522
rect 11736 18470 11774 18522
rect 11774 18470 11786 18522
rect 11786 18470 11792 18522
rect 11816 18470 11838 18522
rect 11838 18470 11850 18522
rect 11850 18470 11872 18522
rect 11896 18470 11902 18522
rect 11902 18470 11914 18522
rect 11914 18470 11952 18522
rect 11976 18470 11978 18522
rect 11978 18470 12030 18522
rect 12030 18470 12032 18522
rect 11656 18468 11712 18470
rect 11736 18468 11792 18470
rect 11816 18468 11872 18470
rect 11896 18468 11952 18470
rect 11976 18468 12032 18470
rect 19656 20698 19712 20700
rect 19736 20698 19792 20700
rect 19816 20698 19872 20700
rect 19896 20698 19952 20700
rect 19976 20698 20032 20700
rect 19656 20646 19658 20698
rect 19658 20646 19710 20698
rect 19710 20646 19712 20698
rect 19736 20646 19774 20698
rect 19774 20646 19786 20698
rect 19786 20646 19792 20698
rect 19816 20646 19838 20698
rect 19838 20646 19850 20698
rect 19850 20646 19872 20698
rect 19896 20646 19902 20698
rect 19902 20646 19914 20698
rect 19914 20646 19952 20698
rect 19976 20646 19978 20698
rect 19978 20646 20030 20698
rect 20030 20646 20032 20698
rect 19656 20644 19712 20646
rect 19736 20644 19792 20646
rect 19816 20644 19872 20646
rect 19896 20644 19952 20646
rect 19976 20644 20032 20646
rect 27656 20698 27712 20700
rect 27736 20698 27792 20700
rect 27816 20698 27872 20700
rect 27896 20698 27952 20700
rect 27976 20698 28032 20700
rect 27656 20646 27658 20698
rect 27658 20646 27710 20698
rect 27710 20646 27712 20698
rect 27736 20646 27774 20698
rect 27774 20646 27786 20698
rect 27786 20646 27792 20698
rect 27816 20646 27838 20698
rect 27838 20646 27850 20698
rect 27850 20646 27872 20698
rect 27896 20646 27902 20698
rect 27902 20646 27914 20698
rect 27914 20646 27952 20698
rect 27976 20646 27978 20698
rect 27978 20646 28030 20698
rect 28030 20646 28032 20698
rect 27656 20644 27712 20646
rect 27736 20644 27792 20646
rect 27816 20644 27872 20646
rect 27896 20644 27952 20646
rect 27976 20644 28032 20646
rect 18916 20154 18972 20156
rect 18996 20154 19052 20156
rect 19076 20154 19132 20156
rect 19156 20154 19212 20156
rect 19236 20154 19292 20156
rect 18916 20102 18918 20154
rect 18918 20102 18970 20154
rect 18970 20102 18972 20154
rect 18996 20102 19034 20154
rect 19034 20102 19046 20154
rect 19046 20102 19052 20154
rect 19076 20102 19098 20154
rect 19098 20102 19110 20154
rect 19110 20102 19132 20154
rect 19156 20102 19162 20154
rect 19162 20102 19174 20154
rect 19174 20102 19212 20154
rect 19236 20102 19238 20154
rect 19238 20102 19290 20154
rect 19290 20102 19292 20154
rect 18916 20100 18972 20102
rect 18996 20100 19052 20102
rect 19076 20100 19132 20102
rect 19156 20100 19212 20102
rect 19236 20100 19292 20102
rect 11656 17434 11712 17436
rect 11736 17434 11792 17436
rect 11816 17434 11872 17436
rect 11896 17434 11952 17436
rect 11976 17434 12032 17436
rect 11656 17382 11658 17434
rect 11658 17382 11710 17434
rect 11710 17382 11712 17434
rect 11736 17382 11774 17434
rect 11774 17382 11786 17434
rect 11786 17382 11792 17434
rect 11816 17382 11838 17434
rect 11838 17382 11850 17434
rect 11850 17382 11872 17434
rect 11896 17382 11902 17434
rect 11902 17382 11914 17434
rect 11914 17382 11952 17434
rect 11976 17382 11978 17434
rect 11978 17382 12030 17434
rect 12030 17382 12032 17434
rect 11656 17380 11712 17382
rect 11736 17380 11792 17382
rect 11816 17380 11872 17382
rect 11896 17380 11952 17382
rect 11976 17380 12032 17382
rect 10916 15802 10972 15804
rect 10996 15802 11052 15804
rect 11076 15802 11132 15804
rect 11156 15802 11212 15804
rect 11236 15802 11292 15804
rect 10916 15750 10918 15802
rect 10918 15750 10970 15802
rect 10970 15750 10972 15802
rect 10996 15750 11034 15802
rect 11034 15750 11046 15802
rect 11046 15750 11052 15802
rect 11076 15750 11098 15802
rect 11098 15750 11110 15802
rect 11110 15750 11132 15802
rect 11156 15750 11162 15802
rect 11162 15750 11174 15802
rect 11174 15750 11212 15802
rect 11236 15750 11238 15802
rect 11238 15750 11290 15802
rect 11290 15750 11292 15802
rect 10916 15748 10972 15750
rect 10996 15748 11052 15750
rect 11076 15748 11132 15750
rect 11156 15748 11212 15750
rect 11236 15748 11292 15750
rect 10916 14714 10972 14716
rect 10996 14714 11052 14716
rect 11076 14714 11132 14716
rect 11156 14714 11212 14716
rect 11236 14714 11292 14716
rect 10916 14662 10918 14714
rect 10918 14662 10970 14714
rect 10970 14662 10972 14714
rect 10996 14662 11034 14714
rect 11034 14662 11046 14714
rect 11046 14662 11052 14714
rect 11076 14662 11098 14714
rect 11098 14662 11110 14714
rect 11110 14662 11132 14714
rect 11156 14662 11162 14714
rect 11162 14662 11174 14714
rect 11174 14662 11212 14714
rect 11236 14662 11238 14714
rect 11238 14662 11290 14714
rect 11290 14662 11292 14714
rect 10916 14660 10972 14662
rect 10996 14660 11052 14662
rect 11076 14660 11132 14662
rect 11156 14660 11212 14662
rect 11236 14660 11292 14662
rect 10916 13626 10972 13628
rect 10996 13626 11052 13628
rect 11076 13626 11132 13628
rect 11156 13626 11212 13628
rect 11236 13626 11292 13628
rect 10916 13574 10918 13626
rect 10918 13574 10970 13626
rect 10970 13574 10972 13626
rect 10996 13574 11034 13626
rect 11034 13574 11046 13626
rect 11046 13574 11052 13626
rect 11076 13574 11098 13626
rect 11098 13574 11110 13626
rect 11110 13574 11132 13626
rect 11156 13574 11162 13626
rect 11162 13574 11174 13626
rect 11174 13574 11212 13626
rect 11236 13574 11238 13626
rect 11238 13574 11290 13626
rect 11290 13574 11292 13626
rect 10916 13572 10972 13574
rect 10996 13572 11052 13574
rect 11076 13572 11132 13574
rect 11156 13572 11212 13574
rect 11236 13572 11292 13574
rect 11656 16346 11712 16348
rect 11736 16346 11792 16348
rect 11816 16346 11872 16348
rect 11896 16346 11952 16348
rect 11976 16346 12032 16348
rect 11656 16294 11658 16346
rect 11658 16294 11710 16346
rect 11710 16294 11712 16346
rect 11736 16294 11774 16346
rect 11774 16294 11786 16346
rect 11786 16294 11792 16346
rect 11816 16294 11838 16346
rect 11838 16294 11850 16346
rect 11850 16294 11872 16346
rect 11896 16294 11902 16346
rect 11902 16294 11914 16346
rect 11914 16294 11952 16346
rect 11976 16294 11978 16346
rect 11978 16294 12030 16346
rect 12030 16294 12032 16346
rect 11656 16292 11712 16294
rect 11736 16292 11792 16294
rect 11816 16292 11872 16294
rect 11896 16292 11952 16294
rect 11976 16292 12032 16294
rect 11656 15258 11712 15260
rect 11736 15258 11792 15260
rect 11816 15258 11872 15260
rect 11896 15258 11952 15260
rect 11976 15258 12032 15260
rect 11656 15206 11658 15258
rect 11658 15206 11710 15258
rect 11710 15206 11712 15258
rect 11736 15206 11774 15258
rect 11774 15206 11786 15258
rect 11786 15206 11792 15258
rect 11816 15206 11838 15258
rect 11838 15206 11850 15258
rect 11850 15206 11872 15258
rect 11896 15206 11902 15258
rect 11902 15206 11914 15258
rect 11914 15206 11952 15258
rect 11976 15206 11978 15258
rect 11978 15206 12030 15258
rect 12030 15206 12032 15258
rect 11656 15204 11712 15206
rect 11736 15204 11792 15206
rect 11816 15204 11872 15206
rect 11896 15204 11952 15206
rect 11976 15204 12032 15206
rect 11656 14170 11712 14172
rect 11736 14170 11792 14172
rect 11816 14170 11872 14172
rect 11896 14170 11952 14172
rect 11976 14170 12032 14172
rect 11656 14118 11658 14170
rect 11658 14118 11710 14170
rect 11710 14118 11712 14170
rect 11736 14118 11774 14170
rect 11774 14118 11786 14170
rect 11786 14118 11792 14170
rect 11816 14118 11838 14170
rect 11838 14118 11850 14170
rect 11850 14118 11872 14170
rect 11896 14118 11902 14170
rect 11902 14118 11914 14170
rect 11914 14118 11952 14170
rect 11976 14118 11978 14170
rect 11978 14118 12030 14170
rect 12030 14118 12032 14170
rect 11656 14116 11712 14118
rect 11736 14116 11792 14118
rect 11816 14116 11872 14118
rect 11896 14116 11952 14118
rect 11976 14116 12032 14118
rect 10916 12538 10972 12540
rect 10996 12538 11052 12540
rect 11076 12538 11132 12540
rect 11156 12538 11212 12540
rect 11236 12538 11292 12540
rect 10916 12486 10918 12538
rect 10918 12486 10970 12538
rect 10970 12486 10972 12538
rect 10996 12486 11034 12538
rect 11034 12486 11046 12538
rect 11046 12486 11052 12538
rect 11076 12486 11098 12538
rect 11098 12486 11110 12538
rect 11110 12486 11132 12538
rect 11156 12486 11162 12538
rect 11162 12486 11174 12538
rect 11174 12486 11212 12538
rect 11236 12486 11238 12538
rect 11238 12486 11290 12538
rect 11290 12486 11292 12538
rect 10916 12484 10972 12486
rect 10996 12484 11052 12486
rect 11076 12484 11132 12486
rect 11156 12484 11212 12486
rect 11236 12484 11292 12486
rect 3656 7642 3712 7644
rect 3736 7642 3792 7644
rect 3816 7642 3872 7644
rect 3896 7642 3952 7644
rect 3976 7642 4032 7644
rect 3656 7590 3658 7642
rect 3658 7590 3710 7642
rect 3710 7590 3712 7642
rect 3736 7590 3774 7642
rect 3774 7590 3786 7642
rect 3786 7590 3792 7642
rect 3816 7590 3838 7642
rect 3838 7590 3850 7642
rect 3850 7590 3872 7642
rect 3896 7590 3902 7642
rect 3902 7590 3914 7642
rect 3914 7590 3952 7642
rect 3976 7590 3978 7642
rect 3978 7590 4030 7642
rect 4030 7590 4032 7642
rect 3656 7588 3712 7590
rect 3736 7588 3792 7590
rect 3816 7588 3872 7590
rect 3896 7588 3952 7590
rect 3976 7588 4032 7590
rect 3656 6554 3712 6556
rect 3736 6554 3792 6556
rect 3816 6554 3872 6556
rect 3896 6554 3952 6556
rect 3976 6554 4032 6556
rect 3656 6502 3658 6554
rect 3658 6502 3710 6554
rect 3710 6502 3712 6554
rect 3736 6502 3774 6554
rect 3774 6502 3786 6554
rect 3786 6502 3792 6554
rect 3816 6502 3838 6554
rect 3838 6502 3850 6554
rect 3850 6502 3872 6554
rect 3896 6502 3902 6554
rect 3902 6502 3914 6554
rect 3914 6502 3952 6554
rect 3976 6502 3978 6554
rect 3978 6502 4030 6554
rect 4030 6502 4032 6554
rect 3656 6500 3712 6502
rect 3736 6500 3792 6502
rect 3816 6500 3872 6502
rect 3896 6500 3952 6502
rect 3976 6500 4032 6502
rect 3656 5466 3712 5468
rect 3736 5466 3792 5468
rect 3816 5466 3872 5468
rect 3896 5466 3952 5468
rect 3976 5466 4032 5468
rect 3656 5414 3658 5466
rect 3658 5414 3710 5466
rect 3710 5414 3712 5466
rect 3736 5414 3774 5466
rect 3774 5414 3786 5466
rect 3786 5414 3792 5466
rect 3816 5414 3838 5466
rect 3838 5414 3850 5466
rect 3850 5414 3872 5466
rect 3896 5414 3902 5466
rect 3902 5414 3914 5466
rect 3914 5414 3952 5466
rect 3976 5414 3978 5466
rect 3978 5414 4030 5466
rect 4030 5414 4032 5466
rect 3656 5412 3712 5414
rect 3736 5412 3792 5414
rect 3816 5412 3872 5414
rect 3896 5412 3952 5414
rect 3976 5412 4032 5414
rect 2916 3834 2972 3836
rect 2996 3834 3052 3836
rect 3076 3834 3132 3836
rect 3156 3834 3212 3836
rect 3236 3834 3292 3836
rect 2916 3782 2918 3834
rect 2918 3782 2970 3834
rect 2970 3782 2972 3834
rect 2996 3782 3034 3834
rect 3034 3782 3046 3834
rect 3046 3782 3052 3834
rect 3076 3782 3098 3834
rect 3098 3782 3110 3834
rect 3110 3782 3132 3834
rect 3156 3782 3162 3834
rect 3162 3782 3174 3834
rect 3174 3782 3212 3834
rect 3236 3782 3238 3834
rect 3238 3782 3290 3834
rect 3290 3782 3292 3834
rect 2916 3780 2972 3782
rect 2996 3780 3052 3782
rect 3076 3780 3132 3782
rect 3156 3780 3212 3782
rect 3236 3780 3292 3782
rect 3656 4378 3712 4380
rect 3736 4378 3792 4380
rect 3816 4378 3872 4380
rect 3896 4378 3952 4380
rect 3976 4378 4032 4380
rect 3656 4326 3658 4378
rect 3658 4326 3710 4378
rect 3710 4326 3712 4378
rect 3736 4326 3774 4378
rect 3774 4326 3786 4378
rect 3786 4326 3792 4378
rect 3816 4326 3838 4378
rect 3838 4326 3850 4378
rect 3850 4326 3872 4378
rect 3896 4326 3902 4378
rect 3902 4326 3914 4378
rect 3914 4326 3952 4378
rect 3976 4326 3978 4378
rect 3978 4326 4030 4378
rect 4030 4326 4032 4378
rect 3656 4324 3712 4326
rect 3736 4324 3792 4326
rect 3816 4324 3872 4326
rect 3896 4324 3952 4326
rect 3976 4324 4032 4326
rect 6182 6180 6238 6216
rect 6182 6160 6184 6180
rect 6184 6160 6236 6180
rect 6236 6160 6238 6180
rect 3656 3290 3712 3292
rect 3736 3290 3792 3292
rect 3816 3290 3872 3292
rect 3896 3290 3952 3292
rect 3976 3290 4032 3292
rect 3656 3238 3658 3290
rect 3658 3238 3710 3290
rect 3710 3238 3712 3290
rect 3736 3238 3774 3290
rect 3774 3238 3786 3290
rect 3786 3238 3792 3290
rect 3816 3238 3838 3290
rect 3838 3238 3850 3290
rect 3850 3238 3872 3290
rect 3896 3238 3902 3290
rect 3902 3238 3914 3290
rect 3914 3238 3952 3290
rect 3976 3238 3978 3290
rect 3978 3238 4030 3290
rect 4030 3238 4032 3290
rect 3656 3236 3712 3238
rect 3736 3236 3792 3238
rect 3816 3236 3872 3238
rect 3896 3236 3952 3238
rect 3976 3236 4032 3238
rect 10916 11450 10972 11452
rect 10996 11450 11052 11452
rect 11076 11450 11132 11452
rect 11156 11450 11212 11452
rect 11236 11450 11292 11452
rect 10916 11398 10918 11450
rect 10918 11398 10970 11450
rect 10970 11398 10972 11450
rect 10996 11398 11034 11450
rect 11034 11398 11046 11450
rect 11046 11398 11052 11450
rect 11076 11398 11098 11450
rect 11098 11398 11110 11450
rect 11110 11398 11132 11450
rect 11156 11398 11162 11450
rect 11162 11398 11174 11450
rect 11174 11398 11212 11450
rect 11236 11398 11238 11450
rect 11238 11398 11290 11450
rect 11290 11398 11292 11450
rect 10916 11396 10972 11398
rect 10996 11396 11052 11398
rect 11076 11396 11132 11398
rect 11156 11396 11212 11398
rect 11236 11396 11292 11398
rect 11656 13082 11712 13084
rect 11736 13082 11792 13084
rect 11816 13082 11872 13084
rect 11896 13082 11952 13084
rect 11976 13082 12032 13084
rect 11656 13030 11658 13082
rect 11658 13030 11710 13082
rect 11710 13030 11712 13082
rect 11736 13030 11774 13082
rect 11774 13030 11786 13082
rect 11786 13030 11792 13082
rect 11816 13030 11838 13082
rect 11838 13030 11850 13082
rect 11850 13030 11872 13082
rect 11896 13030 11902 13082
rect 11902 13030 11914 13082
rect 11914 13030 11952 13082
rect 11976 13030 11978 13082
rect 11978 13030 12030 13082
rect 12030 13030 12032 13082
rect 11656 13028 11712 13030
rect 11736 13028 11792 13030
rect 11816 13028 11872 13030
rect 11896 13028 11952 13030
rect 11976 13028 12032 13030
rect 11656 11994 11712 11996
rect 11736 11994 11792 11996
rect 11816 11994 11872 11996
rect 11896 11994 11952 11996
rect 11976 11994 12032 11996
rect 11656 11942 11658 11994
rect 11658 11942 11710 11994
rect 11710 11942 11712 11994
rect 11736 11942 11774 11994
rect 11774 11942 11786 11994
rect 11786 11942 11792 11994
rect 11816 11942 11838 11994
rect 11838 11942 11850 11994
rect 11850 11942 11872 11994
rect 11896 11942 11902 11994
rect 11902 11942 11914 11994
rect 11914 11942 11952 11994
rect 11976 11942 11978 11994
rect 11978 11942 12030 11994
rect 12030 11942 12032 11994
rect 11656 11940 11712 11942
rect 11736 11940 11792 11942
rect 11816 11940 11872 11942
rect 11896 11940 11952 11942
rect 11976 11940 12032 11942
rect 10916 10362 10972 10364
rect 10996 10362 11052 10364
rect 11076 10362 11132 10364
rect 11156 10362 11212 10364
rect 11236 10362 11292 10364
rect 10916 10310 10918 10362
rect 10918 10310 10970 10362
rect 10970 10310 10972 10362
rect 10996 10310 11034 10362
rect 11034 10310 11046 10362
rect 11046 10310 11052 10362
rect 11076 10310 11098 10362
rect 11098 10310 11110 10362
rect 11110 10310 11132 10362
rect 11156 10310 11162 10362
rect 11162 10310 11174 10362
rect 11174 10310 11212 10362
rect 11236 10310 11238 10362
rect 11238 10310 11290 10362
rect 11290 10310 11292 10362
rect 10916 10308 10972 10310
rect 10996 10308 11052 10310
rect 11076 10308 11132 10310
rect 11156 10308 11212 10310
rect 11236 10308 11292 10310
rect 10916 9274 10972 9276
rect 10996 9274 11052 9276
rect 11076 9274 11132 9276
rect 11156 9274 11212 9276
rect 11236 9274 11292 9276
rect 10916 9222 10918 9274
rect 10918 9222 10970 9274
rect 10970 9222 10972 9274
rect 10996 9222 11034 9274
rect 11034 9222 11046 9274
rect 11046 9222 11052 9274
rect 11076 9222 11098 9274
rect 11098 9222 11110 9274
rect 11110 9222 11132 9274
rect 11156 9222 11162 9274
rect 11162 9222 11174 9274
rect 11174 9222 11212 9274
rect 11236 9222 11238 9274
rect 11238 9222 11290 9274
rect 11290 9222 11292 9274
rect 10916 9220 10972 9222
rect 10996 9220 11052 9222
rect 11076 9220 11132 9222
rect 11156 9220 11212 9222
rect 11236 9220 11292 9222
rect 10916 8186 10972 8188
rect 10996 8186 11052 8188
rect 11076 8186 11132 8188
rect 11156 8186 11212 8188
rect 11236 8186 11292 8188
rect 10916 8134 10918 8186
rect 10918 8134 10970 8186
rect 10970 8134 10972 8186
rect 10996 8134 11034 8186
rect 11034 8134 11046 8186
rect 11046 8134 11052 8186
rect 11076 8134 11098 8186
rect 11098 8134 11110 8186
rect 11110 8134 11132 8186
rect 11156 8134 11162 8186
rect 11162 8134 11174 8186
rect 11174 8134 11212 8186
rect 11236 8134 11238 8186
rect 11238 8134 11290 8186
rect 11290 8134 11292 8186
rect 10916 8132 10972 8134
rect 10996 8132 11052 8134
rect 11076 8132 11132 8134
rect 11156 8132 11212 8134
rect 11236 8132 11292 8134
rect 10916 7098 10972 7100
rect 10996 7098 11052 7100
rect 11076 7098 11132 7100
rect 11156 7098 11212 7100
rect 11236 7098 11292 7100
rect 10916 7046 10918 7098
rect 10918 7046 10970 7098
rect 10970 7046 10972 7098
rect 10996 7046 11034 7098
rect 11034 7046 11046 7098
rect 11046 7046 11052 7098
rect 11076 7046 11098 7098
rect 11098 7046 11110 7098
rect 11110 7046 11132 7098
rect 11156 7046 11162 7098
rect 11162 7046 11174 7098
rect 11174 7046 11212 7098
rect 11236 7046 11238 7098
rect 11238 7046 11290 7098
rect 11290 7046 11292 7098
rect 10916 7044 10972 7046
rect 10996 7044 11052 7046
rect 11076 7044 11132 7046
rect 11156 7044 11212 7046
rect 11236 7044 11292 7046
rect 11656 10906 11712 10908
rect 11736 10906 11792 10908
rect 11816 10906 11872 10908
rect 11896 10906 11952 10908
rect 11976 10906 12032 10908
rect 11656 10854 11658 10906
rect 11658 10854 11710 10906
rect 11710 10854 11712 10906
rect 11736 10854 11774 10906
rect 11774 10854 11786 10906
rect 11786 10854 11792 10906
rect 11816 10854 11838 10906
rect 11838 10854 11850 10906
rect 11850 10854 11872 10906
rect 11896 10854 11902 10906
rect 11902 10854 11914 10906
rect 11914 10854 11952 10906
rect 11976 10854 11978 10906
rect 11978 10854 12030 10906
rect 12030 10854 12032 10906
rect 11656 10852 11712 10854
rect 11736 10852 11792 10854
rect 11816 10852 11872 10854
rect 11896 10852 11952 10854
rect 11976 10852 12032 10854
rect 11656 9818 11712 9820
rect 11736 9818 11792 9820
rect 11816 9818 11872 9820
rect 11896 9818 11952 9820
rect 11976 9818 12032 9820
rect 11656 9766 11658 9818
rect 11658 9766 11710 9818
rect 11710 9766 11712 9818
rect 11736 9766 11774 9818
rect 11774 9766 11786 9818
rect 11786 9766 11792 9818
rect 11816 9766 11838 9818
rect 11838 9766 11850 9818
rect 11850 9766 11872 9818
rect 11896 9766 11902 9818
rect 11902 9766 11914 9818
rect 11914 9766 11952 9818
rect 11976 9766 11978 9818
rect 11978 9766 12030 9818
rect 12030 9766 12032 9818
rect 11656 9764 11712 9766
rect 11736 9764 11792 9766
rect 11816 9764 11872 9766
rect 11896 9764 11952 9766
rect 11976 9764 12032 9766
rect 11656 8730 11712 8732
rect 11736 8730 11792 8732
rect 11816 8730 11872 8732
rect 11896 8730 11952 8732
rect 11976 8730 12032 8732
rect 11656 8678 11658 8730
rect 11658 8678 11710 8730
rect 11710 8678 11712 8730
rect 11736 8678 11774 8730
rect 11774 8678 11786 8730
rect 11786 8678 11792 8730
rect 11816 8678 11838 8730
rect 11838 8678 11850 8730
rect 11850 8678 11872 8730
rect 11896 8678 11902 8730
rect 11902 8678 11914 8730
rect 11914 8678 11952 8730
rect 11976 8678 11978 8730
rect 11978 8678 12030 8730
rect 12030 8678 12032 8730
rect 11656 8676 11712 8678
rect 11736 8676 11792 8678
rect 11816 8676 11872 8678
rect 11896 8676 11952 8678
rect 11976 8676 12032 8678
rect 11656 7642 11712 7644
rect 11736 7642 11792 7644
rect 11816 7642 11872 7644
rect 11896 7642 11952 7644
rect 11976 7642 12032 7644
rect 11656 7590 11658 7642
rect 11658 7590 11710 7642
rect 11710 7590 11712 7642
rect 11736 7590 11774 7642
rect 11774 7590 11786 7642
rect 11786 7590 11792 7642
rect 11816 7590 11838 7642
rect 11838 7590 11850 7642
rect 11850 7590 11872 7642
rect 11896 7590 11902 7642
rect 11902 7590 11914 7642
rect 11914 7590 11952 7642
rect 11976 7590 11978 7642
rect 11978 7590 12030 7642
rect 12030 7590 12032 7642
rect 11656 7588 11712 7590
rect 11736 7588 11792 7590
rect 11816 7588 11872 7590
rect 11896 7588 11952 7590
rect 11976 7588 12032 7590
rect 10916 6010 10972 6012
rect 10996 6010 11052 6012
rect 11076 6010 11132 6012
rect 11156 6010 11212 6012
rect 11236 6010 11292 6012
rect 10916 5958 10918 6010
rect 10918 5958 10970 6010
rect 10970 5958 10972 6010
rect 10996 5958 11034 6010
rect 11034 5958 11046 6010
rect 11046 5958 11052 6010
rect 11076 5958 11098 6010
rect 11098 5958 11110 6010
rect 11110 5958 11132 6010
rect 11156 5958 11162 6010
rect 11162 5958 11174 6010
rect 11174 5958 11212 6010
rect 11236 5958 11238 6010
rect 11238 5958 11290 6010
rect 11290 5958 11292 6010
rect 10916 5956 10972 5958
rect 10996 5956 11052 5958
rect 11076 5956 11132 5958
rect 11156 5956 11212 5958
rect 11236 5956 11292 5958
rect 10916 4922 10972 4924
rect 10996 4922 11052 4924
rect 11076 4922 11132 4924
rect 11156 4922 11212 4924
rect 11236 4922 11292 4924
rect 10916 4870 10918 4922
rect 10918 4870 10970 4922
rect 10970 4870 10972 4922
rect 10996 4870 11034 4922
rect 11034 4870 11046 4922
rect 11046 4870 11052 4922
rect 11076 4870 11098 4922
rect 11098 4870 11110 4922
rect 11110 4870 11132 4922
rect 11156 4870 11162 4922
rect 11162 4870 11174 4922
rect 11174 4870 11212 4922
rect 11236 4870 11238 4922
rect 11238 4870 11290 4922
rect 11290 4870 11292 4922
rect 10916 4868 10972 4870
rect 10996 4868 11052 4870
rect 11076 4868 11132 4870
rect 11156 4868 11212 4870
rect 11236 4868 11292 4870
rect 11656 6554 11712 6556
rect 11736 6554 11792 6556
rect 11816 6554 11872 6556
rect 11896 6554 11952 6556
rect 11976 6554 12032 6556
rect 11656 6502 11658 6554
rect 11658 6502 11710 6554
rect 11710 6502 11712 6554
rect 11736 6502 11774 6554
rect 11774 6502 11786 6554
rect 11786 6502 11792 6554
rect 11816 6502 11838 6554
rect 11838 6502 11850 6554
rect 11850 6502 11872 6554
rect 11896 6502 11902 6554
rect 11902 6502 11914 6554
rect 11914 6502 11952 6554
rect 11976 6502 11978 6554
rect 11978 6502 12030 6554
rect 12030 6502 12032 6554
rect 11656 6500 11712 6502
rect 11736 6500 11792 6502
rect 11816 6500 11872 6502
rect 11896 6500 11952 6502
rect 11976 6500 12032 6502
rect 11656 5466 11712 5468
rect 11736 5466 11792 5468
rect 11816 5466 11872 5468
rect 11896 5466 11952 5468
rect 11976 5466 12032 5468
rect 11656 5414 11658 5466
rect 11658 5414 11710 5466
rect 11710 5414 11712 5466
rect 11736 5414 11774 5466
rect 11774 5414 11786 5466
rect 11786 5414 11792 5466
rect 11816 5414 11838 5466
rect 11838 5414 11850 5466
rect 11850 5414 11872 5466
rect 11896 5414 11902 5466
rect 11902 5414 11914 5466
rect 11914 5414 11952 5466
rect 11976 5414 11978 5466
rect 11978 5414 12030 5466
rect 12030 5414 12032 5466
rect 11656 5412 11712 5414
rect 11736 5412 11792 5414
rect 11816 5412 11872 5414
rect 11896 5412 11952 5414
rect 11976 5412 12032 5414
rect 11656 4378 11712 4380
rect 11736 4378 11792 4380
rect 11816 4378 11872 4380
rect 11896 4378 11952 4380
rect 11976 4378 12032 4380
rect 11656 4326 11658 4378
rect 11658 4326 11710 4378
rect 11710 4326 11712 4378
rect 11736 4326 11774 4378
rect 11774 4326 11786 4378
rect 11786 4326 11792 4378
rect 11816 4326 11838 4378
rect 11838 4326 11850 4378
rect 11850 4326 11872 4378
rect 11896 4326 11902 4378
rect 11902 4326 11914 4378
rect 11914 4326 11952 4378
rect 11976 4326 11978 4378
rect 11978 4326 12030 4378
rect 12030 4326 12032 4378
rect 11656 4324 11712 4326
rect 11736 4324 11792 4326
rect 11816 4324 11872 4326
rect 11896 4324 11952 4326
rect 11976 4324 12032 4326
rect 10916 3834 10972 3836
rect 10996 3834 11052 3836
rect 11076 3834 11132 3836
rect 11156 3834 11212 3836
rect 11236 3834 11292 3836
rect 10916 3782 10918 3834
rect 10918 3782 10970 3834
rect 10970 3782 10972 3834
rect 10996 3782 11034 3834
rect 11034 3782 11046 3834
rect 11046 3782 11052 3834
rect 11076 3782 11098 3834
rect 11098 3782 11110 3834
rect 11110 3782 11132 3834
rect 11156 3782 11162 3834
rect 11162 3782 11174 3834
rect 11174 3782 11212 3834
rect 11236 3782 11238 3834
rect 11238 3782 11290 3834
rect 11290 3782 11292 3834
rect 10916 3780 10972 3782
rect 10996 3780 11052 3782
rect 11076 3780 11132 3782
rect 11156 3780 11212 3782
rect 11236 3780 11292 3782
rect 19656 19610 19712 19612
rect 19736 19610 19792 19612
rect 19816 19610 19872 19612
rect 19896 19610 19952 19612
rect 19976 19610 20032 19612
rect 19656 19558 19658 19610
rect 19658 19558 19710 19610
rect 19710 19558 19712 19610
rect 19736 19558 19774 19610
rect 19774 19558 19786 19610
rect 19786 19558 19792 19610
rect 19816 19558 19838 19610
rect 19838 19558 19850 19610
rect 19850 19558 19872 19610
rect 19896 19558 19902 19610
rect 19902 19558 19914 19610
rect 19914 19558 19952 19610
rect 19976 19558 19978 19610
rect 19978 19558 20030 19610
rect 20030 19558 20032 19610
rect 19656 19556 19712 19558
rect 19736 19556 19792 19558
rect 19816 19556 19872 19558
rect 19896 19556 19952 19558
rect 19976 19556 20032 19558
rect 18916 19066 18972 19068
rect 18996 19066 19052 19068
rect 19076 19066 19132 19068
rect 19156 19066 19212 19068
rect 19236 19066 19292 19068
rect 18916 19014 18918 19066
rect 18918 19014 18970 19066
rect 18970 19014 18972 19066
rect 18996 19014 19034 19066
rect 19034 19014 19046 19066
rect 19046 19014 19052 19066
rect 19076 19014 19098 19066
rect 19098 19014 19110 19066
rect 19110 19014 19132 19066
rect 19156 19014 19162 19066
rect 19162 19014 19174 19066
rect 19174 19014 19212 19066
rect 19236 19014 19238 19066
rect 19238 19014 19290 19066
rect 19290 19014 19292 19066
rect 18916 19012 18972 19014
rect 18996 19012 19052 19014
rect 19076 19012 19132 19014
rect 19156 19012 19212 19014
rect 19236 19012 19292 19014
rect 19656 18522 19712 18524
rect 19736 18522 19792 18524
rect 19816 18522 19872 18524
rect 19896 18522 19952 18524
rect 19976 18522 20032 18524
rect 19656 18470 19658 18522
rect 19658 18470 19710 18522
rect 19710 18470 19712 18522
rect 19736 18470 19774 18522
rect 19774 18470 19786 18522
rect 19786 18470 19792 18522
rect 19816 18470 19838 18522
rect 19838 18470 19850 18522
rect 19850 18470 19872 18522
rect 19896 18470 19902 18522
rect 19902 18470 19914 18522
rect 19914 18470 19952 18522
rect 19976 18470 19978 18522
rect 19978 18470 20030 18522
rect 20030 18470 20032 18522
rect 19656 18468 19712 18470
rect 19736 18468 19792 18470
rect 19816 18468 19872 18470
rect 19896 18468 19952 18470
rect 19976 18468 20032 18470
rect 18916 17978 18972 17980
rect 18996 17978 19052 17980
rect 19076 17978 19132 17980
rect 19156 17978 19212 17980
rect 19236 17978 19292 17980
rect 18916 17926 18918 17978
rect 18918 17926 18970 17978
rect 18970 17926 18972 17978
rect 18996 17926 19034 17978
rect 19034 17926 19046 17978
rect 19046 17926 19052 17978
rect 19076 17926 19098 17978
rect 19098 17926 19110 17978
rect 19110 17926 19132 17978
rect 19156 17926 19162 17978
rect 19162 17926 19174 17978
rect 19174 17926 19212 17978
rect 19236 17926 19238 17978
rect 19238 17926 19290 17978
rect 19290 17926 19292 17978
rect 18916 17924 18972 17926
rect 18996 17924 19052 17926
rect 19076 17924 19132 17926
rect 19156 17924 19212 17926
rect 19236 17924 19292 17926
rect 19656 17434 19712 17436
rect 19736 17434 19792 17436
rect 19816 17434 19872 17436
rect 19896 17434 19952 17436
rect 19976 17434 20032 17436
rect 19656 17382 19658 17434
rect 19658 17382 19710 17434
rect 19710 17382 19712 17434
rect 19736 17382 19774 17434
rect 19774 17382 19786 17434
rect 19786 17382 19792 17434
rect 19816 17382 19838 17434
rect 19838 17382 19850 17434
rect 19850 17382 19872 17434
rect 19896 17382 19902 17434
rect 19902 17382 19914 17434
rect 19914 17382 19952 17434
rect 19976 17382 19978 17434
rect 19978 17382 20030 17434
rect 20030 17382 20032 17434
rect 19656 17380 19712 17382
rect 19736 17380 19792 17382
rect 19816 17380 19872 17382
rect 19896 17380 19952 17382
rect 19976 17380 20032 17382
rect 18916 16890 18972 16892
rect 18996 16890 19052 16892
rect 19076 16890 19132 16892
rect 19156 16890 19212 16892
rect 19236 16890 19292 16892
rect 18916 16838 18918 16890
rect 18918 16838 18970 16890
rect 18970 16838 18972 16890
rect 18996 16838 19034 16890
rect 19034 16838 19046 16890
rect 19046 16838 19052 16890
rect 19076 16838 19098 16890
rect 19098 16838 19110 16890
rect 19110 16838 19132 16890
rect 19156 16838 19162 16890
rect 19162 16838 19174 16890
rect 19174 16838 19212 16890
rect 19236 16838 19238 16890
rect 19238 16838 19290 16890
rect 19290 16838 19292 16890
rect 18916 16836 18972 16838
rect 18996 16836 19052 16838
rect 19076 16836 19132 16838
rect 19156 16836 19212 16838
rect 19236 16836 19292 16838
rect 19656 16346 19712 16348
rect 19736 16346 19792 16348
rect 19816 16346 19872 16348
rect 19896 16346 19952 16348
rect 19976 16346 20032 16348
rect 19656 16294 19658 16346
rect 19658 16294 19710 16346
rect 19710 16294 19712 16346
rect 19736 16294 19774 16346
rect 19774 16294 19786 16346
rect 19786 16294 19792 16346
rect 19816 16294 19838 16346
rect 19838 16294 19850 16346
rect 19850 16294 19872 16346
rect 19896 16294 19902 16346
rect 19902 16294 19914 16346
rect 19914 16294 19952 16346
rect 19976 16294 19978 16346
rect 19978 16294 20030 16346
rect 20030 16294 20032 16346
rect 19656 16292 19712 16294
rect 19736 16292 19792 16294
rect 19816 16292 19872 16294
rect 19896 16292 19952 16294
rect 19976 16292 20032 16294
rect 11656 3290 11712 3292
rect 11736 3290 11792 3292
rect 11816 3290 11872 3292
rect 11896 3290 11952 3292
rect 11976 3290 12032 3292
rect 11656 3238 11658 3290
rect 11658 3238 11710 3290
rect 11710 3238 11712 3290
rect 11736 3238 11774 3290
rect 11774 3238 11786 3290
rect 11786 3238 11792 3290
rect 11816 3238 11838 3290
rect 11838 3238 11850 3290
rect 11850 3238 11872 3290
rect 11896 3238 11902 3290
rect 11902 3238 11914 3290
rect 11914 3238 11952 3290
rect 11976 3238 11978 3290
rect 11978 3238 12030 3290
rect 12030 3238 12032 3290
rect 11656 3236 11712 3238
rect 11736 3236 11792 3238
rect 11816 3236 11872 3238
rect 11896 3236 11952 3238
rect 11976 3236 12032 3238
rect 14278 6160 14334 6216
rect 18916 15802 18972 15804
rect 18996 15802 19052 15804
rect 19076 15802 19132 15804
rect 19156 15802 19212 15804
rect 19236 15802 19292 15804
rect 18916 15750 18918 15802
rect 18918 15750 18970 15802
rect 18970 15750 18972 15802
rect 18996 15750 19034 15802
rect 19034 15750 19046 15802
rect 19046 15750 19052 15802
rect 19076 15750 19098 15802
rect 19098 15750 19110 15802
rect 19110 15750 19132 15802
rect 19156 15750 19162 15802
rect 19162 15750 19174 15802
rect 19174 15750 19212 15802
rect 19236 15750 19238 15802
rect 19238 15750 19290 15802
rect 19290 15750 19292 15802
rect 18916 15748 18972 15750
rect 18996 15748 19052 15750
rect 19076 15748 19132 15750
rect 19156 15748 19212 15750
rect 19236 15748 19292 15750
rect 18916 14714 18972 14716
rect 18996 14714 19052 14716
rect 19076 14714 19132 14716
rect 19156 14714 19212 14716
rect 19236 14714 19292 14716
rect 18916 14662 18918 14714
rect 18918 14662 18970 14714
rect 18970 14662 18972 14714
rect 18996 14662 19034 14714
rect 19034 14662 19046 14714
rect 19046 14662 19052 14714
rect 19076 14662 19098 14714
rect 19098 14662 19110 14714
rect 19110 14662 19132 14714
rect 19156 14662 19162 14714
rect 19162 14662 19174 14714
rect 19174 14662 19212 14714
rect 19236 14662 19238 14714
rect 19238 14662 19290 14714
rect 19290 14662 19292 14714
rect 18916 14660 18972 14662
rect 18996 14660 19052 14662
rect 19076 14660 19132 14662
rect 19156 14660 19212 14662
rect 19236 14660 19292 14662
rect 18916 13626 18972 13628
rect 18996 13626 19052 13628
rect 19076 13626 19132 13628
rect 19156 13626 19212 13628
rect 19236 13626 19292 13628
rect 18916 13574 18918 13626
rect 18918 13574 18970 13626
rect 18970 13574 18972 13626
rect 18996 13574 19034 13626
rect 19034 13574 19046 13626
rect 19046 13574 19052 13626
rect 19076 13574 19098 13626
rect 19098 13574 19110 13626
rect 19110 13574 19132 13626
rect 19156 13574 19162 13626
rect 19162 13574 19174 13626
rect 19174 13574 19212 13626
rect 19236 13574 19238 13626
rect 19238 13574 19290 13626
rect 19290 13574 19292 13626
rect 18916 13572 18972 13574
rect 18996 13572 19052 13574
rect 19076 13572 19132 13574
rect 19156 13572 19212 13574
rect 19236 13572 19292 13574
rect 18916 12538 18972 12540
rect 18996 12538 19052 12540
rect 19076 12538 19132 12540
rect 19156 12538 19212 12540
rect 19236 12538 19292 12540
rect 18916 12486 18918 12538
rect 18918 12486 18970 12538
rect 18970 12486 18972 12538
rect 18996 12486 19034 12538
rect 19034 12486 19046 12538
rect 19046 12486 19052 12538
rect 19076 12486 19098 12538
rect 19098 12486 19110 12538
rect 19110 12486 19132 12538
rect 19156 12486 19162 12538
rect 19162 12486 19174 12538
rect 19174 12486 19212 12538
rect 19236 12486 19238 12538
rect 19238 12486 19290 12538
rect 19290 12486 19292 12538
rect 18916 12484 18972 12486
rect 18996 12484 19052 12486
rect 19076 12484 19132 12486
rect 19156 12484 19212 12486
rect 19236 12484 19292 12486
rect 19656 15258 19712 15260
rect 19736 15258 19792 15260
rect 19816 15258 19872 15260
rect 19896 15258 19952 15260
rect 19976 15258 20032 15260
rect 19656 15206 19658 15258
rect 19658 15206 19710 15258
rect 19710 15206 19712 15258
rect 19736 15206 19774 15258
rect 19774 15206 19786 15258
rect 19786 15206 19792 15258
rect 19816 15206 19838 15258
rect 19838 15206 19850 15258
rect 19850 15206 19872 15258
rect 19896 15206 19902 15258
rect 19902 15206 19914 15258
rect 19914 15206 19952 15258
rect 19976 15206 19978 15258
rect 19978 15206 20030 15258
rect 20030 15206 20032 15258
rect 19656 15204 19712 15206
rect 19736 15204 19792 15206
rect 19816 15204 19872 15206
rect 19896 15204 19952 15206
rect 19976 15204 20032 15206
rect 19656 14170 19712 14172
rect 19736 14170 19792 14172
rect 19816 14170 19872 14172
rect 19896 14170 19952 14172
rect 19976 14170 20032 14172
rect 19656 14118 19658 14170
rect 19658 14118 19710 14170
rect 19710 14118 19712 14170
rect 19736 14118 19774 14170
rect 19774 14118 19786 14170
rect 19786 14118 19792 14170
rect 19816 14118 19838 14170
rect 19838 14118 19850 14170
rect 19850 14118 19872 14170
rect 19896 14118 19902 14170
rect 19902 14118 19914 14170
rect 19914 14118 19952 14170
rect 19976 14118 19978 14170
rect 19978 14118 20030 14170
rect 20030 14118 20032 14170
rect 19656 14116 19712 14118
rect 19736 14116 19792 14118
rect 19816 14116 19872 14118
rect 19896 14116 19952 14118
rect 19976 14116 20032 14118
rect 19656 13082 19712 13084
rect 19736 13082 19792 13084
rect 19816 13082 19872 13084
rect 19896 13082 19952 13084
rect 19976 13082 20032 13084
rect 19656 13030 19658 13082
rect 19658 13030 19710 13082
rect 19710 13030 19712 13082
rect 19736 13030 19774 13082
rect 19774 13030 19786 13082
rect 19786 13030 19792 13082
rect 19816 13030 19838 13082
rect 19838 13030 19850 13082
rect 19850 13030 19872 13082
rect 19896 13030 19902 13082
rect 19902 13030 19914 13082
rect 19914 13030 19952 13082
rect 19976 13030 19978 13082
rect 19978 13030 20030 13082
rect 20030 13030 20032 13082
rect 19656 13028 19712 13030
rect 19736 13028 19792 13030
rect 19816 13028 19872 13030
rect 19896 13028 19952 13030
rect 19976 13028 20032 13030
rect 19656 11994 19712 11996
rect 19736 11994 19792 11996
rect 19816 11994 19872 11996
rect 19896 11994 19952 11996
rect 19976 11994 20032 11996
rect 19656 11942 19658 11994
rect 19658 11942 19710 11994
rect 19710 11942 19712 11994
rect 19736 11942 19774 11994
rect 19774 11942 19786 11994
rect 19786 11942 19792 11994
rect 19816 11942 19838 11994
rect 19838 11942 19850 11994
rect 19850 11942 19872 11994
rect 19896 11942 19902 11994
rect 19902 11942 19914 11994
rect 19914 11942 19952 11994
rect 19976 11942 19978 11994
rect 19978 11942 20030 11994
rect 20030 11942 20032 11994
rect 19656 11940 19712 11942
rect 19736 11940 19792 11942
rect 19816 11940 19872 11942
rect 19896 11940 19952 11942
rect 19976 11940 20032 11942
rect 18916 11450 18972 11452
rect 18996 11450 19052 11452
rect 19076 11450 19132 11452
rect 19156 11450 19212 11452
rect 19236 11450 19292 11452
rect 18916 11398 18918 11450
rect 18918 11398 18970 11450
rect 18970 11398 18972 11450
rect 18996 11398 19034 11450
rect 19034 11398 19046 11450
rect 19046 11398 19052 11450
rect 19076 11398 19098 11450
rect 19098 11398 19110 11450
rect 19110 11398 19132 11450
rect 19156 11398 19162 11450
rect 19162 11398 19174 11450
rect 19174 11398 19212 11450
rect 19236 11398 19238 11450
rect 19238 11398 19290 11450
rect 19290 11398 19292 11450
rect 18916 11396 18972 11398
rect 18996 11396 19052 11398
rect 19076 11396 19132 11398
rect 19156 11396 19212 11398
rect 19236 11396 19292 11398
rect 18916 10362 18972 10364
rect 18996 10362 19052 10364
rect 19076 10362 19132 10364
rect 19156 10362 19212 10364
rect 19236 10362 19292 10364
rect 18916 10310 18918 10362
rect 18918 10310 18970 10362
rect 18970 10310 18972 10362
rect 18996 10310 19034 10362
rect 19034 10310 19046 10362
rect 19046 10310 19052 10362
rect 19076 10310 19098 10362
rect 19098 10310 19110 10362
rect 19110 10310 19132 10362
rect 19156 10310 19162 10362
rect 19162 10310 19174 10362
rect 19174 10310 19212 10362
rect 19236 10310 19238 10362
rect 19238 10310 19290 10362
rect 19290 10310 19292 10362
rect 18916 10308 18972 10310
rect 18996 10308 19052 10310
rect 19076 10308 19132 10310
rect 19156 10308 19212 10310
rect 19236 10308 19292 10310
rect 18916 9274 18972 9276
rect 18996 9274 19052 9276
rect 19076 9274 19132 9276
rect 19156 9274 19212 9276
rect 19236 9274 19292 9276
rect 18916 9222 18918 9274
rect 18918 9222 18970 9274
rect 18970 9222 18972 9274
rect 18996 9222 19034 9274
rect 19034 9222 19046 9274
rect 19046 9222 19052 9274
rect 19076 9222 19098 9274
rect 19098 9222 19110 9274
rect 19110 9222 19132 9274
rect 19156 9222 19162 9274
rect 19162 9222 19174 9274
rect 19174 9222 19212 9274
rect 19236 9222 19238 9274
rect 19238 9222 19290 9274
rect 19290 9222 19292 9274
rect 18916 9220 18972 9222
rect 18996 9220 19052 9222
rect 19076 9220 19132 9222
rect 19156 9220 19212 9222
rect 19236 9220 19292 9222
rect 19656 10906 19712 10908
rect 19736 10906 19792 10908
rect 19816 10906 19872 10908
rect 19896 10906 19952 10908
rect 19976 10906 20032 10908
rect 19656 10854 19658 10906
rect 19658 10854 19710 10906
rect 19710 10854 19712 10906
rect 19736 10854 19774 10906
rect 19774 10854 19786 10906
rect 19786 10854 19792 10906
rect 19816 10854 19838 10906
rect 19838 10854 19850 10906
rect 19850 10854 19872 10906
rect 19896 10854 19902 10906
rect 19902 10854 19914 10906
rect 19914 10854 19952 10906
rect 19976 10854 19978 10906
rect 19978 10854 20030 10906
rect 20030 10854 20032 10906
rect 19656 10852 19712 10854
rect 19736 10852 19792 10854
rect 19816 10852 19872 10854
rect 19896 10852 19952 10854
rect 19976 10852 20032 10854
rect 19656 9818 19712 9820
rect 19736 9818 19792 9820
rect 19816 9818 19872 9820
rect 19896 9818 19952 9820
rect 19976 9818 20032 9820
rect 19656 9766 19658 9818
rect 19658 9766 19710 9818
rect 19710 9766 19712 9818
rect 19736 9766 19774 9818
rect 19774 9766 19786 9818
rect 19786 9766 19792 9818
rect 19816 9766 19838 9818
rect 19838 9766 19850 9818
rect 19850 9766 19872 9818
rect 19896 9766 19902 9818
rect 19902 9766 19914 9818
rect 19914 9766 19952 9818
rect 19976 9766 19978 9818
rect 19978 9766 20030 9818
rect 20030 9766 20032 9818
rect 19656 9764 19712 9766
rect 19736 9764 19792 9766
rect 19816 9764 19872 9766
rect 19896 9764 19952 9766
rect 19976 9764 20032 9766
rect 18916 8186 18972 8188
rect 18996 8186 19052 8188
rect 19076 8186 19132 8188
rect 19156 8186 19212 8188
rect 19236 8186 19292 8188
rect 18916 8134 18918 8186
rect 18918 8134 18970 8186
rect 18970 8134 18972 8186
rect 18996 8134 19034 8186
rect 19034 8134 19046 8186
rect 19046 8134 19052 8186
rect 19076 8134 19098 8186
rect 19098 8134 19110 8186
rect 19110 8134 19132 8186
rect 19156 8134 19162 8186
rect 19162 8134 19174 8186
rect 19174 8134 19212 8186
rect 19236 8134 19238 8186
rect 19238 8134 19290 8186
rect 19290 8134 19292 8186
rect 18916 8132 18972 8134
rect 18996 8132 19052 8134
rect 19076 8132 19132 8134
rect 19156 8132 19212 8134
rect 19236 8132 19292 8134
rect 19656 8730 19712 8732
rect 19736 8730 19792 8732
rect 19816 8730 19872 8732
rect 19896 8730 19952 8732
rect 19976 8730 20032 8732
rect 19656 8678 19658 8730
rect 19658 8678 19710 8730
rect 19710 8678 19712 8730
rect 19736 8678 19774 8730
rect 19774 8678 19786 8730
rect 19786 8678 19792 8730
rect 19816 8678 19838 8730
rect 19838 8678 19850 8730
rect 19850 8678 19872 8730
rect 19896 8678 19902 8730
rect 19902 8678 19914 8730
rect 19914 8678 19952 8730
rect 19976 8678 19978 8730
rect 19978 8678 20030 8730
rect 20030 8678 20032 8730
rect 19656 8676 19712 8678
rect 19736 8676 19792 8678
rect 19816 8676 19872 8678
rect 19896 8676 19952 8678
rect 19976 8676 20032 8678
rect 26916 20154 26972 20156
rect 26996 20154 27052 20156
rect 27076 20154 27132 20156
rect 27156 20154 27212 20156
rect 27236 20154 27292 20156
rect 26916 20102 26918 20154
rect 26918 20102 26970 20154
rect 26970 20102 26972 20154
rect 26996 20102 27034 20154
rect 27034 20102 27046 20154
rect 27046 20102 27052 20154
rect 27076 20102 27098 20154
rect 27098 20102 27110 20154
rect 27110 20102 27132 20154
rect 27156 20102 27162 20154
rect 27162 20102 27174 20154
rect 27174 20102 27212 20154
rect 27236 20102 27238 20154
rect 27238 20102 27290 20154
rect 27290 20102 27292 20154
rect 26916 20100 26972 20102
rect 26996 20100 27052 20102
rect 27076 20100 27132 20102
rect 27156 20100 27212 20102
rect 27236 20100 27292 20102
rect 28354 22344 28410 22400
rect 27656 19610 27712 19612
rect 27736 19610 27792 19612
rect 27816 19610 27872 19612
rect 27896 19610 27952 19612
rect 27976 19610 28032 19612
rect 27656 19558 27658 19610
rect 27658 19558 27710 19610
rect 27710 19558 27712 19610
rect 27736 19558 27774 19610
rect 27774 19558 27786 19610
rect 27786 19558 27792 19610
rect 27816 19558 27838 19610
rect 27838 19558 27850 19610
rect 27850 19558 27872 19610
rect 27896 19558 27902 19610
rect 27902 19558 27914 19610
rect 27914 19558 27952 19610
rect 27976 19558 27978 19610
rect 27978 19558 28030 19610
rect 28030 19558 28032 19610
rect 27656 19556 27712 19558
rect 27736 19556 27792 19558
rect 27816 19556 27872 19558
rect 27896 19556 27952 19558
rect 27976 19556 28032 19558
rect 26916 19066 26972 19068
rect 26996 19066 27052 19068
rect 27076 19066 27132 19068
rect 27156 19066 27212 19068
rect 27236 19066 27292 19068
rect 26916 19014 26918 19066
rect 26918 19014 26970 19066
rect 26970 19014 26972 19066
rect 26996 19014 27034 19066
rect 27034 19014 27046 19066
rect 27046 19014 27052 19066
rect 27076 19014 27098 19066
rect 27098 19014 27110 19066
rect 27110 19014 27132 19066
rect 27156 19014 27162 19066
rect 27162 19014 27174 19066
rect 27174 19014 27212 19066
rect 27236 19014 27238 19066
rect 27238 19014 27290 19066
rect 27290 19014 27292 19066
rect 26916 19012 26972 19014
rect 26996 19012 27052 19014
rect 27076 19012 27132 19014
rect 27156 19012 27212 19014
rect 27236 19012 27292 19014
rect 18916 7098 18972 7100
rect 18996 7098 19052 7100
rect 19076 7098 19132 7100
rect 19156 7098 19212 7100
rect 19236 7098 19292 7100
rect 18916 7046 18918 7098
rect 18918 7046 18970 7098
rect 18970 7046 18972 7098
rect 18996 7046 19034 7098
rect 19034 7046 19046 7098
rect 19046 7046 19052 7098
rect 19076 7046 19098 7098
rect 19098 7046 19110 7098
rect 19110 7046 19132 7098
rect 19156 7046 19162 7098
rect 19162 7046 19174 7098
rect 19174 7046 19212 7098
rect 19236 7046 19238 7098
rect 19238 7046 19290 7098
rect 19290 7046 19292 7098
rect 18916 7044 18972 7046
rect 18996 7044 19052 7046
rect 19076 7044 19132 7046
rect 19156 7044 19212 7046
rect 19236 7044 19292 7046
rect 19656 7642 19712 7644
rect 19736 7642 19792 7644
rect 19816 7642 19872 7644
rect 19896 7642 19952 7644
rect 19976 7642 20032 7644
rect 19656 7590 19658 7642
rect 19658 7590 19710 7642
rect 19710 7590 19712 7642
rect 19736 7590 19774 7642
rect 19774 7590 19786 7642
rect 19786 7590 19792 7642
rect 19816 7590 19838 7642
rect 19838 7590 19850 7642
rect 19850 7590 19872 7642
rect 19896 7590 19902 7642
rect 19902 7590 19914 7642
rect 19914 7590 19952 7642
rect 19976 7590 19978 7642
rect 19978 7590 20030 7642
rect 20030 7590 20032 7642
rect 19656 7588 19712 7590
rect 19736 7588 19792 7590
rect 19816 7588 19872 7590
rect 19896 7588 19952 7590
rect 19976 7588 20032 7590
rect 18916 6010 18972 6012
rect 18996 6010 19052 6012
rect 19076 6010 19132 6012
rect 19156 6010 19212 6012
rect 19236 6010 19292 6012
rect 18916 5958 18918 6010
rect 18918 5958 18970 6010
rect 18970 5958 18972 6010
rect 18996 5958 19034 6010
rect 19034 5958 19046 6010
rect 19046 5958 19052 6010
rect 19076 5958 19098 6010
rect 19098 5958 19110 6010
rect 19110 5958 19132 6010
rect 19156 5958 19162 6010
rect 19162 5958 19174 6010
rect 19174 5958 19212 6010
rect 19236 5958 19238 6010
rect 19238 5958 19290 6010
rect 19290 5958 19292 6010
rect 18916 5956 18972 5958
rect 18996 5956 19052 5958
rect 19076 5956 19132 5958
rect 19156 5956 19212 5958
rect 19236 5956 19292 5958
rect 19656 6554 19712 6556
rect 19736 6554 19792 6556
rect 19816 6554 19872 6556
rect 19896 6554 19952 6556
rect 19976 6554 20032 6556
rect 19656 6502 19658 6554
rect 19658 6502 19710 6554
rect 19710 6502 19712 6554
rect 19736 6502 19774 6554
rect 19774 6502 19786 6554
rect 19786 6502 19792 6554
rect 19816 6502 19838 6554
rect 19838 6502 19850 6554
rect 19850 6502 19872 6554
rect 19896 6502 19902 6554
rect 19902 6502 19914 6554
rect 19914 6502 19952 6554
rect 19976 6502 19978 6554
rect 19978 6502 20030 6554
rect 20030 6502 20032 6554
rect 19656 6500 19712 6502
rect 19736 6500 19792 6502
rect 19816 6500 19872 6502
rect 19896 6500 19952 6502
rect 19976 6500 20032 6502
rect 27656 18522 27712 18524
rect 27736 18522 27792 18524
rect 27816 18522 27872 18524
rect 27896 18522 27952 18524
rect 27976 18522 28032 18524
rect 27656 18470 27658 18522
rect 27658 18470 27710 18522
rect 27710 18470 27712 18522
rect 27736 18470 27774 18522
rect 27774 18470 27786 18522
rect 27786 18470 27792 18522
rect 27816 18470 27838 18522
rect 27838 18470 27850 18522
rect 27850 18470 27872 18522
rect 27896 18470 27902 18522
rect 27902 18470 27914 18522
rect 27914 18470 27952 18522
rect 27976 18470 27978 18522
rect 27978 18470 28030 18522
rect 28030 18470 28032 18522
rect 27656 18468 27712 18470
rect 27736 18468 27792 18470
rect 27816 18468 27872 18470
rect 27896 18468 27952 18470
rect 27976 18468 28032 18470
rect 26916 17978 26972 17980
rect 26996 17978 27052 17980
rect 27076 17978 27132 17980
rect 27156 17978 27212 17980
rect 27236 17978 27292 17980
rect 26916 17926 26918 17978
rect 26918 17926 26970 17978
rect 26970 17926 26972 17978
rect 26996 17926 27034 17978
rect 27034 17926 27046 17978
rect 27046 17926 27052 17978
rect 27076 17926 27098 17978
rect 27098 17926 27110 17978
rect 27110 17926 27132 17978
rect 27156 17926 27162 17978
rect 27162 17926 27174 17978
rect 27174 17926 27212 17978
rect 27236 17926 27238 17978
rect 27238 17926 27290 17978
rect 27290 17926 27292 17978
rect 26916 17924 26972 17926
rect 26996 17924 27052 17926
rect 27076 17924 27132 17926
rect 27156 17924 27212 17926
rect 27236 17924 27292 17926
rect 27656 17434 27712 17436
rect 27736 17434 27792 17436
rect 27816 17434 27872 17436
rect 27896 17434 27952 17436
rect 27976 17434 28032 17436
rect 27656 17382 27658 17434
rect 27658 17382 27710 17434
rect 27710 17382 27712 17434
rect 27736 17382 27774 17434
rect 27774 17382 27786 17434
rect 27786 17382 27792 17434
rect 27816 17382 27838 17434
rect 27838 17382 27850 17434
rect 27850 17382 27872 17434
rect 27896 17382 27902 17434
rect 27902 17382 27914 17434
rect 27914 17382 27952 17434
rect 27976 17382 27978 17434
rect 27978 17382 28030 17434
rect 28030 17382 28032 17434
rect 27656 17380 27712 17382
rect 27736 17380 27792 17382
rect 27816 17380 27872 17382
rect 27896 17380 27952 17382
rect 27976 17380 28032 17382
rect 26916 16890 26972 16892
rect 26996 16890 27052 16892
rect 27076 16890 27132 16892
rect 27156 16890 27212 16892
rect 27236 16890 27292 16892
rect 26916 16838 26918 16890
rect 26918 16838 26970 16890
rect 26970 16838 26972 16890
rect 26996 16838 27034 16890
rect 27034 16838 27046 16890
rect 27046 16838 27052 16890
rect 27076 16838 27098 16890
rect 27098 16838 27110 16890
rect 27110 16838 27132 16890
rect 27156 16838 27162 16890
rect 27162 16838 27174 16890
rect 27174 16838 27212 16890
rect 27236 16838 27238 16890
rect 27238 16838 27290 16890
rect 27290 16838 27292 16890
rect 26916 16836 26972 16838
rect 26996 16836 27052 16838
rect 27076 16836 27132 16838
rect 27156 16836 27212 16838
rect 27236 16836 27292 16838
rect 27656 16346 27712 16348
rect 27736 16346 27792 16348
rect 27816 16346 27872 16348
rect 27896 16346 27952 16348
rect 27976 16346 28032 16348
rect 27656 16294 27658 16346
rect 27658 16294 27710 16346
rect 27710 16294 27712 16346
rect 27736 16294 27774 16346
rect 27774 16294 27786 16346
rect 27786 16294 27792 16346
rect 27816 16294 27838 16346
rect 27838 16294 27850 16346
rect 27850 16294 27872 16346
rect 27896 16294 27902 16346
rect 27902 16294 27914 16346
rect 27914 16294 27952 16346
rect 27976 16294 27978 16346
rect 27978 16294 28030 16346
rect 28030 16294 28032 16346
rect 27656 16292 27712 16294
rect 27736 16292 27792 16294
rect 27816 16292 27872 16294
rect 27896 16292 27952 16294
rect 27976 16292 28032 16294
rect 26916 15802 26972 15804
rect 26996 15802 27052 15804
rect 27076 15802 27132 15804
rect 27156 15802 27212 15804
rect 27236 15802 27292 15804
rect 26916 15750 26918 15802
rect 26918 15750 26970 15802
rect 26970 15750 26972 15802
rect 26996 15750 27034 15802
rect 27034 15750 27046 15802
rect 27046 15750 27052 15802
rect 27076 15750 27098 15802
rect 27098 15750 27110 15802
rect 27110 15750 27132 15802
rect 27156 15750 27162 15802
rect 27162 15750 27174 15802
rect 27174 15750 27212 15802
rect 27236 15750 27238 15802
rect 27238 15750 27290 15802
rect 27290 15750 27292 15802
rect 26916 15748 26972 15750
rect 26996 15748 27052 15750
rect 27076 15748 27132 15750
rect 27156 15748 27212 15750
rect 27236 15748 27292 15750
rect 27656 15258 27712 15260
rect 27736 15258 27792 15260
rect 27816 15258 27872 15260
rect 27896 15258 27952 15260
rect 27976 15258 28032 15260
rect 27656 15206 27658 15258
rect 27658 15206 27710 15258
rect 27710 15206 27712 15258
rect 27736 15206 27774 15258
rect 27774 15206 27786 15258
rect 27786 15206 27792 15258
rect 27816 15206 27838 15258
rect 27838 15206 27850 15258
rect 27850 15206 27872 15258
rect 27896 15206 27902 15258
rect 27902 15206 27914 15258
rect 27914 15206 27952 15258
rect 27976 15206 27978 15258
rect 27978 15206 28030 15258
rect 28030 15206 28032 15258
rect 27656 15204 27712 15206
rect 27736 15204 27792 15206
rect 27816 15204 27872 15206
rect 27896 15204 27952 15206
rect 27976 15204 28032 15206
rect 26916 14714 26972 14716
rect 26996 14714 27052 14716
rect 27076 14714 27132 14716
rect 27156 14714 27212 14716
rect 27236 14714 27292 14716
rect 26916 14662 26918 14714
rect 26918 14662 26970 14714
rect 26970 14662 26972 14714
rect 26996 14662 27034 14714
rect 27034 14662 27046 14714
rect 27046 14662 27052 14714
rect 27076 14662 27098 14714
rect 27098 14662 27110 14714
rect 27110 14662 27132 14714
rect 27156 14662 27162 14714
rect 27162 14662 27174 14714
rect 27174 14662 27212 14714
rect 27236 14662 27238 14714
rect 27238 14662 27290 14714
rect 27290 14662 27292 14714
rect 26916 14660 26972 14662
rect 26996 14660 27052 14662
rect 27076 14660 27132 14662
rect 27156 14660 27212 14662
rect 27236 14660 27292 14662
rect 27656 14170 27712 14172
rect 27736 14170 27792 14172
rect 27816 14170 27872 14172
rect 27896 14170 27952 14172
rect 27976 14170 28032 14172
rect 27656 14118 27658 14170
rect 27658 14118 27710 14170
rect 27710 14118 27712 14170
rect 27736 14118 27774 14170
rect 27774 14118 27786 14170
rect 27786 14118 27792 14170
rect 27816 14118 27838 14170
rect 27838 14118 27850 14170
rect 27850 14118 27872 14170
rect 27896 14118 27902 14170
rect 27902 14118 27914 14170
rect 27914 14118 27952 14170
rect 27976 14118 27978 14170
rect 27978 14118 28030 14170
rect 28030 14118 28032 14170
rect 27656 14116 27712 14118
rect 27736 14116 27792 14118
rect 27816 14116 27872 14118
rect 27896 14116 27952 14118
rect 27976 14116 28032 14118
rect 26916 13626 26972 13628
rect 26996 13626 27052 13628
rect 27076 13626 27132 13628
rect 27156 13626 27212 13628
rect 27236 13626 27292 13628
rect 26916 13574 26918 13626
rect 26918 13574 26970 13626
rect 26970 13574 26972 13626
rect 26996 13574 27034 13626
rect 27034 13574 27046 13626
rect 27046 13574 27052 13626
rect 27076 13574 27098 13626
rect 27098 13574 27110 13626
rect 27110 13574 27132 13626
rect 27156 13574 27162 13626
rect 27162 13574 27174 13626
rect 27174 13574 27212 13626
rect 27236 13574 27238 13626
rect 27238 13574 27290 13626
rect 27290 13574 27292 13626
rect 26916 13572 26972 13574
rect 26996 13572 27052 13574
rect 27076 13572 27132 13574
rect 27156 13572 27212 13574
rect 27236 13572 27292 13574
rect 27656 13082 27712 13084
rect 27736 13082 27792 13084
rect 27816 13082 27872 13084
rect 27896 13082 27952 13084
rect 27976 13082 28032 13084
rect 27656 13030 27658 13082
rect 27658 13030 27710 13082
rect 27710 13030 27712 13082
rect 27736 13030 27774 13082
rect 27774 13030 27786 13082
rect 27786 13030 27792 13082
rect 27816 13030 27838 13082
rect 27838 13030 27850 13082
rect 27850 13030 27872 13082
rect 27896 13030 27902 13082
rect 27902 13030 27914 13082
rect 27914 13030 27952 13082
rect 27976 13030 27978 13082
rect 27978 13030 28030 13082
rect 28030 13030 28032 13082
rect 27656 13028 27712 13030
rect 27736 13028 27792 13030
rect 27816 13028 27872 13030
rect 27896 13028 27952 13030
rect 27976 13028 28032 13030
rect 26916 12538 26972 12540
rect 26996 12538 27052 12540
rect 27076 12538 27132 12540
rect 27156 12538 27212 12540
rect 27236 12538 27292 12540
rect 26916 12486 26918 12538
rect 26918 12486 26970 12538
rect 26970 12486 26972 12538
rect 26996 12486 27034 12538
rect 27034 12486 27046 12538
rect 27046 12486 27052 12538
rect 27076 12486 27098 12538
rect 27098 12486 27110 12538
rect 27110 12486 27132 12538
rect 27156 12486 27162 12538
rect 27162 12486 27174 12538
rect 27174 12486 27212 12538
rect 27236 12486 27238 12538
rect 27238 12486 27290 12538
rect 27290 12486 27292 12538
rect 26916 12484 26972 12486
rect 26996 12484 27052 12486
rect 27076 12484 27132 12486
rect 27156 12484 27212 12486
rect 27236 12484 27292 12486
rect 19656 5466 19712 5468
rect 19736 5466 19792 5468
rect 19816 5466 19872 5468
rect 19896 5466 19952 5468
rect 19976 5466 20032 5468
rect 19656 5414 19658 5466
rect 19658 5414 19710 5466
rect 19710 5414 19712 5466
rect 19736 5414 19774 5466
rect 19774 5414 19786 5466
rect 19786 5414 19792 5466
rect 19816 5414 19838 5466
rect 19838 5414 19850 5466
rect 19850 5414 19872 5466
rect 19896 5414 19902 5466
rect 19902 5414 19914 5466
rect 19914 5414 19952 5466
rect 19976 5414 19978 5466
rect 19978 5414 20030 5466
rect 20030 5414 20032 5466
rect 19656 5412 19712 5414
rect 19736 5412 19792 5414
rect 19816 5412 19872 5414
rect 19896 5412 19952 5414
rect 19976 5412 20032 5414
rect 18916 4922 18972 4924
rect 18996 4922 19052 4924
rect 19076 4922 19132 4924
rect 19156 4922 19212 4924
rect 19236 4922 19292 4924
rect 18916 4870 18918 4922
rect 18918 4870 18970 4922
rect 18970 4870 18972 4922
rect 18996 4870 19034 4922
rect 19034 4870 19046 4922
rect 19046 4870 19052 4922
rect 19076 4870 19098 4922
rect 19098 4870 19110 4922
rect 19110 4870 19132 4922
rect 19156 4870 19162 4922
rect 19162 4870 19174 4922
rect 19174 4870 19212 4922
rect 19236 4870 19238 4922
rect 19238 4870 19290 4922
rect 19290 4870 19292 4922
rect 18916 4868 18972 4870
rect 18996 4868 19052 4870
rect 19076 4868 19132 4870
rect 19156 4868 19212 4870
rect 19236 4868 19292 4870
rect 19656 4378 19712 4380
rect 19736 4378 19792 4380
rect 19816 4378 19872 4380
rect 19896 4378 19952 4380
rect 19976 4378 20032 4380
rect 19656 4326 19658 4378
rect 19658 4326 19710 4378
rect 19710 4326 19712 4378
rect 19736 4326 19774 4378
rect 19774 4326 19786 4378
rect 19786 4326 19792 4378
rect 19816 4326 19838 4378
rect 19838 4326 19850 4378
rect 19850 4326 19872 4378
rect 19896 4326 19902 4378
rect 19902 4326 19914 4378
rect 19914 4326 19952 4378
rect 19976 4326 19978 4378
rect 19978 4326 20030 4378
rect 20030 4326 20032 4378
rect 19656 4324 19712 4326
rect 19736 4324 19792 4326
rect 19816 4324 19872 4326
rect 19896 4324 19952 4326
rect 19976 4324 20032 4326
rect 18916 3834 18972 3836
rect 18996 3834 19052 3836
rect 19076 3834 19132 3836
rect 19156 3834 19212 3836
rect 19236 3834 19292 3836
rect 18916 3782 18918 3834
rect 18918 3782 18970 3834
rect 18970 3782 18972 3834
rect 18996 3782 19034 3834
rect 19034 3782 19046 3834
rect 19046 3782 19052 3834
rect 19076 3782 19098 3834
rect 19098 3782 19110 3834
rect 19110 3782 19132 3834
rect 19156 3782 19162 3834
rect 19162 3782 19174 3834
rect 19174 3782 19212 3834
rect 19236 3782 19238 3834
rect 19238 3782 19290 3834
rect 19290 3782 19292 3834
rect 18916 3780 18972 3782
rect 18996 3780 19052 3782
rect 19076 3780 19132 3782
rect 19156 3780 19212 3782
rect 19236 3780 19292 3782
rect 19656 3290 19712 3292
rect 19736 3290 19792 3292
rect 19816 3290 19872 3292
rect 19896 3290 19952 3292
rect 19976 3290 20032 3292
rect 19656 3238 19658 3290
rect 19658 3238 19710 3290
rect 19710 3238 19712 3290
rect 19736 3238 19774 3290
rect 19774 3238 19786 3290
rect 19786 3238 19792 3290
rect 19816 3238 19838 3290
rect 19838 3238 19850 3290
rect 19850 3238 19872 3290
rect 19896 3238 19902 3290
rect 19902 3238 19914 3290
rect 19914 3238 19952 3290
rect 19976 3238 19978 3290
rect 19978 3238 20030 3290
rect 20030 3238 20032 3290
rect 19656 3236 19712 3238
rect 19736 3236 19792 3238
rect 19816 3236 19872 3238
rect 19896 3236 19952 3238
rect 19976 3236 20032 3238
rect 27656 11994 27712 11996
rect 27736 11994 27792 11996
rect 27816 11994 27872 11996
rect 27896 11994 27952 11996
rect 27976 11994 28032 11996
rect 27656 11942 27658 11994
rect 27658 11942 27710 11994
rect 27710 11942 27712 11994
rect 27736 11942 27774 11994
rect 27774 11942 27786 11994
rect 27786 11942 27792 11994
rect 27816 11942 27838 11994
rect 27838 11942 27850 11994
rect 27850 11942 27872 11994
rect 27896 11942 27902 11994
rect 27902 11942 27914 11994
rect 27914 11942 27952 11994
rect 27976 11942 27978 11994
rect 27978 11942 28030 11994
rect 28030 11942 28032 11994
rect 27656 11940 27712 11942
rect 27736 11940 27792 11942
rect 27816 11940 27872 11942
rect 27896 11940 27952 11942
rect 27976 11940 28032 11942
rect 26916 11450 26972 11452
rect 26996 11450 27052 11452
rect 27076 11450 27132 11452
rect 27156 11450 27212 11452
rect 27236 11450 27292 11452
rect 26916 11398 26918 11450
rect 26918 11398 26970 11450
rect 26970 11398 26972 11450
rect 26996 11398 27034 11450
rect 27034 11398 27046 11450
rect 27046 11398 27052 11450
rect 27076 11398 27098 11450
rect 27098 11398 27110 11450
rect 27110 11398 27132 11450
rect 27156 11398 27162 11450
rect 27162 11398 27174 11450
rect 27174 11398 27212 11450
rect 27236 11398 27238 11450
rect 27238 11398 27290 11450
rect 27290 11398 27292 11450
rect 26916 11396 26972 11398
rect 26996 11396 27052 11398
rect 27076 11396 27132 11398
rect 27156 11396 27212 11398
rect 27236 11396 27292 11398
rect 27656 10906 27712 10908
rect 27736 10906 27792 10908
rect 27816 10906 27872 10908
rect 27896 10906 27952 10908
rect 27976 10906 28032 10908
rect 27656 10854 27658 10906
rect 27658 10854 27710 10906
rect 27710 10854 27712 10906
rect 27736 10854 27774 10906
rect 27774 10854 27786 10906
rect 27786 10854 27792 10906
rect 27816 10854 27838 10906
rect 27838 10854 27850 10906
rect 27850 10854 27872 10906
rect 27896 10854 27902 10906
rect 27902 10854 27914 10906
rect 27914 10854 27952 10906
rect 27976 10854 27978 10906
rect 27978 10854 28030 10906
rect 28030 10854 28032 10906
rect 27656 10852 27712 10854
rect 27736 10852 27792 10854
rect 27816 10852 27872 10854
rect 27896 10852 27952 10854
rect 27976 10852 28032 10854
rect 26916 10362 26972 10364
rect 26996 10362 27052 10364
rect 27076 10362 27132 10364
rect 27156 10362 27212 10364
rect 27236 10362 27292 10364
rect 26916 10310 26918 10362
rect 26918 10310 26970 10362
rect 26970 10310 26972 10362
rect 26996 10310 27034 10362
rect 27034 10310 27046 10362
rect 27046 10310 27052 10362
rect 27076 10310 27098 10362
rect 27098 10310 27110 10362
rect 27110 10310 27132 10362
rect 27156 10310 27162 10362
rect 27162 10310 27174 10362
rect 27174 10310 27212 10362
rect 27236 10310 27238 10362
rect 27238 10310 27290 10362
rect 27290 10310 27292 10362
rect 26916 10308 26972 10310
rect 26996 10308 27052 10310
rect 27076 10308 27132 10310
rect 27156 10308 27212 10310
rect 27236 10308 27292 10310
rect 27656 9818 27712 9820
rect 27736 9818 27792 9820
rect 27816 9818 27872 9820
rect 27896 9818 27952 9820
rect 27976 9818 28032 9820
rect 27656 9766 27658 9818
rect 27658 9766 27710 9818
rect 27710 9766 27712 9818
rect 27736 9766 27774 9818
rect 27774 9766 27786 9818
rect 27786 9766 27792 9818
rect 27816 9766 27838 9818
rect 27838 9766 27850 9818
rect 27850 9766 27872 9818
rect 27896 9766 27902 9818
rect 27902 9766 27914 9818
rect 27914 9766 27952 9818
rect 27976 9766 27978 9818
rect 27978 9766 28030 9818
rect 28030 9766 28032 9818
rect 27656 9764 27712 9766
rect 27736 9764 27792 9766
rect 27816 9764 27872 9766
rect 27896 9764 27952 9766
rect 27976 9764 28032 9766
rect 26916 9274 26972 9276
rect 26996 9274 27052 9276
rect 27076 9274 27132 9276
rect 27156 9274 27212 9276
rect 27236 9274 27292 9276
rect 26916 9222 26918 9274
rect 26918 9222 26970 9274
rect 26970 9222 26972 9274
rect 26996 9222 27034 9274
rect 27034 9222 27046 9274
rect 27046 9222 27052 9274
rect 27076 9222 27098 9274
rect 27098 9222 27110 9274
rect 27110 9222 27132 9274
rect 27156 9222 27162 9274
rect 27162 9222 27174 9274
rect 27174 9222 27212 9274
rect 27236 9222 27238 9274
rect 27238 9222 27290 9274
rect 27290 9222 27292 9274
rect 26916 9220 26972 9222
rect 26996 9220 27052 9222
rect 27076 9220 27132 9222
rect 27156 9220 27212 9222
rect 27236 9220 27292 9222
rect 27656 8730 27712 8732
rect 27736 8730 27792 8732
rect 27816 8730 27872 8732
rect 27896 8730 27952 8732
rect 27976 8730 28032 8732
rect 27656 8678 27658 8730
rect 27658 8678 27710 8730
rect 27710 8678 27712 8730
rect 27736 8678 27774 8730
rect 27774 8678 27786 8730
rect 27786 8678 27792 8730
rect 27816 8678 27838 8730
rect 27838 8678 27850 8730
rect 27850 8678 27872 8730
rect 27896 8678 27902 8730
rect 27902 8678 27914 8730
rect 27914 8678 27952 8730
rect 27976 8678 27978 8730
rect 27978 8678 28030 8730
rect 28030 8678 28032 8730
rect 27656 8676 27712 8678
rect 27736 8676 27792 8678
rect 27816 8676 27872 8678
rect 27896 8676 27952 8678
rect 27976 8676 28032 8678
rect 26916 8186 26972 8188
rect 26996 8186 27052 8188
rect 27076 8186 27132 8188
rect 27156 8186 27212 8188
rect 27236 8186 27292 8188
rect 26916 8134 26918 8186
rect 26918 8134 26970 8186
rect 26970 8134 26972 8186
rect 26996 8134 27034 8186
rect 27034 8134 27046 8186
rect 27046 8134 27052 8186
rect 27076 8134 27098 8186
rect 27098 8134 27110 8186
rect 27110 8134 27132 8186
rect 27156 8134 27162 8186
rect 27162 8134 27174 8186
rect 27174 8134 27212 8186
rect 27236 8134 27238 8186
rect 27238 8134 27290 8186
rect 27290 8134 27292 8186
rect 26916 8132 26972 8134
rect 26996 8132 27052 8134
rect 27076 8132 27132 8134
rect 27156 8132 27212 8134
rect 27236 8132 27292 8134
rect 27656 7642 27712 7644
rect 27736 7642 27792 7644
rect 27816 7642 27872 7644
rect 27896 7642 27952 7644
rect 27976 7642 28032 7644
rect 27656 7590 27658 7642
rect 27658 7590 27710 7642
rect 27710 7590 27712 7642
rect 27736 7590 27774 7642
rect 27774 7590 27786 7642
rect 27786 7590 27792 7642
rect 27816 7590 27838 7642
rect 27838 7590 27850 7642
rect 27850 7590 27872 7642
rect 27896 7590 27902 7642
rect 27902 7590 27914 7642
rect 27914 7590 27952 7642
rect 27976 7590 27978 7642
rect 27978 7590 28030 7642
rect 28030 7590 28032 7642
rect 27656 7588 27712 7590
rect 27736 7588 27792 7590
rect 27816 7588 27872 7590
rect 27896 7588 27952 7590
rect 27976 7588 28032 7590
rect 28354 7384 28410 7440
rect 26916 7098 26972 7100
rect 26996 7098 27052 7100
rect 27076 7098 27132 7100
rect 27156 7098 27212 7100
rect 27236 7098 27292 7100
rect 26916 7046 26918 7098
rect 26918 7046 26970 7098
rect 26970 7046 26972 7098
rect 26996 7046 27034 7098
rect 27034 7046 27046 7098
rect 27046 7046 27052 7098
rect 27076 7046 27098 7098
rect 27098 7046 27110 7098
rect 27110 7046 27132 7098
rect 27156 7046 27162 7098
rect 27162 7046 27174 7098
rect 27174 7046 27212 7098
rect 27236 7046 27238 7098
rect 27238 7046 27290 7098
rect 27290 7046 27292 7098
rect 26916 7044 26972 7046
rect 26996 7044 27052 7046
rect 27076 7044 27132 7046
rect 27156 7044 27212 7046
rect 27236 7044 27292 7046
rect 27656 6554 27712 6556
rect 27736 6554 27792 6556
rect 27816 6554 27872 6556
rect 27896 6554 27952 6556
rect 27976 6554 28032 6556
rect 27656 6502 27658 6554
rect 27658 6502 27710 6554
rect 27710 6502 27712 6554
rect 27736 6502 27774 6554
rect 27774 6502 27786 6554
rect 27786 6502 27792 6554
rect 27816 6502 27838 6554
rect 27838 6502 27850 6554
rect 27850 6502 27872 6554
rect 27896 6502 27902 6554
rect 27902 6502 27914 6554
rect 27914 6502 27952 6554
rect 27976 6502 27978 6554
rect 27978 6502 28030 6554
rect 28030 6502 28032 6554
rect 27656 6500 27712 6502
rect 27736 6500 27792 6502
rect 27816 6500 27872 6502
rect 27896 6500 27952 6502
rect 27976 6500 28032 6502
rect 26916 6010 26972 6012
rect 26996 6010 27052 6012
rect 27076 6010 27132 6012
rect 27156 6010 27212 6012
rect 27236 6010 27292 6012
rect 26916 5958 26918 6010
rect 26918 5958 26970 6010
rect 26970 5958 26972 6010
rect 26996 5958 27034 6010
rect 27034 5958 27046 6010
rect 27046 5958 27052 6010
rect 27076 5958 27098 6010
rect 27098 5958 27110 6010
rect 27110 5958 27132 6010
rect 27156 5958 27162 6010
rect 27162 5958 27174 6010
rect 27174 5958 27212 6010
rect 27236 5958 27238 6010
rect 27238 5958 27290 6010
rect 27290 5958 27292 6010
rect 26916 5956 26972 5958
rect 26996 5956 27052 5958
rect 27076 5956 27132 5958
rect 27156 5956 27212 5958
rect 27236 5956 27292 5958
rect 27656 5466 27712 5468
rect 27736 5466 27792 5468
rect 27816 5466 27872 5468
rect 27896 5466 27952 5468
rect 27976 5466 28032 5468
rect 27656 5414 27658 5466
rect 27658 5414 27710 5466
rect 27710 5414 27712 5466
rect 27736 5414 27774 5466
rect 27774 5414 27786 5466
rect 27786 5414 27792 5466
rect 27816 5414 27838 5466
rect 27838 5414 27850 5466
rect 27850 5414 27872 5466
rect 27896 5414 27902 5466
rect 27902 5414 27914 5466
rect 27914 5414 27952 5466
rect 27976 5414 27978 5466
rect 27978 5414 28030 5466
rect 28030 5414 28032 5466
rect 27656 5412 27712 5414
rect 27736 5412 27792 5414
rect 27816 5412 27872 5414
rect 27896 5412 27952 5414
rect 27976 5412 28032 5414
rect 26916 4922 26972 4924
rect 26996 4922 27052 4924
rect 27076 4922 27132 4924
rect 27156 4922 27212 4924
rect 27236 4922 27292 4924
rect 26916 4870 26918 4922
rect 26918 4870 26970 4922
rect 26970 4870 26972 4922
rect 26996 4870 27034 4922
rect 27034 4870 27046 4922
rect 27046 4870 27052 4922
rect 27076 4870 27098 4922
rect 27098 4870 27110 4922
rect 27110 4870 27132 4922
rect 27156 4870 27162 4922
rect 27162 4870 27174 4922
rect 27174 4870 27212 4922
rect 27236 4870 27238 4922
rect 27238 4870 27290 4922
rect 27290 4870 27292 4922
rect 26916 4868 26972 4870
rect 26996 4868 27052 4870
rect 27076 4868 27132 4870
rect 27156 4868 27212 4870
rect 27236 4868 27292 4870
rect 27656 4378 27712 4380
rect 27736 4378 27792 4380
rect 27816 4378 27872 4380
rect 27896 4378 27952 4380
rect 27976 4378 28032 4380
rect 27656 4326 27658 4378
rect 27658 4326 27710 4378
rect 27710 4326 27712 4378
rect 27736 4326 27774 4378
rect 27774 4326 27786 4378
rect 27786 4326 27792 4378
rect 27816 4326 27838 4378
rect 27838 4326 27850 4378
rect 27850 4326 27872 4378
rect 27896 4326 27902 4378
rect 27902 4326 27914 4378
rect 27914 4326 27952 4378
rect 27976 4326 27978 4378
rect 27978 4326 28030 4378
rect 28030 4326 28032 4378
rect 27656 4324 27712 4326
rect 27736 4324 27792 4326
rect 27816 4324 27872 4326
rect 27896 4324 27952 4326
rect 27976 4324 28032 4326
rect 26916 3834 26972 3836
rect 26996 3834 27052 3836
rect 27076 3834 27132 3836
rect 27156 3834 27212 3836
rect 27236 3834 27292 3836
rect 26916 3782 26918 3834
rect 26918 3782 26970 3834
rect 26970 3782 26972 3834
rect 26996 3782 27034 3834
rect 27034 3782 27046 3834
rect 27046 3782 27052 3834
rect 27076 3782 27098 3834
rect 27098 3782 27110 3834
rect 27110 3782 27132 3834
rect 27156 3782 27162 3834
rect 27162 3782 27174 3834
rect 27174 3782 27212 3834
rect 27236 3782 27238 3834
rect 27238 3782 27290 3834
rect 27290 3782 27292 3834
rect 26916 3780 26972 3782
rect 26996 3780 27052 3782
rect 27076 3780 27132 3782
rect 27156 3780 27212 3782
rect 27236 3780 27292 3782
rect 27656 3290 27712 3292
rect 27736 3290 27792 3292
rect 27816 3290 27872 3292
rect 27896 3290 27952 3292
rect 27976 3290 28032 3292
rect 27656 3238 27658 3290
rect 27658 3238 27710 3290
rect 27710 3238 27712 3290
rect 27736 3238 27774 3290
rect 27774 3238 27786 3290
rect 27786 3238 27792 3290
rect 27816 3238 27838 3290
rect 27838 3238 27850 3290
rect 27850 3238 27872 3290
rect 27896 3238 27902 3290
rect 27902 3238 27914 3290
rect 27914 3238 27952 3290
rect 27976 3238 27978 3290
rect 27978 3238 28030 3290
rect 28030 3238 28032 3290
rect 27656 3236 27712 3238
rect 27736 3236 27792 3238
rect 27816 3236 27872 3238
rect 27896 3236 27952 3238
rect 27976 3236 28032 3238
rect 2916 2746 2972 2748
rect 2996 2746 3052 2748
rect 3076 2746 3132 2748
rect 3156 2746 3212 2748
rect 3236 2746 3292 2748
rect 2916 2694 2918 2746
rect 2918 2694 2970 2746
rect 2970 2694 2972 2746
rect 2996 2694 3034 2746
rect 3034 2694 3046 2746
rect 3046 2694 3052 2746
rect 3076 2694 3098 2746
rect 3098 2694 3110 2746
rect 3110 2694 3132 2746
rect 3156 2694 3162 2746
rect 3162 2694 3174 2746
rect 3174 2694 3212 2746
rect 3236 2694 3238 2746
rect 3238 2694 3290 2746
rect 3290 2694 3292 2746
rect 2916 2692 2972 2694
rect 2996 2692 3052 2694
rect 3076 2692 3132 2694
rect 3156 2692 3212 2694
rect 3236 2692 3292 2694
rect 10916 2746 10972 2748
rect 10996 2746 11052 2748
rect 11076 2746 11132 2748
rect 11156 2746 11212 2748
rect 11236 2746 11292 2748
rect 10916 2694 10918 2746
rect 10918 2694 10970 2746
rect 10970 2694 10972 2746
rect 10996 2694 11034 2746
rect 11034 2694 11046 2746
rect 11046 2694 11052 2746
rect 11076 2694 11098 2746
rect 11098 2694 11110 2746
rect 11110 2694 11132 2746
rect 11156 2694 11162 2746
rect 11162 2694 11174 2746
rect 11174 2694 11212 2746
rect 11236 2694 11238 2746
rect 11238 2694 11290 2746
rect 11290 2694 11292 2746
rect 10916 2692 10972 2694
rect 10996 2692 11052 2694
rect 11076 2692 11132 2694
rect 11156 2692 11212 2694
rect 11236 2692 11292 2694
rect 18916 2746 18972 2748
rect 18996 2746 19052 2748
rect 19076 2746 19132 2748
rect 19156 2746 19212 2748
rect 19236 2746 19292 2748
rect 18916 2694 18918 2746
rect 18918 2694 18970 2746
rect 18970 2694 18972 2746
rect 18996 2694 19034 2746
rect 19034 2694 19046 2746
rect 19046 2694 19052 2746
rect 19076 2694 19098 2746
rect 19098 2694 19110 2746
rect 19110 2694 19132 2746
rect 19156 2694 19162 2746
rect 19162 2694 19174 2746
rect 19174 2694 19212 2746
rect 19236 2694 19238 2746
rect 19238 2694 19290 2746
rect 19290 2694 19292 2746
rect 18916 2692 18972 2694
rect 18996 2692 19052 2694
rect 19076 2692 19132 2694
rect 19156 2692 19212 2694
rect 19236 2692 19292 2694
rect 26916 2746 26972 2748
rect 26996 2746 27052 2748
rect 27076 2746 27132 2748
rect 27156 2746 27212 2748
rect 27236 2746 27292 2748
rect 26916 2694 26918 2746
rect 26918 2694 26970 2746
rect 26970 2694 26972 2746
rect 26996 2694 27034 2746
rect 27034 2694 27046 2746
rect 27046 2694 27052 2746
rect 27076 2694 27098 2746
rect 27098 2694 27110 2746
rect 27110 2694 27132 2746
rect 27156 2694 27162 2746
rect 27162 2694 27174 2746
rect 27174 2694 27212 2746
rect 27236 2694 27238 2746
rect 27238 2694 27290 2746
rect 27290 2694 27292 2746
rect 26916 2692 26972 2694
rect 26996 2692 27052 2694
rect 27076 2692 27132 2694
rect 27156 2692 27212 2694
rect 27236 2692 27292 2694
rect 3656 2202 3712 2204
rect 3736 2202 3792 2204
rect 3816 2202 3872 2204
rect 3896 2202 3952 2204
rect 3976 2202 4032 2204
rect 3656 2150 3658 2202
rect 3658 2150 3710 2202
rect 3710 2150 3712 2202
rect 3736 2150 3774 2202
rect 3774 2150 3786 2202
rect 3786 2150 3792 2202
rect 3816 2150 3838 2202
rect 3838 2150 3850 2202
rect 3850 2150 3872 2202
rect 3896 2150 3902 2202
rect 3902 2150 3914 2202
rect 3914 2150 3952 2202
rect 3976 2150 3978 2202
rect 3978 2150 4030 2202
rect 4030 2150 4032 2202
rect 3656 2148 3712 2150
rect 3736 2148 3792 2150
rect 3816 2148 3872 2150
rect 3896 2148 3952 2150
rect 3976 2148 4032 2150
rect 11656 2202 11712 2204
rect 11736 2202 11792 2204
rect 11816 2202 11872 2204
rect 11896 2202 11952 2204
rect 11976 2202 12032 2204
rect 11656 2150 11658 2202
rect 11658 2150 11710 2202
rect 11710 2150 11712 2202
rect 11736 2150 11774 2202
rect 11774 2150 11786 2202
rect 11786 2150 11792 2202
rect 11816 2150 11838 2202
rect 11838 2150 11850 2202
rect 11850 2150 11872 2202
rect 11896 2150 11902 2202
rect 11902 2150 11914 2202
rect 11914 2150 11952 2202
rect 11976 2150 11978 2202
rect 11978 2150 12030 2202
rect 12030 2150 12032 2202
rect 11656 2148 11712 2150
rect 11736 2148 11792 2150
rect 11816 2148 11872 2150
rect 11896 2148 11952 2150
rect 11976 2148 12032 2150
rect 19656 2202 19712 2204
rect 19736 2202 19792 2204
rect 19816 2202 19872 2204
rect 19896 2202 19952 2204
rect 19976 2202 20032 2204
rect 19656 2150 19658 2202
rect 19658 2150 19710 2202
rect 19710 2150 19712 2202
rect 19736 2150 19774 2202
rect 19774 2150 19786 2202
rect 19786 2150 19792 2202
rect 19816 2150 19838 2202
rect 19838 2150 19850 2202
rect 19850 2150 19872 2202
rect 19896 2150 19902 2202
rect 19902 2150 19914 2202
rect 19914 2150 19952 2202
rect 19976 2150 19978 2202
rect 19978 2150 20030 2202
rect 20030 2150 20032 2202
rect 19656 2148 19712 2150
rect 19736 2148 19792 2150
rect 19816 2148 19872 2150
rect 19896 2148 19952 2150
rect 19976 2148 20032 2150
rect 27656 2202 27712 2204
rect 27736 2202 27792 2204
rect 27816 2202 27872 2204
rect 27896 2202 27952 2204
rect 27976 2202 28032 2204
rect 27656 2150 27658 2202
rect 27658 2150 27710 2202
rect 27710 2150 27712 2202
rect 27736 2150 27774 2202
rect 27774 2150 27786 2202
rect 27786 2150 27792 2202
rect 27816 2150 27838 2202
rect 27838 2150 27850 2202
rect 27850 2150 27872 2202
rect 27896 2150 27902 2202
rect 27902 2150 27914 2202
rect 27914 2150 27952 2202
rect 27976 2150 27978 2202
rect 27978 2150 28030 2202
rect 28030 2150 28032 2202
rect 27656 2148 27712 2150
rect 27736 2148 27792 2150
rect 27816 2148 27872 2150
rect 27896 2148 27952 2150
rect 27976 2148 28032 2150
<< metal3 >>
rect 2906 27776 3302 27777
rect 2906 27712 2912 27776
rect 2976 27712 2992 27776
rect 3056 27712 3072 27776
rect 3136 27712 3152 27776
rect 3216 27712 3232 27776
rect 3296 27712 3302 27776
rect 2906 27711 3302 27712
rect 10906 27776 11302 27777
rect 10906 27712 10912 27776
rect 10976 27712 10992 27776
rect 11056 27712 11072 27776
rect 11136 27712 11152 27776
rect 11216 27712 11232 27776
rect 11296 27712 11302 27776
rect 10906 27711 11302 27712
rect 18906 27776 19302 27777
rect 18906 27712 18912 27776
rect 18976 27712 18992 27776
rect 19056 27712 19072 27776
rect 19136 27712 19152 27776
rect 19216 27712 19232 27776
rect 19296 27712 19302 27776
rect 18906 27711 19302 27712
rect 26906 27776 27302 27777
rect 26906 27712 26912 27776
rect 26976 27712 26992 27776
rect 27056 27712 27072 27776
rect 27136 27712 27152 27776
rect 27216 27712 27232 27776
rect 27296 27712 27302 27776
rect 26906 27711 27302 27712
rect 3646 27232 4042 27233
rect 3646 27168 3652 27232
rect 3716 27168 3732 27232
rect 3796 27168 3812 27232
rect 3876 27168 3892 27232
rect 3956 27168 3972 27232
rect 4036 27168 4042 27232
rect 3646 27167 4042 27168
rect 11646 27232 12042 27233
rect 11646 27168 11652 27232
rect 11716 27168 11732 27232
rect 11796 27168 11812 27232
rect 11876 27168 11892 27232
rect 11956 27168 11972 27232
rect 12036 27168 12042 27232
rect 11646 27167 12042 27168
rect 19646 27232 20042 27233
rect 19646 27168 19652 27232
rect 19716 27168 19732 27232
rect 19796 27168 19812 27232
rect 19876 27168 19892 27232
rect 19956 27168 19972 27232
rect 20036 27168 20042 27232
rect 19646 27167 20042 27168
rect 27646 27232 28042 27233
rect 27646 27168 27652 27232
rect 27716 27168 27732 27232
rect 27796 27168 27812 27232
rect 27876 27168 27892 27232
rect 27956 27168 27972 27232
rect 28036 27168 28042 27232
rect 27646 27167 28042 27168
rect 2906 26688 3302 26689
rect 2906 26624 2912 26688
rect 2976 26624 2992 26688
rect 3056 26624 3072 26688
rect 3136 26624 3152 26688
rect 3216 26624 3232 26688
rect 3296 26624 3302 26688
rect 2906 26623 3302 26624
rect 10906 26688 11302 26689
rect 10906 26624 10912 26688
rect 10976 26624 10992 26688
rect 11056 26624 11072 26688
rect 11136 26624 11152 26688
rect 11216 26624 11232 26688
rect 11296 26624 11302 26688
rect 10906 26623 11302 26624
rect 18906 26688 19302 26689
rect 18906 26624 18912 26688
rect 18976 26624 18992 26688
rect 19056 26624 19072 26688
rect 19136 26624 19152 26688
rect 19216 26624 19232 26688
rect 19296 26624 19302 26688
rect 18906 26623 19302 26624
rect 26906 26688 27302 26689
rect 26906 26624 26912 26688
rect 26976 26624 26992 26688
rect 27056 26624 27072 26688
rect 27136 26624 27152 26688
rect 27216 26624 27232 26688
rect 27296 26624 27302 26688
rect 26906 26623 27302 26624
rect 3646 26144 4042 26145
rect 3646 26080 3652 26144
rect 3716 26080 3732 26144
rect 3796 26080 3812 26144
rect 3876 26080 3892 26144
rect 3956 26080 3972 26144
rect 4036 26080 4042 26144
rect 3646 26079 4042 26080
rect 11646 26144 12042 26145
rect 11646 26080 11652 26144
rect 11716 26080 11732 26144
rect 11796 26080 11812 26144
rect 11876 26080 11892 26144
rect 11956 26080 11972 26144
rect 12036 26080 12042 26144
rect 11646 26079 12042 26080
rect 19646 26144 20042 26145
rect 19646 26080 19652 26144
rect 19716 26080 19732 26144
rect 19796 26080 19812 26144
rect 19876 26080 19892 26144
rect 19956 26080 19972 26144
rect 20036 26080 20042 26144
rect 19646 26079 20042 26080
rect 27646 26144 28042 26145
rect 27646 26080 27652 26144
rect 27716 26080 27732 26144
rect 27796 26080 27812 26144
rect 27876 26080 27892 26144
rect 27956 26080 27972 26144
rect 28036 26080 28042 26144
rect 27646 26079 28042 26080
rect 2906 25600 3302 25601
rect 2906 25536 2912 25600
rect 2976 25536 2992 25600
rect 3056 25536 3072 25600
rect 3136 25536 3152 25600
rect 3216 25536 3232 25600
rect 3296 25536 3302 25600
rect 2906 25535 3302 25536
rect 10906 25600 11302 25601
rect 10906 25536 10912 25600
rect 10976 25536 10992 25600
rect 11056 25536 11072 25600
rect 11136 25536 11152 25600
rect 11216 25536 11232 25600
rect 11296 25536 11302 25600
rect 10906 25535 11302 25536
rect 18906 25600 19302 25601
rect 18906 25536 18912 25600
rect 18976 25536 18992 25600
rect 19056 25536 19072 25600
rect 19136 25536 19152 25600
rect 19216 25536 19232 25600
rect 19296 25536 19302 25600
rect 18906 25535 19302 25536
rect 26906 25600 27302 25601
rect 26906 25536 26912 25600
rect 26976 25536 26992 25600
rect 27056 25536 27072 25600
rect 27136 25536 27152 25600
rect 27216 25536 27232 25600
rect 27296 25536 27302 25600
rect 26906 25535 27302 25536
rect 0 25122 800 25152
rect 1209 25122 1275 25125
rect 0 25120 1275 25122
rect 0 25064 1214 25120
rect 1270 25064 1275 25120
rect 0 25062 1275 25064
rect 0 25032 800 25062
rect 1209 25059 1275 25062
rect 3646 25056 4042 25057
rect 3646 24992 3652 25056
rect 3716 24992 3732 25056
rect 3796 24992 3812 25056
rect 3876 24992 3892 25056
rect 3956 24992 3972 25056
rect 4036 24992 4042 25056
rect 3646 24991 4042 24992
rect 11646 25056 12042 25057
rect 11646 24992 11652 25056
rect 11716 24992 11732 25056
rect 11796 24992 11812 25056
rect 11876 24992 11892 25056
rect 11956 24992 11972 25056
rect 12036 24992 12042 25056
rect 11646 24991 12042 24992
rect 19646 25056 20042 25057
rect 19646 24992 19652 25056
rect 19716 24992 19732 25056
rect 19796 24992 19812 25056
rect 19876 24992 19892 25056
rect 19956 24992 19972 25056
rect 20036 24992 20042 25056
rect 19646 24991 20042 24992
rect 27646 25056 28042 25057
rect 27646 24992 27652 25056
rect 27716 24992 27732 25056
rect 27796 24992 27812 25056
rect 27876 24992 27892 25056
rect 27956 24992 27972 25056
rect 28036 24992 28042 25056
rect 27646 24991 28042 24992
rect 0 24578 800 24608
rect 1301 24578 1367 24581
rect 0 24576 1367 24578
rect 0 24520 1306 24576
rect 1362 24520 1367 24576
rect 0 24518 1367 24520
rect 0 24488 800 24518
rect 1301 24515 1367 24518
rect 2906 24512 3302 24513
rect 2906 24448 2912 24512
rect 2976 24448 2992 24512
rect 3056 24448 3072 24512
rect 3136 24448 3152 24512
rect 3216 24448 3232 24512
rect 3296 24448 3302 24512
rect 2906 24447 3302 24448
rect 10906 24512 11302 24513
rect 10906 24448 10912 24512
rect 10976 24448 10992 24512
rect 11056 24448 11072 24512
rect 11136 24448 11152 24512
rect 11216 24448 11232 24512
rect 11296 24448 11302 24512
rect 10906 24447 11302 24448
rect 18906 24512 19302 24513
rect 18906 24448 18912 24512
rect 18976 24448 18992 24512
rect 19056 24448 19072 24512
rect 19136 24448 19152 24512
rect 19216 24448 19232 24512
rect 19296 24448 19302 24512
rect 18906 24447 19302 24448
rect 26906 24512 27302 24513
rect 26906 24448 26912 24512
rect 26976 24448 26992 24512
rect 27056 24448 27072 24512
rect 27136 24448 27152 24512
rect 27216 24448 27232 24512
rect 27296 24448 27302 24512
rect 26906 24447 27302 24448
rect 0 24034 800 24064
rect 1301 24034 1367 24037
rect 0 24032 1367 24034
rect 0 23976 1306 24032
rect 1362 23976 1367 24032
rect 0 23974 1367 23976
rect 0 23944 800 23974
rect 1301 23971 1367 23974
rect 3646 23968 4042 23969
rect 3646 23904 3652 23968
rect 3716 23904 3732 23968
rect 3796 23904 3812 23968
rect 3876 23904 3892 23968
rect 3956 23904 3972 23968
rect 4036 23904 4042 23968
rect 3646 23903 4042 23904
rect 11646 23968 12042 23969
rect 11646 23904 11652 23968
rect 11716 23904 11732 23968
rect 11796 23904 11812 23968
rect 11876 23904 11892 23968
rect 11956 23904 11972 23968
rect 12036 23904 12042 23968
rect 11646 23903 12042 23904
rect 19646 23968 20042 23969
rect 19646 23904 19652 23968
rect 19716 23904 19732 23968
rect 19796 23904 19812 23968
rect 19876 23904 19892 23968
rect 19956 23904 19972 23968
rect 20036 23904 20042 23968
rect 19646 23903 20042 23904
rect 27646 23968 28042 23969
rect 27646 23904 27652 23968
rect 27716 23904 27732 23968
rect 27796 23904 27812 23968
rect 27876 23904 27892 23968
rect 27956 23904 27972 23968
rect 28036 23904 28042 23968
rect 27646 23903 28042 23904
rect 0 23490 800 23520
rect 1301 23490 1367 23493
rect 0 23488 1367 23490
rect 0 23432 1306 23488
rect 1362 23432 1367 23488
rect 0 23430 1367 23432
rect 0 23400 800 23430
rect 1301 23427 1367 23430
rect 2906 23424 3302 23425
rect 2906 23360 2912 23424
rect 2976 23360 2992 23424
rect 3056 23360 3072 23424
rect 3136 23360 3152 23424
rect 3216 23360 3232 23424
rect 3296 23360 3302 23424
rect 2906 23359 3302 23360
rect 10906 23424 11302 23425
rect 10906 23360 10912 23424
rect 10976 23360 10992 23424
rect 11056 23360 11072 23424
rect 11136 23360 11152 23424
rect 11216 23360 11232 23424
rect 11296 23360 11302 23424
rect 10906 23359 11302 23360
rect 18906 23424 19302 23425
rect 18906 23360 18912 23424
rect 18976 23360 18992 23424
rect 19056 23360 19072 23424
rect 19136 23360 19152 23424
rect 19216 23360 19232 23424
rect 19296 23360 19302 23424
rect 18906 23359 19302 23360
rect 26906 23424 27302 23425
rect 26906 23360 26912 23424
rect 26976 23360 26992 23424
rect 27056 23360 27072 23424
rect 27136 23360 27152 23424
rect 27216 23360 27232 23424
rect 27296 23360 27302 23424
rect 26906 23359 27302 23360
rect 3785 23082 3851 23085
rect 3785 23080 4170 23082
rect 3785 23024 3790 23080
rect 3846 23024 4170 23080
rect 3785 23022 4170 23024
rect 3785 23019 3851 23022
rect 0 22946 800 22976
rect 1393 22946 1459 22949
rect 0 22944 1459 22946
rect 0 22888 1398 22944
rect 1454 22888 1459 22944
rect 0 22886 1459 22888
rect 0 22856 800 22886
rect 1393 22883 1459 22886
rect 3646 22880 4042 22881
rect 3646 22816 3652 22880
rect 3716 22816 3732 22880
rect 3796 22816 3812 22880
rect 3876 22816 3892 22880
rect 3956 22816 3972 22880
rect 4036 22816 4042 22880
rect 3646 22815 4042 22816
rect 4110 22541 4170 23022
rect 11646 22880 12042 22881
rect 11646 22816 11652 22880
rect 11716 22816 11732 22880
rect 11796 22816 11812 22880
rect 11876 22816 11892 22880
rect 11956 22816 11972 22880
rect 12036 22816 12042 22880
rect 11646 22815 12042 22816
rect 19646 22880 20042 22881
rect 19646 22816 19652 22880
rect 19716 22816 19732 22880
rect 19796 22816 19812 22880
rect 19876 22816 19892 22880
rect 19956 22816 19972 22880
rect 20036 22816 20042 22880
rect 19646 22815 20042 22816
rect 27646 22880 28042 22881
rect 27646 22816 27652 22880
rect 27716 22816 27732 22880
rect 27796 22816 27812 22880
rect 27876 22816 27892 22880
rect 27956 22816 27972 22880
rect 28036 22816 28042 22880
rect 27646 22815 28042 22816
rect 4061 22536 4170 22541
rect 4061 22480 4066 22536
rect 4122 22480 4170 22536
rect 4061 22478 4170 22480
rect 4061 22475 4127 22478
rect 0 22402 800 22432
rect 1209 22402 1275 22405
rect 0 22400 1275 22402
rect 0 22344 1214 22400
rect 1270 22344 1275 22400
rect 0 22342 1275 22344
rect 0 22312 800 22342
rect 1209 22339 1275 22342
rect 28349 22402 28415 22405
rect 29200 22402 30000 22432
rect 28349 22400 30000 22402
rect 28349 22344 28354 22400
rect 28410 22344 30000 22400
rect 28349 22342 30000 22344
rect 28349 22339 28415 22342
rect 2906 22336 3302 22337
rect 2906 22272 2912 22336
rect 2976 22272 2992 22336
rect 3056 22272 3072 22336
rect 3136 22272 3152 22336
rect 3216 22272 3232 22336
rect 3296 22272 3302 22336
rect 2906 22271 3302 22272
rect 10906 22336 11302 22337
rect 10906 22272 10912 22336
rect 10976 22272 10992 22336
rect 11056 22272 11072 22336
rect 11136 22272 11152 22336
rect 11216 22272 11232 22336
rect 11296 22272 11302 22336
rect 10906 22271 11302 22272
rect 18906 22336 19302 22337
rect 18906 22272 18912 22336
rect 18976 22272 18992 22336
rect 19056 22272 19072 22336
rect 19136 22272 19152 22336
rect 19216 22272 19232 22336
rect 19296 22272 19302 22336
rect 18906 22271 19302 22272
rect 26906 22336 27302 22337
rect 26906 22272 26912 22336
rect 26976 22272 26992 22336
rect 27056 22272 27072 22336
rect 27136 22272 27152 22336
rect 27216 22272 27232 22336
rect 27296 22272 27302 22336
rect 29200 22312 30000 22342
rect 26906 22271 27302 22272
rect 3366 21932 3372 21996
rect 3436 21994 3442 21996
rect 3969 21994 4035 21997
rect 3436 21992 4035 21994
rect 3436 21936 3974 21992
rect 4030 21936 4035 21992
rect 3436 21934 4035 21936
rect 3436 21932 3442 21934
rect 3969 21931 4035 21934
rect 0 21858 800 21888
rect 1209 21858 1275 21861
rect 0 21856 1275 21858
rect 0 21800 1214 21856
rect 1270 21800 1275 21856
rect 0 21798 1275 21800
rect 0 21768 800 21798
rect 1209 21795 1275 21798
rect 3646 21792 4042 21793
rect 3646 21728 3652 21792
rect 3716 21728 3732 21792
rect 3796 21728 3812 21792
rect 3876 21728 3892 21792
rect 3956 21728 3972 21792
rect 4036 21728 4042 21792
rect 3646 21727 4042 21728
rect 11646 21792 12042 21793
rect 11646 21728 11652 21792
rect 11716 21728 11732 21792
rect 11796 21728 11812 21792
rect 11876 21728 11892 21792
rect 11956 21728 11972 21792
rect 12036 21728 12042 21792
rect 11646 21727 12042 21728
rect 19646 21792 20042 21793
rect 19646 21728 19652 21792
rect 19716 21728 19732 21792
rect 19796 21728 19812 21792
rect 19876 21728 19892 21792
rect 19956 21728 19972 21792
rect 20036 21728 20042 21792
rect 19646 21727 20042 21728
rect 27646 21792 28042 21793
rect 27646 21728 27652 21792
rect 27716 21728 27732 21792
rect 27796 21728 27812 21792
rect 27876 21728 27892 21792
rect 27956 21728 27972 21792
rect 28036 21728 28042 21792
rect 27646 21727 28042 21728
rect 0 21314 800 21344
rect 1301 21314 1367 21317
rect 0 21312 1367 21314
rect 0 21256 1306 21312
rect 1362 21256 1367 21312
rect 0 21254 1367 21256
rect 0 21224 800 21254
rect 1301 21251 1367 21254
rect 1710 21252 1716 21316
rect 1780 21314 1786 21316
rect 2405 21314 2471 21317
rect 1780 21312 2471 21314
rect 1780 21256 2410 21312
rect 2466 21256 2471 21312
rect 1780 21254 2471 21256
rect 1780 21252 1786 21254
rect 2405 21251 2471 21254
rect 2906 21248 3302 21249
rect 2906 21184 2912 21248
rect 2976 21184 2992 21248
rect 3056 21184 3072 21248
rect 3136 21184 3152 21248
rect 3216 21184 3232 21248
rect 3296 21184 3302 21248
rect 2906 21183 3302 21184
rect 10906 21248 11302 21249
rect 10906 21184 10912 21248
rect 10976 21184 10992 21248
rect 11056 21184 11072 21248
rect 11136 21184 11152 21248
rect 11216 21184 11232 21248
rect 11296 21184 11302 21248
rect 10906 21183 11302 21184
rect 18906 21248 19302 21249
rect 18906 21184 18912 21248
rect 18976 21184 18992 21248
rect 19056 21184 19072 21248
rect 19136 21184 19152 21248
rect 19216 21184 19232 21248
rect 19296 21184 19302 21248
rect 18906 21183 19302 21184
rect 26906 21248 27302 21249
rect 26906 21184 26912 21248
rect 26976 21184 26992 21248
rect 27056 21184 27072 21248
rect 27136 21184 27152 21248
rect 27216 21184 27232 21248
rect 27296 21184 27302 21248
rect 26906 21183 27302 21184
rect 0 20770 800 20800
rect 1301 20770 1367 20773
rect 0 20768 1367 20770
rect 0 20712 1306 20768
rect 1362 20712 1367 20768
rect 0 20710 1367 20712
rect 0 20680 800 20710
rect 1301 20707 1367 20710
rect 1577 20770 1643 20773
rect 2630 20770 2636 20772
rect 1577 20768 2636 20770
rect 1577 20712 1582 20768
rect 1638 20712 2636 20768
rect 1577 20710 2636 20712
rect 1577 20707 1643 20710
rect 2630 20708 2636 20710
rect 2700 20708 2706 20772
rect 3646 20704 4042 20705
rect 3646 20640 3652 20704
rect 3716 20640 3732 20704
rect 3796 20640 3812 20704
rect 3876 20640 3892 20704
rect 3956 20640 3972 20704
rect 4036 20640 4042 20704
rect 3646 20639 4042 20640
rect 11646 20704 12042 20705
rect 11646 20640 11652 20704
rect 11716 20640 11732 20704
rect 11796 20640 11812 20704
rect 11876 20640 11892 20704
rect 11956 20640 11972 20704
rect 12036 20640 12042 20704
rect 11646 20639 12042 20640
rect 19646 20704 20042 20705
rect 19646 20640 19652 20704
rect 19716 20640 19732 20704
rect 19796 20640 19812 20704
rect 19876 20640 19892 20704
rect 19956 20640 19972 20704
rect 20036 20640 20042 20704
rect 19646 20639 20042 20640
rect 27646 20704 28042 20705
rect 27646 20640 27652 20704
rect 27716 20640 27732 20704
rect 27796 20640 27812 20704
rect 27876 20640 27892 20704
rect 27956 20640 27972 20704
rect 28036 20640 28042 20704
rect 27646 20639 28042 20640
rect 2957 20362 3023 20365
rect 2638 20360 3023 20362
rect 2638 20304 2962 20360
rect 3018 20304 3023 20360
rect 2638 20302 3023 20304
rect 0 20226 800 20256
rect 1301 20226 1367 20229
rect 0 20224 1367 20226
rect 0 20168 1306 20224
rect 1362 20168 1367 20224
rect 0 20166 1367 20168
rect 0 20136 800 20166
rect 1301 20163 1367 20166
rect 2638 19954 2698 20302
rect 2957 20299 3023 20302
rect 2906 20160 3302 20161
rect 2906 20096 2912 20160
rect 2976 20096 2992 20160
rect 3056 20096 3072 20160
rect 3136 20096 3152 20160
rect 3216 20096 3232 20160
rect 3296 20096 3302 20160
rect 2906 20095 3302 20096
rect 10906 20160 11302 20161
rect 10906 20096 10912 20160
rect 10976 20096 10992 20160
rect 11056 20096 11072 20160
rect 11136 20096 11152 20160
rect 11216 20096 11232 20160
rect 11296 20096 11302 20160
rect 10906 20095 11302 20096
rect 18906 20160 19302 20161
rect 18906 20096 18912 20160
rect 18976 20096 18992 20160
rect 19056 20096 19072 20160
rect 19136 20096 19152 20160
rect 19216 20096 19232 20160
rect 19296 20096 19302 20160
rect 18906 20095 19302 20096
rect 26906 20160 27302 20161
rect 26906 20096 26912 20160
rect 26976 20096 26992 20160
rect 27056 20096 27072 20160
rect 27136 20096 27152 20160
rect 27216 20096 27232 20160
rect 27296 20096 27302 20160
rect 26906 20095 27302 20096
rect 2957 19954 3023 19957
rect 2638 19952 3023 19954
rect 2638 19896 2962 19952
rect 3018 19896 3023 19952
rect 2638 19894 3023 19896
rect 2957 19891 3023 19894
rect 0 19682 800 19712
rect 1301 19682 1367 19685
rect 0 19680 1367 19682
rect 0 19624 1306 19680
rect 1362 19624 1367 19680
rect 0 19622 1367 19624
rect 0 19592 800 19622
rect 1301 19619 1367 19622
rect 3646 19616 4042 19617
rect 3646 19552 3652 19616
rect 3716 19552 3732 19616
rect 3796 19552 3812 19616
rect 3876 19552 3892 19616
rect 3956 19552 3972 19616
rect 4036 19552 4042 19616
rect 3646 19551 4042 19552
rect 11646 19616 12042 19617
rect 11646 19552 11652 19616
rect 11716 19552 11732 19616
rect 11796 19552 11812 19616
rect 11876 19552 11892 19616
rect 11956 19552 11972 19616
rect 12036 19552 12042 19616
rect 11646 19551 12042 19552
rect 19646 19616 20042 19617
rect 19646 19552 19652 19616
rect 19716 19552 19732 19616
rect 19796 19552 19812 19616
rect 19876 19552 19892 19616
rect 19956 19552 19972 19616
rect 20036 19552 20042 19616
rect 19646 19551 20042 19552
rect 27646 19616 28042 19617
rect 27646 19552 27652 19616
rect 27716 19552 27732 19616
rect 27796 19552 27812 19616
rect 27876 19552 27892 19616
rect 27956 19552 27972 19616
rect 28036 19552 28042 19616
rect 27646 19551 28042 19552
rect 2078 19348 2084 19412
rect 2148 19410 2154 19412
rect 2865 19410 2931 19413
rect 3366 19410 3372 19412
rect 2148 19408 3372 19410
rect 2148 19352 2870 19408
rect 2926 19352 3372 19408
rect 2148 19350 3372 19352
rect 2148 19348 2154 19350
rect 2865 19347 2931 19350
rect 3366 19348 3372 19350
rect 3436 19348 3442 19412
rect 3877 19410 3943 19413
rect 4245 19410 4311 19413
rect 5809 19410 5875 19413
rect 3877 19408 5875 19410
rect 3877 19352 3882 19408
rect 3938 19352 4250 19408
rect 4306 19352 5814 19408
rect 5870 19352 5875 19408
rect 3877 19350 5875 19352
rect 3877 19347 3943 19350
rect 4245 19347 4311 19350
rect 5809 19347 5875 19350
rect 2589 19274 2655 19277
rect 5625 19274 5691 19277
rect 2589 19272 5691 19274
rect 2589 19216 2594 19272
rect 2650 19216 5630 19272
rect 5686 19216 5691 19272
rect 2589 19214 5691 19216
rect 2589 19211 2655 19214
rect 5625 19211 5691 19214
rect 0 19138 800 19168
rect 1393 19138 1459 19141
rect 0 19136 1459 19138
rect 0 19080 1398 19136
rect 1454 19080 1459 19136
rect 0 19078 1459 19080
rect 0 19048 800 19078
rect 1393 19075 1459 19078
rect 2906 19072 3302 19073
rect 2906 19008 2912 19072
rect 2976 19008 2992 19072
rect 3056 19008 3072 19072
rect 3136 19008 3152 19072
rect 3216 19008 3232 19072
rect 3296 19008 3302 19072
rect 2906 19007 3302 19008
rect 10906 19072 11302 19073
rect 10906 19008 10912 19072
rect 10976 19008 10992 19072
rect 11056 19008 11072 19072
rect 11136 19008 11152 19072
rect 11216 19008 11232 19072
rect 11296 19008 11302 19072
rect 10906 19007 11302 19008
rect 18906 19072 19302 19073
rect 18906 19008 18912 19072
rect 18976 19008 18992 19072
rect 19056 19008 19072 19072
rect 19136 19008 19152 19072
rect 19216 19008 19232 19072
rect 19296 19008 19302 19072
rect 18906 19007 19302 19008
rect 26906 19072 27302 19073
rect 26906 19008 26912 19072
rect 26976 19008 26992 19072
rect 27056 19008 27072 19072
rect 27136 19008 27152 19072
rect 27216 19008 27232 19072
rect 27296 19008 27302 19072
rect 26906 19007 27302 19008
rect 3049 18866 3115 18869
rect 3693 18866 3759 18869
rect 3049 18864 3759 18866
rect 3049 18808 3054 18864
rect 3110 18808 3698 18864
rect 3754 18808 3759 18864
rect 3049 18806 3759 18808
rect 3049 18803 3115 18806
rect 3693 18803 3759 18806
rect 3325 18730 3391 18733
rect 3877 18730 3943 18733
rect 3325 18728 3943 18730
rect 3325 18672 3330 18728
rect 3386 18672 3882 18728
rect 3938 18672 3943 18728
rect 3325 18670 3943 18672
rect 3325 18667 3391 18670
rect 3877 18667 3943 18670
rect 0 18594 800 18624
rect 1301 18594 1367 18597
rect 0 18592 1367 18594
rect 0 18536 1306 18592
rect 1362 18536 1367 18592
rect 0 18534 1367 18536
rect 0 18504 800 18534
rect 1301 18531 1367 18534
rect 3646 18528 4042 18529
rect 3646 18464 3652 18528
rect 3716 18464 3732 18528
rect 3796 18464 3812 18528
rect 3876 18464 3892 18528
rect 3956 18464 3972 18528
rect 4036 18464 4042 18528
rect 3646 18463 4042 18464
rect 11646 18528 12042 18529
rect 11646 18464 11652 18528
rect 11716 18464 11732 18528
rect 11796 18464 11812 18528
rect 11876 18464 11892 18528
rect 11956 18464 11972 18528
rect 12036 18464 12042 18528
rect 11646 18463 12042 18464
rect 19646 18528 20042 18529
rect 19646 18464 19652 18528
rect 19716 18464 19732 18528
rect 19796 18464 19812 18528
rect 19876 18464 19892 18528
rect 19956 18464 19972 18528
rect 20036 18464 20042 18528
rect 19646 18463 20042 18464
rect 27646 18528 28042 18529
rect 27646 18464 27652 18528
rect 27716 18464 27732 18528
rect 27796 18464 27812 18528
rect 27876 18464 27892 18528
rect 27956 18464 27972 18528
rect 28036 18464 28042 18528
rect 27646 18463 28042 18464
rect 0 18050 800 18080
rect 1301 18050 1367 18053
rect 0 18048 1367 18050
rect 0 17992 1306 18048
rect 1362 17992 1367 18048
rect 0 17990 1367 17992
rect 0 17960 800 17990
rect 1301 17987 1367 17990
rect 2906 17984 3302 17985
rect 2906 17920 2912 17984
rect 2976 17920 2992 17984
rect 3056 17920 3072 17984
rect 3136 17920 3152 17984
rect 3216 17920 3232 17984
rect 3296 17920 3302 17984
rect 2906 17919 3302 17920
rect 10906 17984 11302 17985
rect 10906 17920 10912 17984
rect 10976 17920 10992 17984
rect 11056 17920 11072 17984
rect 11136 17920 11152 17984
rect 11216 17920 11232 17984
rect 11296 17920 11302 17984
rect 10906 17919 11302 17920
rect 18906 17984 19302 17985
rect 18906 17920 18912 17984
rect 18976 17920 18992 17984
rect 19056 17920 19072 17984
rect 19136 17920 19152 17984
rect 19216 17920 19232 17984
rect 19296 17920 19302 17984
rect 18906 17919 19302 17920
rect 26906 17984 27302 17985
rect 26906 17920 26912 17984
rect 26976 17920 26992 17984
rect 27056 17920 27072 17984
rect 27136 17920 27152 17984
rect 27216 17920 27232 17984
rect 27296 17920 27302 17984
rect 26906 17919 27302 17920
rect 0 17506 800 17536
rect 1209 17506 1275 17509
rect 0 17504 1275 17506
rect 0 17448 1214 17504
rect 1270 17448 1275 17504
rect 0 17446 1275 17448
rect 0 17416 800 17446
rect 1209 17443 1275 17446
rect 3646 17440 4042 17441
rect 3646 17376 3652 17440
rect 3716 17376 3732 17440
rect 3796 17376 3812 17440
rect 3876 17376 3892 17440
rect 3956 17376 3972 17440
rect 4036 17376 4042 17440
rect 3646 17375 4042 17376
rect 11646 17440 12042 17441
rect 11646 17376 11652 17440
rect 11716 17376 11732 17440
rect 11796 17376 11812 17440
rect 11876 17376 11892 17440
rect 11956 17376 11972 17440
rect 12036 17376 12042 17440
rect 11646 17375 12042 17376
rect 19646 17440 20042 17441
rect 19646 17376 19652 17440
rect 19716 17376 19732 17440
rect 19796 17376 19812 17440
rect 19876 17376 19892 17440
rect 19956 17376 19972 17440
rect 20036 17376 20042 17440
rect 19646 17375 20042 17376
rect 27646 17440 28042 17441
rect 27646 17376 27652 17440
rect 27716 17376 27732 17440
rect 27796 17376 27812 17440
rect 27876 17376 27892 17440
rect 27956 17376 27972 17440
rect 28036 17376 28042 17440
rect 27646 17375 28042 17376
rect 3049 17098 3115 17101
rect 3366 17098 3372 17100
rect 3049 17096 3372 17098
rect 3049 17040 3054 17096
rect 3110 17040 3372 17096
rect 3049 17038 3372 17040
rect 3049 17035 3115 17038
rect 3366 17036 3372 17038
rect 3436 17036 3442 17100
rect 0 16962 800 16992
rect 1301 16962 1367 16965
rect 0 16960 1367 16962
rect 0 16904 1306 16960
rect 1362 16904 1367 16960
rect 0 16902 1367 16904
rect 0 16872 800 16902
rect 1301 16899 1367 16902
rect 2906 16896 3302 16897
rect 2906 16832 2912 16896
rect 2976 16832 2992 16896
rect 3056 16832 3072 16896
rect 3136 16832 3152 16896
rect 3216 16832 3232 16896
rect 3296 16832 3302 16896
rect 2906 16831 3302 16832
rect 10906 16896 11302 16897
rect 10906 16832 10912 16896
rect 10976 16832 10992 16896
rect 11056 16832 11072 16896
rect 11136 16832 11152 16896
rect 11216 16832 11232 16896
rect 11296 16832 11302 16896
rect 10906 16831 11302 16832
rect 18906 16896 19302 16897
rect 18906 16832 18912 16896
rect 18976 16832 18992 16896
rect 19056 16832 19072 16896
rect 19136 16832 19152 16896
rect 19216 16832 19232 16896
rect 19296 16832 19302 16896
rect 18906 16831 19302 16832
rect 26906 16896 27302 16897
rect 26906 16832 26912 16896
rect 26976 16832 26992 16896
rect 27056 16832 27072 16896
rect 27136 16832 27152 16896
rect 27216 16832 27232 16896
rect 27296 16832 27302 16896
rect 26906 16831 27302 16832
rect 2630 16492 2636 16556
rect 2700 16554 2706 16556
rect 5901 16554 5967 16557
rect 2700 16552 5967 16554
rect 2700 16496 5906 16552
rect 5962 16496 5967 16552
rect 2700 16494 5967 16496
rect 2700 16492 2706 16494
rect 5901 16491 5967 16494
rect 0 16418 800 16448
rect 1485 16418 1551 16421
rect 0 16416 1551 16418
rect 0 16360 1490 16416
rect 1546 16360 1551 16416
rect 0 16358 1551 16360
rect 0 16328 800 16358
rect 1485 16355 1551 16358
rect 3646 16352 4042 16353
rect 3646 16288 3652 16352
rect 3716 16288 3732 16352
rect 3796 16288 3812 16352
rect 3876 16288 3892 16352
rect 3956 16288 3972 16352
rect 4036 16288 4042 16352
rect 3646 16287 4042 16288
rect 11646 16352 12042 16353
rect 11646 16288 11652 16352
rect 11716 16288 11732 16352
rect 11796 16288 11812 16352
rect 11876 16288 11892 16352
rect 11956 16288 11972 16352
rect 12036 16288 12042 16352
rect 11646 16287 12042 16288
rect 19646 16352 20042 16353
rect 19646 16288 19652 16352
rect 19716 16288 19732 16352
rect 19796 16288 19812 16352
rect 19876 16288 19892 16352
rect 19956 16288 19972 16352
rect 20036 16288 20042 16352
rect 19646 16287 20042 16288
rect 27646 16352 28042 16353
rect 27646 16288 27652 16352
rect 27716 16288 27732 16352
rect 27796 16288 27812 16352
rect 27876 16288 27892 16352
rect 27956 16288 27972 16352
rect 28036 16288 28042 16352
rect 27646 16287 28042 16288
rect 1577 16282 1643 16285
rect 1710 16282 1716 16284
rect 1577 16280 1716 16282
rect 1577 16224 1582 16280
rect 1638 16224 1716 16280
rect 1577 16222 1716 16224
rect 1577 16219 1643 16222
rect 1710 16220 1716 16222
rect 1780 16220 1786 16284
rect 0 15874 800 15904
rect 1301 15874 1367 15877
rect 0 15872 1367 15874
rect 0 15816 1306 15872
rect 1362 15816 1367 15872
rect 0 15814 1367 15816
rect 0 15784 800 15814
rect 1301 15811 1367 15814
rect 2906 15808 3302 15809
rect 2906 15744 2912 15808
rect 2976 15744 2992 15808
rect 3056 15744 3072 15808
rect 3136 15744 3152 15808
rect 3216 15744 3232 15808
rect 3296 15744 3302 15808
rect 2906 15743 3302 15744
rect 10906 15808 11302 15809
rect 10906 15744 10912 15808
rect 10976 15744 10992 15808
rect 11056 15744 11072 15808
rect 11136 15744 11152 15808
rect 11216 15744 11232 15808
rect 11296 15744 11302 15808
rect 10906 15743 11302 15744
rect 18906 15808 19302 15809
rect 18906 15744 18912 15808
rect 18976 15744 18992 15808
rect 19056 15744 19072 15808
rect 19136 15744 19152 15808
rect 19216 15744 19232 15808
rect 19296 15744 19302 15808
rect 18906 15743 19302 15744
rect 26906 15808 27302 15809
rect 26906 15744 26912 15808
rect 26976 15744 26992 15808
rect 27056 15744 27072 15808
rect 27136 15744 27152 15808
rect 27216 15744 27232 15808
rect 27296 15744 27302 15808
rect 26906 15743 27302 15744
rect 0 15330 800 15360
rect 1393 15330 1459 15333
rect 0 15328 1459 15330
rect 0 15272 1398 15328
rect 1454 15272 1459 15328
rect 0 15270 1459 15272
rect 0 15240 800 15270
rect 1393 15267 1459 15270
rect 3646 15264 4042 15265
rect 3646 15200 3652 15264
rect 3716 15200 3732 15264
rect 3796 15200 3812 15264
rect 3876 15200 3892 15264
rect 3956 15200 3972 15264
rect 4036 15200 4042 15264
rect 3646 15199 4042 15200
rect 11646 15264 12042 15265
rect 11646 15200 11652 15264
rect 11716 15200 11732 15264
rect 11796 15200 11812 15264
rect 11876 15200 11892 15264
rect 11956 15200 11972 15264
rect 12036 15200 12042 15264
rect 11646 15199 12042 15200
rect 19646 15264 20042 15265
rect 19646 15200 19652 15264
rect 19716 15200 19732 15264
rect 19796 15200 19812 15264
rect 19876 15200 19892 15264
rect 19956 15200 19972 15264
rect 20036 15200 20042 15264
rect 19646 15199 20042 15200
rect 27646 15264 28042 15265
rect 27646 15200 27652 15264
rect 27716 15200 27732 15264
rect 27796 15200 27812 15264
rect 27876 15200 27892 15264
rect 27956 15200 27972 15264
rect 28036 15200 28042 15264
rect 27646 15199 28042 15200
rect 2630 14996 2636 15060
rect 2700 15058 2706 15060
rect 2957 15058 3023 15061
rect 2700 15056 3023 15058
rect 2700 15000 2962 15056
rect 3018 15000 3023 15056
rect 2700 14998 3023 15000
rect 2700 14996 2706 14998
rect 2957 14995 3023 14998
rect 0 14786 800 14816
rect 1301 14786 1367 14789
rect 0 14784 1367 14786
rect 0 14728 1306 14784
rect 1362 14728 1367 14784
rect 0 14726 1367 14728
rect 0 14696 800 14726
rect 1301 14723 1367 14726
rect 2906 14720 3302 14721
rect 2906 14656 2912 14720
rect 2976 14656 2992 14720
rect 3056 14656 3072 14720
rect 3136 14656 3152 14720
rect 3216 14656 3232 14720
rect 3296 14656 3302 14720
rect 2906 14655 3302 14656
rect 10906 14720 11302 14721
rect 10906 14656 10912 14720
rect 10976 14656 10992 14720
rect 11056 14656 11072 14720
rect 11136 14656 11152 14720
rect 11216 14656 11232 14720
rect 11296 14656 11302 14720
rect 10906 14655 11302 14656
rect 18906 14720 19302 14721
rect 18906 14656 18912 14720
rect 18976 14656 18992 14720
rect 19056 14656 19072 14720
rect 19136 14656 19152 14720
rect 19216 14656 19232 14720
rect 19296 14656 19302 14720
rect 18906 14655 19302 14656
rect 26906 14720 27302 14721
rect 26906 14656 26912 14720
rect 26976 14656 26992 14720
rect 27056 14656 27072 14720
rect 27136 14656 27152 14720
rect 27216 14656 27232 14720
rect 27296 14656 27302 14720
rect 26906 14655 27302 14656
rect 0 14242 800 14272
rect 1301 14242 1367 14245
rect 0 14240 1367 14242
rect 0 14184 1306 14240
rect 1362 14184 1367 14240
rect 0 14182 1367 14184
rect 0 14152 800 14182
rect 1301 14179 1367 14182
rect 3646 14176 4042 14177
rect 3646 14112 3652 14176
rect 3716 14112 3732 14176
rect 3796 14112 3812 14176
rect 3876 14112 3892 14176
rect 3956 14112 3972 14176
rect 4036 14112 4042 14176
rect 3646 14111 4042 14112
rect 11646 14176 12042 14177
rect 11646 14112 11652 14176
rect 11716 14112 11732 14176
rect 11796 14112 11812 14176
rect 11876 14112 11892 14176
rect 11956 14112 11972 14176
rect 12036 14112 12042 14176
rect 11646 14111 12042 14112
rect 19646 14176 20042 14177
rect 19646 14112 19652 14176
rect 19716 14112 19732 14176
rect 19796 14112 19812 14176
rect 19876 14112 19892 14176
rect 19956 14112 19972 14176
rect 20036 14112 20042 14176
rect 19646 14111 20042 14112
rect 27646 14176 28042 14177
rect 27646 14112 27652 14176
rect 27716 14112 27732 14176
rect 27796 14112 27812 14176
rect 27876 14112 27892 14176
rect 27956 14112 27972 14176
rect 28036 14112 28042 14176
rect 27646 14111 28042 14112
rect 2957 13970 3023 13973
rect 3509 13970 3575 13973
rect 3877 13970 3943 13973
rect 2957 13968 3943 13970
rect 2957 13912 2962 13968
rect 3018 13912 3514 13968
rect 3570 13912 3882 13968
rect 3938 13912 3943 13968
rect 2957 13910 3943 13912
rect 2957 13907 3023 13910
rect 3509 13907 3575 13910
rect 3877 13907 3943 13910
rect 0 13698 800 13728
rect 1301 13698 1367 13701
rect 0 13696 1367 13698
rect 0 13640 1306 13696
rect 1362 13640 1367 13696
rect 0 13638 1367 13640
rect 0 13608 800 13638
rect 1301 13635 1367 13638
rect 2906 13632 3302 13633
rect 2906 13568 2912 13632
rect 2976 13568 2992 13632
rect 3056 13568 3072 13632
rect 3136 13568 3152 13632
rect 3216 13568 3232 13632
rect 3296 13568 3302 13632
rect 2906 13567 3302 13568
rect 10906 13632 11302 13633
rect 10906 13568 10912 13632
rect 10976 13568 10992 13632
rect 11056 13568 11072 13632
rect 11136 13568 11152 13632
rect 11216 13568 11232 13632
rect 11296 13568 11302 13632
rect 10906 13567 11302 13568
rect 18906 13632 19302 13633
rect 18906 13568 18912 13632
rect 18976 13568 18992 13632
rect 19056 13568 19072 13632
rect 19136 13568 19152 13632
rect 19216 13568 19232 13632
rect 19296 13568 19302 13632
rect 18906 13567 19302 13568
rect 26906 13632 27302 13633
rect 26906 13568 26912 13632
rect 26976 13568 26992 13632
rect 27056 13568 27072 13632
rect 27136 13568 27152 13632
rect 27216 13568 27232 13632
rect 27296 13568 27302 13632
rect 26906 13567 27302 13568
rect 0 13154 800 13184
rect 1209 13154 1275 13157
rect 0 13152 1275 13154
rect 0 13096 1214 13152
rect 1270 13096 1275 13152
rect 0 13094 1275 13096
rect 0 13064 800 13094
rect 1209 13091 1275 13094
rect 3646 13088 4042 13089
rect 3646 13024 3652 13088
rect 3716 13024 3732 13088
rect 3796 13024 3812 13088
rect 3876 13024 3892 13088
rect 3956 13024 3972 13088
rect 4036 13024 4042 13088
rect 3646 13023 4042 13024
rect 11646 13088 12042 13089
rect 11646 13024 11652 13088
rect 11716 13024 11732 13088
rect 11796 13024 11812 13088
rect 11876 13024 11892 13088
rect 11956 13024 11972 13088
rect 12036 13024 12042 13088
rect 11646 13023 12042 13024
rect 19646 13088 20042 13089
rect 19646 13024 19652 13088
rect 19716 13024 19732 13088
rect 19796 13024 19812 13088
rect 19876 13024 19892 13088
rect 19956 13024 19972 13088
rect 20036 13024 20042 13088
rect 19646 13023 20042 13024
rect 27646 13088 28042 13089
rect 27646 13024 27652 13088
rect 27716 13024 27732 13088
rect 27796 13024 27812 13088
rect 27876 13024 27892 13088
rect 27956 13024 27972 13088
rect 28036 13024 28042 13088
rect 27646 13023 28042 13024
rect 0 12610 800 12640
rect 1301 12610 1367 12613
rect 0 12608 1367 12610
rect 0 12552 1306 12608
rect 1362 12552 1367 12608
rect 0 12550 1367 12552
rect 0 12520 800 12550
rect 1301 12547 1367 12550
rect 2906 12544 3302 12545
rect 2906 12480 2912 12544
rect 2976 12480 2992 12544
rect 3056 12480 3072 12544
rect 3136 12480 3152 12544
rect 3216 12480 3232 12544
rect 3296 12480 3302 12544
rect 2906 12479 3302 12480
rect 10906 12544 11302 12545
rect 10906 12480 10912 12544
rect 10976 12480 10992 12544
rect 11056 12480 11072 12544
rect 11136 12480 11152 12544
rect 11216 12480 11232 12544
rect 11296 12480 11302 12544
rect 10906 12479 11302 12480
rect 18906 12544 19302 12545
rect 18906 12480 18912 12544
rect 18976 12480 18992 12544
rect 19056 12480 19072 12544
rect 19136 12480 19152 12544
rect 19216 12480 19232 12544
rect 19296 12480 19302 12544
rect 18906 12479 19302 12480
rect 26906 12544 27302 12545
rect 26906 12480 26912 12544
rect 26976 12480 26992 12544
rect 27056 12480 27072 12544
rect 27136 12480 27152 12544
rect 27216 12480 27232 12544
rect 27296 12480 27302 12544
rect 26906 12479 27302 12480
rect 0 12066 800 12096
rect 1301 12066 1367 12069
rect 0 12064 1367 12066
rect 0 12008 1306 12064
rect 1362 12008 1367 12064
rect 0 12006 1367 12008
rect 0 11976 800 12006
rect 1301 12003 1367 12006
rect 1945 12066 2011 12069
rect 2078 12066 2084 12068
rect 1945 12064 2084 12066
rect 1945 12008 1950 12064
rect 2006 12008 2084 12064
rect 1945 12006 2084 12008
rect 1945 12003 2011 12006
rect 2078 12004 2084 12006
rect 2148 12004 2154 12068
rect 3646 12000 4042 12001
rect 3646 11936 3652 12000
rect 3716 11936 3732 12000
rect 3796 11936 3812 12000
rect 3876 11936 3892 12000
rect 3956 11936 3972 12000
rect 4036 11936 4042 12000
rect 3646 11935 4042 11936
rect 11646 12000 12042 12001
rect 11646 11936 11652 12000
rect 11716 11936 11732 12000
rect 11796 11936 11812 12000
rect 11876 11936 11892 12000
rect 11956 11936 11972 12000
rect 12036 11936 12042 12000
rect 11646 11935 12042 11936
rect 19646 12000 20042 12001
rect 19646 11936 19652 12000
rect 19716 11936 19732 12000
rect 19796 11936 19812 12000
rect 19876 11936 19892 12000
rect 19956 11936 19972 12000
rect 20036 11936 20042 12000
rect 19646 11935 20042 11936
rect 27646 12000 28042 12001
rect 27646 11936 27652 12000
rect 27716 11936 27732 12000
rect 27796 11936 27812 12000
rect 27876 11936 27892 12000
rect 27956 11936 27972 12000
rect 28036 11936 28042 12000
rect 27646 11935 28042 11936
rect 0 11522 800 11552
rect 1301 11522 1367 11525
rect 0 11520 1367 11522
rect 0 11464 1306 11520
rect 1362 11464 1367 11520
rect 0 11462 1367 11464
rect 0 11432 800 11462
rect 1301 11459 1367 11462
rect 2906 11456 3302 11457
rect 2906 11392 2912 11456
rect 2976 11392 2992 11456
rect 3056 11392 3072 11456
rect 3136 11392 3152 11456
rect 3216 11392 3232 11456
rect 3296 11392 3302 11456
rect 2906 11391 3302 11392
rect 10906 11456 11302 11457
rect 10906 11392 10912 11456
rect 10976 11392 10992 11456
rect 11056 11392 11072 11456
rect 11136 11392 11152 11456
rect 11216 11392 11232 11456
rect 11296 11392 11302 11456
rect 10906 11391 11302 11392
rect 18906 11456 19302 11457
rect 18906 11392 18912 11456
rect 18976 11392 18992 11456
rect 19056 11392 19072 11456
rect 19136 11392 19152 11456
rect 19216 11392 19232 11456
rect 19296 11392 19302 11456
rect 18906 11391 19302 11392
rect 26906 11456 27302 11457
rect 26906 11392 26912 11456
rect 26976 11392 26992 11456
rect 27056 11392 27072 11456
rect 27136 11392 27152 11456
rect 27216 11392 27232 11456
rect 27296 11392 27302 11456
rect 26906 11391 27302 11392
rect 3366 11324 3372 11388
rect 3436 11386 3442 11388
rect 3785 11386 3851 11389
rect 3436 11384 3851 11386
rect 3436 11328 3790 11384
rect 3846 11328 3851 11384
rect 3436 11326 3851 11328
rect 3436 11324 3442 11326
rect 3785 11323 3851 11326
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 3646 10912 4042 10913
rect 3646 10848 3652 10912
rect 3716 10848 3732 10912
rect 3796 10848 3812 10912
rect 3876 10848 3892 10912
rect 3956 10848 3972 10912
rect 4036 10848 4042 10912
rect 3646 10847 4042 10848
rect 11646 10912 12042 10913
rect 11646 10848 11652 10912
rect 11716 10848 11732 10912
rect 11796 10848 11812 10912
rect 11876 10848 11892 10912
rect 11956 10848 11972 10912
rect 12036 10848 12042 10912
rect 11646 10847 12042 10848
rect 19646 10912 20042 10913
rect 19646 10848 19652 10912
rect 19716 10848 19732 10912
rect 19796 10848 19812 10912
rect 19876 10848 19892 10912
rect 19956 10848 19972 10912
rect 20036 10848 20042 10912
rect 19646 10847 20042 10848
rect 27646 10912 28042 10913
rect 27646 10848 27652 10912
rect 27716 10848 27732 10912
rect 27796 10848 27812 10912
rect 27876 10848 27892 10912
rect 27956 10848 27972 10912
rect 28036 10848 28042 10912
rect 27646 10847 28042 10848
rect 0 10434 800 10464
rect 1301 10434 1367 10437
rect 0 10432 1367 10434
rect 0 10376 1306 10432
rect 1362 10376 1367 10432
rect 0 10374 1367 10376
rect 0 10344 800 10374
rect 1301 10371 1367 10374
rect 2906 10368 3302 10369
rect 2906 10304 2912 10368
rect 2976 10304 2992 10368
rect 3056 10304 3072 10368
rect 3136 10304 3152 10368
rect 3216 10304 3232 10368
rect 3296 10304 3302 10368
rect 2906 10303 3302 10304
rect 10906 10368 11302 10369
rect 10906 10304 10912 10368
rect 10976 10304 10992 10368
rect 11056 10304 11072 10368
rect 11136 10304 11152 10368
rect 11216 10304 11232 10368
rect 11296 10304 11302 10368
rect 10906 10303 11302 10304
rect 18906 10368 19302 10369
rect 18906 10304 18912 10368
rect 18976 10304 18992 10368
rect 19056 10304 19072 10368
rect 19136 10304 19152 10368
rect 19216 10304 19232 10368
rect 19296 10304 19302 10368
rect 18906 10303 19302 10304
rect 26906 10368 27302 10369
rect 26906 10304 26912 10368
rect 26976 10304 26992 10368
rect 27056 10304 27072 10368
rect 27136 10304 27152 10368
rect 27216 10304 27232 10368
rect 27296 10304 27302 10368
rect 26906 10303 27302 10304
rect 0 9890 800 9920
rect 1301 9890 1367 9893
rect 0 9888 1367 9890
rect 0 9832 1306 9888
rect 1362 9832 1367 9888
rect 0 9830 1367 9832
rect 0 9800 800 9830
rect 1301 9827 1367 9830
rect 3646 9824 4042 9825
rect 3646 9760 3652 9824
rect 3716 9760 3732 9824
rect 3796 9760 3812 9824
rect 3876 9760 3892 9824
rect 3956 9760 3972 9824
rect 4036 9760 4042 9824
rect 3646 9759 4042 9760
rect 11646 9824 12042 9825
rect 11646 9760 11652 9824
rect 11716 9760 11732 9824
rect 11796 9760 11812 9824
rect 11876 9760 11892 9824
rect 11956 9760 11972 9824
rect 12036 9760 12042 9824
rect 11646 9759 12042 9760
rect 19646 9824 20042 9825
rect 19646 9760 19652 9824
rect 19716 9760 19732 9824
rect 19796 9760 19812 9824
rect 19876 9760 19892 9824
rect 19956 9760 19972 9824
rect 20036 9760 20042 9824
rect 19646 9759 20042 9760
rect 27646 9824 28042 9825
rect 27646 9760 27652 9824
rect 27716 9760 27732 9824
rect 27796 9760 27812 9824
rect 27876 9760 27892 9824
rect 27956 9760 27972 9824
rect 28036 9760 28042 9824
rect 27646 9759 28042 9760
rect 0 9346 800 9376
rect 1301 9346 1367 9349
rect 0 9344 1367 9346
rect 0 9288 1306 9344
rect 1362 9288 1367 9344
rect 0 9286 1367 9288
rect 0 9256 800 9286
rect 1301 9283 1367 9286
rect 2906 9280 3302 9281
rect 2906 9216 2912 9280
rect 2976 9216 2992 9280
rect 3056 9216 3072 9280
rect 3136 9216 3152 9280
rect 3216 9216 3232 9280
rect 3296 9216 3302 9280
rect 2906 9215 3302 9216
rect 10906 9280 11302 9281
rect 10906 9216 10912 9280
rect 10976 9216 10992 9280
rect 11056 9216 11072 9280
rect 11136 9216 11152 9280
rect 11216 9216 11232 9280
rect 11296 9216 11302 9280
rect 10906 9215 11302 9216
rect 18906 9280 19302 9281
rect 18906 9216 18912 9280
rect 18976 9216 18992 9280
rect 19056 9216 19072 9280
rect 19136 9216 19152 9280
rect 19216 9216 19232 9280
rect 19296 9216 19302 9280
rect 18906 9215 19302 9216
rect 26906 9280 27302 9281
rect 26906 9216 26912 9280
rect 26976 9216 26992 9280
rect 27056 9216 27072 9280
rect 27136 9216 27152 9280
rect 27216 9216 27232 9280
rect 27296 9216 27302 9280
rect 26906 9215 27302 9216
rect 0 8802 800 8832
rect 1301 8802 1367 8805
rect 0 8800 1367 8802
rect 0 8744 1306 8800
rect 1362 8744 1367 8800
rect 0 8742 1367 8744
rect 0 8712 800 8742
rect 1301 8739 1367 8742
rect 3646 8736 4042 8737
rect 3646 8672 3652 8736
rect 3716 8672 3732 8736
rect 3796 8672 3812 8736
rect 3876 8672 3892 8736
rect 3956 8672 3972 8736
rect 4036 8672 4042 8736
rect 3646 8671 4042 8672
rect 11646 8736 12042 8737
rect 11646 8672 11652 8736
rect 11716 8672 11732 8736
rect 11796 8672 11812 8736
rect 11876 8672 11892 8736
rect 11956 8672 11972 8736
rect 12036 8672 12042 8736
rect 11646 8671 12042 8672
rect 19646 8736 20042 8737
rect 19646 8672 19652 8736
rect 19716 8672 19732 8736
rect 19796 8672 19812 8736
rect 19876 8672 19892 8736
rect 19956 8672 19972 8736
rect 20036 8672 20042 8736
rect 19646 8671 20042 8672
rect 27646 8736 28042 8737
rect 27646 8672 27652 8736
rect 27716 8672 27732 8736
rect 27796 8672 27812 8736
rect 27876 8672 27892 8736
rect 27956 8672 27972 8736
rect 28036 8672 28042 8736
rect 27646 8671 28042 8672
rect 0 8258 800 8288
rect 1301 8258 1367 8261
rect 0 8256 1367 8258
rect 0 8200 1306 8256
rect 1362 8200 1367 8256
rect 0 8198 1367 8200
rect 0 8168 800 8198
rect 1301 8195 1367 8198
rect 2906 8192 3302 8193
rect 2906 8128 2912 8192
rect 2976 8128 2992 8192
rect 3056 8128 3072 8192
rect 3136 8128 3152 8192
rect 3216 8128 3232 8192
rect 3296 8128 3302 8192
rect 2906 8127 3302 8128
rect 10906 8192 11302 8193
rect 10906 8128 10912 8192
rect 10976 8128 10992 8192
rect 11056 8128 11072 8192
rect 11136 8128 11152 8192
rect 11216 8128 11232 8192
rect 11296 8128 11302 8192
rect 10906 8127 11302 8128
rect 18906 8192 19302 8193
rect 18906 8128 18912 8192
rect 18976 8128 18992 8192
rect 19056 8128 19072 8192
rect 19136 8128 19152 8192
rect 19216 8128 19232 8192
rect 19296 8128 19302 8192
rect 18906 8127 19302 8128
rect 26906 8192 27302 8193
rect 26906 8128 26912 8192
rect 26976 8128 26992 8192
rect 27056 8128 27072 8192
rect 27136 8128 27152 8192
rect 27216 8128 27232 8192
rect 27296 8128 27302 8192
rect 26906 8127 27302 8128
rect 0 7714 800 7744
rect 1209 7714 1275 7717
rect 0 7712 1275 7714
rect 0 7656 1214 7712
rect 1270 7656 1275 7712
rect 0 7654 1275 7656
rect 0 7624 800 7654
rect 1209 7651 1275 7654
rect 3646 7648 4042 7649
rect 3646 7584 3652 7648
rect 3716 7584 3732 7648
rect 3796 7584 3812 7648
rect 3876 7584 3892 7648
rect 3956 7584 3972 7648
rect 4036 7584 4042 7648
rect 3646 7583 4042 7584
rect 11646 7648 12042 7649
rect 11646 7584 11652 7648
rect 11716 7584 11732 7648
rect 11796 7584 11812 7648
rect 11876 7584 11892 7648
rect 11956 7584 11972 7648
rect 12036 7584 12042 7648
rect 11646 7583 12042 7584
rect 19646 7648 20042 7649
rect 19646 7584 19652 7648
rect 19716 7584 19732 7648
rect 19796 7584 19812 7648
rect 19876 7584 19892 7648
rect 19956 7584 19972 7648
rect 20036 7584 20042 7648
rect 19646 7583 20042 7584
rect 27646 7648 28042 7649
rect 27646 7584 27652 7648
rect 27716 7584 27732 7648
rect 27796 7584 27812 7648
rect 27876 7584 27892 7648
rect 27956 7584 27972 7648
rect 28036 7584 28042 7648
rect 27646 7583 28042 7584
rect 28349 7442 28415 7445
rect 29200 7442 30000 7472
rect 28349 7440 30000 7442
rect 28349 7384 28354 7440
rect 28410 7384 30000 7440
rect 28349 7382 30000 7384
rect 28349 7379 28415 7382
rect 29200 7352 30000 7382
rect 0 7170 800 7200
rect 1209 7170 1275 7173
rect 0 7168 1275 7170
rect 0 7112 1214 7168
rect 1270 7112 1275 7168
rect 0 7110 1275 7112
rect 0 7080 800 7110
rect 1209 7107 1275 7110
rect 2906 7104 3302 7105
rect 2906 7040 2912 7104
rect 2976 7040 2992 7104
rect 3056 7040 3072 7104
rect 3136 7040 3152 7104
rect 3216 7040 3232 7104
rect 3296 7040 3302 7104
rect 2906 7039 3302 7040
rect 10906 7104 11302 7105
rect 10906 7040 10912 7104
rect 10976 7040 10992 7104
rect 11056 7040 11072 7104
rect 11136 7040 11152 7104
rect 11216 7040 11232 7104
rect 11296 7040 11302 7104
rect 10906 7039 11302 7040
rect 18906 7104 19302 7105
rect 18906 7040 18912 7104
rect 18976 7040 18992 7104
rect 19056 7040 19072 7104
rect 19136 7040 19152 7104
rect 19216 7040 19232 7104
rect 19296 7040 19302 7104
rect 18906 7039 19302 7040
rect 26906 7104 27302 7105
rect 26906 7040 26912 7104
rect 26976 7040 26992 7104
rect 27056 7040 27072 7104
rect 27136 7040 27152 7104
rect 27216 7040 27232 7104
rect 27296 7040 27302 7104
rect 26906 7039 27302 7040
rect 0 6626 800 6656
rect 1301 6626 1367 6629
rect 0 6624 1367 6626
rect 0 6568 1306 6624
rect 1362 6568 1367 6624
rect 0 6566 1367 6568
rect 0 6536 800 6566
rect 1301 6563 1367 6566
rect 3646 6560 4042 6561
rect 3646 6496 3652 6560
rect 3716 6496 3732 6560
rect 3796 6496 3812 6560
rect 3876 6496 3892 6560
rect 3956 6496 3972 6560
rect 4036 6496 4042 6560
rect 3646 6495 4042 6496
rect 11646 6560 12042 6561
rect 11646 6496 11652 6560
rect 11716 6496 11732 6560
rect 11796 6496 11812 6560
rect 11876 6496 11892 6560
rect 11956 6496 11972 6560
rect 12036 6496 12042 6560
rect 11646 6495 12042 6496
rect 19646 6560 20042 6561
rect 19646 6496 19652 6560
rect 19716 6496 19732 6560
rect 19796 6496 19812 6560
rect 19876 6496 19892 6560
rect 19956 6496 19972 6560
rect 20036 6496 20042 6560
rect 19646 6495 20042 6496
rect 27646 6560 28042 6561
rect 27646 6496 27652 6560
rect 27716 6496 27732 6560
rect 27796 6496 27812 6560
rect 27876 6496 27892 6560
rect 27956 6496 27972 6560
rect 28036 6496 28042 6560
rect 27646 6495 28042 6496
rect 6177 6218 6243 6221
rect 14273 6218 14339 6221
rect 6177 6216 14339 6218
rect 6177 6160 6182 6216
rect 6238 6160 14278 6216
rect 14334 6160 14339 6216
rect 6177 6158 14339 6160
rect 6177 6155 6243 6158
rect 14273 6155 14339 6158
rect 0 6082 800 6112
rect 1301 6082 1367 6085
rect 0 6080 1367 6082
rect 0 6024 1306 6080
rect 1362 6024 1367 6080
rect 0 6022 1367 6024
rect 0 5992 800 6022
rect 1301 6019 1367 6022
rect 2906 6016 3302 6017
rect 2906 5952 2912 6016
rect 2976 5952 2992 6016
rect 3056 5952 3072 6016
rect 3136 5952 3152 6016
rect 3216 5952 3232 6016
rect 3296 5952 3302 6016
rect 2906 5951 3302 5952
rect 10906 6016 11302 6017
rect 10906 5952 10912 6016
rect 10976 5952 10992 6016
rect 11056 5952 11072 6016
rect 11136 5952 11152 6016
rect 11216 5952 11232 6016
rect 11296 5952 11302 6016
rect 10906 5951 11302 5952
rect 18906 6016 19302 6017
rect 18906 5952 18912 6016
rect 18976 5952 18992 6016
rect 19056 5952 19072 6016
rect 19136 5952 19152 6016
rect 19216 5952 19232 6016
rect 19296 5952 19302 6016
rect 18906 5951 19302 5952
rect 26906 6016 27302 6017
rect 26906 5952 26912 6016
rect 26976 5952 26992 6016
rect 27056 5952 27072 6016
rect 27136 5952 27152 6016
rect 27216 5952 27232 6016
rect 27296 5952 27302 6016
rect 26906 5951 27302 5952
rect 0 5538 800 5568
rect 1301 5538 1367 5541
rect 0 5536 1367 5538
rect 0 5480 1306 5536
rect 1362 5480 1367 5536
rect 0 5478 1367 5480
rect 0 5448 800 5478
rect 1301 5475 1367 5478
rect 3646 5472 4042 5473
rect 3646 5408 3652 5472
rect 3716 5408 3732 5472
rect 3796 5408 3812 5472
rect 3876 5408 3892 5472
rect 3956 5408 3972 5472
rect 4036 5408 4042 5472
rect 3646 5407 4042 5408
rect 11646 5472 12042 5473
rect 11646 5408 11652 5472
rect 11716 5408 11732 5472
rect 11796 5408 11812 5472
rect 11876 5408 11892 5472
rect 11956 5408 11972 5472
rect 12036 5408 12042 5472
rect 11646 5407 12042 5408
rect 19646 5472 20042 5473
rect 19646 5408 19652 5472
rect 19716 5408 19732 5472
rect 19796 5408 19812 5472
rect 19876 5408 19892 5472
rect 19956 5408 19972 5472
rect 20036 5408 20042 5472
rect 19646 5407 20042 5408
rect 27646 5472 28042 5473
rect 27646 5408 27652 5472
rect 27716 5408 27732 5472
rect 27796 5408 27812 5472
rect 27876 5408 27892 5472
rect 27956 5408 27972 5472
rect 28036 5408 28042 5472
rect 27646 5407 28042 5408
rect 0 4994 800 5024
rect 1301 4994 1367 4997
rect 0 4992 1367 4994
rect 0 4936 1306 4992
rect 1362 4936 1367 4992
rect 0 4934 1367 4936
rect 0 4904 800 4934
rect 1301 4931 1367 4934
rect 2906 4928 3302 4929
rect 2906 4864 2912 4928
rect 2976 4864 2992 4928
rect 3056 4864 3072 4928
rect 3136 4864 3152 4928
rect 3216 4864 3232 4928
rect 3296 4864 3302 4928
rect 2906 4863 3302 4864
rect 10906 4928 11302 4929
rect 10906 4864 10912 4928
rect 10976 4864 10992 4928
rect 11056 4864 11072 4928
rect 11136 4864 11152 4928
rect 11216 4864 11232 4928
rect 11296 4864 11302 4928
rect 10906 4863 11302 4864
rect 18906 4928 19302 4929
rect 18906 4864 18912 4928
rect 18976 4864 18992 4928
rect 19056 4864 19072 4928
rect 19136 4864 19152 4928
rect 19216 4864 19232 4928
rect 19296 4864 19302 4928
rect 18906 4863 19302 4864
rect 26906 4928 27302 4929
rect 26906 4864 26912 4928
rect 26976 4864 26992 4928
rect 27056 4864 27072 4928
rect 27136 4864 27152 4928
rect 27216 4864 27232 4928
rect 27296 4864 27302 4928
rect 26906 4863 27302 4864
rect 0 4450 800 4480
rect 1025 4450 1091 4453
rect 0 4448 1091 4450
rect 0 4392 1030 4448
rect 1086 4392 1091 4448
rect 0 4390 1091 4392
rect 0 4360 800 4390
rect 1025 4387 1091 4390
rect 3646 4384 4042 4385
rect 3646 4320 3652 4384
rect 3716 4320 3732 4384
rect 3796 4320 3812 4384
rect 3876 4320 3892 4384
rect 3956 4320 3972 4384
rect 4036 4320 4042 4384
rect 3646 4319 4042 4320
rect 11646 4384 12042 4385
rect 11646 4320 11652 4384
rect 11716 4320 11732 4384
rect 11796 4320 11812 4384
rect 11876 4320 11892 4384
rect 11956 4320 11972 4384
rect 12036 4320 12042 4384
rect 11646 4319 12042 4320
rect 19646 4384 20042 4385
rect 19646 4320 19652 4384
rect 19716 4320 19732 4384
rect 19796 4320 19812 4384
rect 19876 4320 19892 4384
rect 19956 4320 19972 4384
rect 20036 4320 20042 4384
rect 19646 4319 20042 4320
rect 27646 4384 28042 4385
rect 27646 4320 27652 4384
rect 27716 4320 27732 4384
rect 27796 4320 27812 4384
rect 27876 4320 27892 4384
rect 27956 4320 27972 4384
rect 28036 4320 28042 4384
rect 27646 4319 28042 4320
rect 2906 3840 3302 3841
rect 2906 3776 2912 3840
rect 2976 3776 2992 3840
rect 3056 3776 3072 3840
rect 3136 3776 3152 3840
rect 3216 3776 3232 3840
rect 3296 3776 3302 3840
rect 2906 3775 3302 3776
rect 10906 3840 11302 3841
rect 10906 3776 10912 3840
rect 10976 3776 10992 3840
rect 11056 3776 11072 3840
rect 11136 3776 11152 3840
rect 11216 3776 11232 3840
rect 11296 3776 11302 3840
rect 10906 3775 11302 3776
rect 18906 3840 19302 3841
rect 18906 3776 18912 3840
rect 18976 3776 18992 3840
rect 19056 3776 19072 3840
rect 19136 3776 19152 3840
rect 19216 3776 19232 3840
rect 19296 3776 19302 3840
rect 18906 3775 19302 3776
rect 26906 3840 27302 3841
rect 26906 3776 26912 3840
rect 26976 3776 26992 3840
rect 27056 3776 27072 3840
rect 27136 3776 27152 3840
rect 27216 3776 27232 3840
rect 27296 3776 27302 3840
rect 26906 3775 27302 3776
rect 3646 3296 4042 3297
rect 3646 3232 3652 3296
rect 3716 3232 3732 3296
rect 3796 3232 3812 3296
rect 3876 3232 3892 3296
rect 3956 3232 3972 3296
rect 4036 3232 4042 3296
rect 3646 3231 4042 3232
rect 11646 3296 12042 3297
rect 11646 3232 11652 3296
rect 11716 3232 11732 3296
rect 11796 3232 11812 3296
rect 11876 3232 11892 3296
rect 11956 3232 11972 3296
rect 12036 3232 12042 3296
rect 11646 3231 12042 3232
rect 19646 3296 20042 3297
rect 19646 3232 19652 3296
rect 19716 3232 19732 3296
rect 19796 3232 19812 3296
rect 19876 3232 19892 3296
rect 19956 3232 19972 3296
rect 20036 3232 20042 3296
rect 19646 3231 20042 3232
rect 27646 3296 28042 3297
rect 27646 3232 27652 3296
rect 27716 3232 27732 3296
rect 27796 3232 27812 3296
rect 27876 3232 27892 3296
rect 27956 3232 27972 3296
rect 28036 3232 28042 3296
rect 27646 3231 28042 3232
rect 2906 2752 3302 2753
rect 2906 2688 2912 2752
rect 2976 2688 2992 2752
rect 3056 2688 3072 2752
rect 3136 2688 3152 2752
rect 3216 2688 3232 2752
rect 3296 2688 3302 2752
rect 2906 2687 3302 2688
rect 10906 2752 11302 2753
rect 10906 2688 10912 2752
rect 10976 2688 10992 2752
rect 11056 2688 11072 2752
rect 11136 2688 11152 2752
rect 11216 2688 11232 2752
rect 11296 2688 11302 2752
rect 10906 2687 11302 2688
rect 18906 2752 19302 2753
rect 18906 2688 18912 2752
rect 18976 2688 18992 2752
rect 19056 2688 19072 2752
rect 19136 2688 19152 2752
rect 19216 2688 19232 2752
rect 19296 2688 19302 2752
rect 18906 2687 19302 2688
rect 26906 2752 27302 2753
rect 26906 2688 26912 2752
rect 26976 2688 26992 2752
rect 27056 2688 27072 2752
rect 27136 2688 27152 2752
rect 27216 2688 27232 2752
rect 27296 2688 27302 2752
rect 26906 2687 27302 2688
rect 3646 2208 4042 2209
rect 3646 2144 3652 2208
rect 3716 2144 3732 2208
rect 3796 2144 3812 2208
rect 3876 2144 3892 2208
rect 3956 2144 3972 2208
rect 4036 2144 4042 2208
rect 3646 2143 4042 2144
rect 11646 2208 12042 2209
rect 11646 2144 11652 2208
rect 11716 2144 11732 2208
rect 11796 2144 11812 2208
rect 11876 2144 11892 2208
rect 11956 2144 11972 2208
rect 12036 2144 12042 2208
rect 11646 2143 12042 2144
rect 19646 2208 20042 2209
rect 19646 2144 19652 2208
rect 19716 2144 19732 2208
rect 19796 2144 19812 2208
rect 19876 2144 19892 2208
rect 19956 2144 19972 2208
rect 20036 2144 20042 2208
rect 19646 2143 20042 2144
rect 27646 2208 28042 2209
rect 27646 2144 27652 2208
rect 27716 2144 27732 2208
rect 27796 2144 27812 2208
rect 27876 2144 27892 2208
rect 27956 2144 27972 2208
rect 28036 2144 28042 2208
rect 27646 2143 28042 2144
<< via3 >>
rect 2912 27772 2976 27776
rect 2912 27716 2916 27772
rect 2916 27716 2972 27772
rect 2972 27716 2976 27772
rect 2912 27712 2976 27716
rect 2992 27772 3056 27776
rect 2992 27716 2996 27772
rect 2996 27716 3052 27772
rect 3052 27716 3056 27772
rect 2992 27712 3056 27716
rect 3072 27772 3136 27776
rect 3072 27716 3076 27772
rect 3076 27716 3132 27772
rect 3132 27716 3136 27772
rect 3072 27712 3136 27716
rect 3152 27772 3216 27776
rect 3152 27716 3156 27772
rect 3156 27716 3212 27772
rect 3212 27716 3216 27772
rect 3152 27712 3216 27716
rect 3232 27772 3296 27776
rect 3232 27716 3236 27772
rect 3236 27716 3292 27772
rect 3292 27716 3296 27772
rect 3232 27712 3296 27716
rect 10912 27772 10976 27776
rect 10912 27716 10916 27772
rect 10916 27716 10972 27772
rect 10972 27716 10976 27772
rect 10912 27712 10976 27716
rect 10992 27772 11056 27776
rect 10992 27716 10996 27772
rect 10996 27716 11052 27772
rect 11052 27716 11056 27772
rect 10992 27712 11056 27716
rect 11072 27772 11136 27776
rect 11072 27716 11076 27772
rect 11076 27716 11132 27772
rect 11132 27716 11136 27772
rect 11072 27712 11136 27716
rect 11152 27772 11216 27776
rect 11152 27716 11156 27772
rect 11156 27716 11212 27772
rect 11212 27716 11216 27772
rect 11152 27712 11216 27716
rect 11232 27772 11296 27776
rect 11232 27716 11236 27772
rect 11236 27716 11292 27772
rect 11292 27716 11296 27772
rect 11232 27712 11296 27716
rect 18912 27772 18976 27776
rect 18912 27716 18916 27772
rect 18916 27716 18972 27772
rect 18972 27716 18976 27772
rect 18912 27712 18976 27716
rect 18992 27772 19056 27776
rect 18992 27716 18996 27772
rect 18996 27716 19052 27772
rect 19052 27716 19056 27772
rect 18992 27712 19056 27716
rect 19072 27772 19136 27776
rect 19072 27716 19076 27772
rect 19076 27716 19132 27772
rect 19132 27716 19136 27772
rect 19072 27712 19136 27716
rect 19152 27772 19216 27776
rect 19152 27716 19156 27772
rect 19156 27716 19212 27772
rect 19212 27716 19216 27772
rect 19152 27712 19216 27716
rect 19232 27772 19296 27776
rect 19232 27716 19236 27772
rect 19236 27716 19292 27772
rect 19292 27716 19296 27772
rect 19232 27712 19296 27716
rect 26912 27772 26976 27776
rect 26912 27716 26916 27772
rect 26916 27716 26972 27772
rect 26972 27716 26976 27772
rect 26912 27712 26976 27716
rect 26992 27772 27056 27776
rect 26992 27716 26996 27772
rect 26996 27716 27052 27772
rect 27052 27716 27056 27772
rect 26992 27712 27056 27716
rect 27072 27772 27136 27776
rect 27072 27716 27076 27772
rect 27076 27716 27132 27772
rect 27132 27716 27136 27772
rect 27072 27712 27136 27716
rect 27152 27772 27216 27776
rect 27152 27716 27156 27772
rect 27156 27716 27212 27772
rect 27212 27716 27216 27772
rect 27152 27712 27216 27716
rect 27232 27772 27296 27776
rect 27232 27716 27236 27772
rect 27236 27716 27292 27772
rect 27292 27716 27296 27772
rect 27232 27712 27296 27716
rect 3652 27228 3716 27232
rect 3652 27172 3656 27228
rect 3656 27172 3712 27228
rect 3712 27172 3716 27228
rect 3652 27168 3716 27172
rect 3732 27228 3796 27232
rect 3732 27172 3736 27228
rect 3736 27172 3792 27228
rect 3792 27172 3796 27228
rect 3732 27168 3796 27172
rect 3812 27228 3876 27232
rect 3812 27172 3816 27228
rect 3816 27172 3872 27228
rect 3872 27172 3876 27228
rect 3812 27168 3876 27172
rect 3892 27228 3956 27232
rect 3892 27172 3896 27228
rect 3896 27172 3952 27228
rect 3952 27172 3956 27228
rect 3892 27168 3956 27172
rect 3972 27228 4036 27232
rect 3972 27172 3976 27228
rect 3976 27172 4032 27228
rect 4032 27172 4036 27228
rect 3972 27168 4036 27172
rect 11652 27228 11716 27232
rect 11652 27172 11656 27228
rect 11656 27172 11712 27228
rect 11712 27172 11716 27228
rect 11652 27168 11716 27172
rect 11732 27228 11796 27232
rect 11732 27172 11736 27228
rect 11736 27172 11792 27228
rect 11792 27172 11796 27228
rect 11732 27168 11796 27172
rect 11812 27228 11876 27232
rect 11812 27172 11816 27228
rect 11816 27172 11872 27228
rect 11872 27172 11876 27228
rect 11812 27168 11876 27172
rect 11892 27228 11956 27232
rect 11892 27172 11896 27228
rect 11896 27172 11952 27228
rect 11952 27172 11956 27228
rect 11892 27168 11956 27172
rect 11972 27228 12036 27232
rect 11972 27172 11976 27228
rect 11976 27172 12032 27228
rect 12032 27172 12036 27228
rect 11972 27168 12036 27172
rect 19652 27228 19716 27232
rect 19652 27172 19656 27228
rect 19656 27172 19712 27228
rect 19712 27172 19716 27228
rect 19652 27168 19716 27172
rect 19732 27228 19796 27232
rect 19732 27172 19736 27228
rect 19736 27172 19792 27228
rect 19792 27172 19796 27228
rect 19732 27168 19796 27172
rect 19812 27228 19876 27232
rect 19812 27172 19816 27228
rect 19816 27172 19872 27228
rect 19872 27172 19876 27228
rect 19812 27168 19876 27172
rect 19892 27228 19956 27232
rect 19892 27172 19896 27228
rect 19896 27172 19952 27228
rect 19952 27172 19956 27228
rect 19892 27168 19956 27172
rect 19972 27228 20036 27232
rect 19972 27172 19976 27228
rect 19976 27172 20032 27228
rect 20032 27172 20036 27228
rect 19972 27168 20036 27172
rect 27652 27228 27716 27232
rect 27652 27172 27656 27228
rect 27656 27172 27712 27228
rect 27712 27172 27716 27228
rect 27652 27168 27716 27172
rect 27732 27228 27796 27232
rect 27732 27172 27736 27228
rect 27736 27172 27792 27228
rect 27792 27172 27796 27228
rect 27732 27168 27796 27172
rect 27812 27228 27876 27232
rect 27812 27172 27816 27228
rect 27816 27172 27872 27228
rect 27872 27172 27876 27228
rect 27812 27168 27876 27172
rect 27892 27228 27956 27232
rect 27892 27172 27896 27228
rect 27896 27172 27952 27228
rect 27952 27172 27956 27228
rect 27892 27168 27956 27172
rect 27972 27228 28036 27232
rect 27972 27172 27976 27228
rect 27976 27172 28032 27228
rect 28032 27172 28036 27228
rect 27972 27168 28036 27172
rect 2912 26684 2976 26688
rect 2912 26628 2916 26684
rect 2916 26628 2972 26684
rect 2972 26628 2976 26684
rect 2912 26624 2976 26628
rect 2992 26684 3056 26688
rect 2992 26628 2996 26684
rect 2996 26628 3052 26684
rect 3052 26628 3056 26684
rect 2992 26624 3056 26628
rect 3072 26684 3136 26688
rect 3072 26628 3076 26684
rect 3076 26628 3132 26684
rect 3132 26628 3136 26684
rect 3072 26624 3136 26628
rect 3152 26684 3216 26688
rect 3152 26628 3156 26684
rect 3156 26628 3212 26684
rect 3212 26628 3216 26684
rect 3152 26624 3216 26628
rect 3232 26684 3296 26688
rect 3232 26628 3236 26684
rect 3236 26628 3292 26684
rect 3292 26628 3296 26684
rect 3232 26624 3296 26628
rect 10912 26684 10976 26688
rect 10912 26628 10916 26684
rect 10916 26628 10972 26684
rect 10972 26628 10976 26684
rect 10912 26624 10976 26628
rect 10992 26684 11056 26688
rect 10992 26628 10996 26684
rect 10996 26628 11052 26684
rect 11052 26628 11056 26684
rect 10992 26624 11056 26628
rect 11072 26684 11136 26688
rect 11072 26628 11076 26684
rect 11076 26628 11132 26684
rect 11132 26628 11136 26684
rect 11072 26624 11136 26628
rect 11152 26684 11216 26688
rect 11152 26628 11156 26684
rect 11156 26628 11212 26684
rect 11212 26628 11216 26684
rect 11152 26624 11216 26628
rect 11232 26684 11296 26688
rect 11232 26628 11236 26684
rect 11236 26628 11292 26684
rect 11292 26628 11296 26684
rect 11232 26624 11296 26628
rect 18912 26684 18976 26688
rect 18912 26628 18916 26684
rect 18916 26628 18972 26684
rect 18972 26628 18976 26684
rect 18912 26624 18976 26628
rect 18992 26684 19056 26688
rect 18992 26628 18996 26684
rect 18996 26628 19052 26684
rect 19052 26628 19056 26684
rect 18992 26624 19056 26628
rect 19072 26684 19136 26688
rect 19072 26628 19076 26684
rect 19076 26628 19132 26684
rect 19132 26628 19136 26684
rect 19072 26624 19136 26628
rect 19152 26684 19216 26688
rect 19152 26628 19156 26684
rect 19156 26628 19212 26684
rect 19212 26628 19216 26684
rect 19152 26624 19216 26628
rect 19232 26684 19296 26688
rect 19232 26628 19236 26684
rect 19236 26628 19292 26684
rect 19292 26628 19296 26684
rect 19232 26624 19296 26628
rect 26912 26684 26976 26688
rect 26912 26628 26916 26684
rect 26916 26628 26972 26684
rect 26972 26628 26976 26684
rect 26912 26624 26976 26628
rect 26992 26684 27056 26688
rect 26992 26628 26996 26684
rect 26996 26628 27052 26684
rect 27052 26628 27056 26684
rect 26992 26624 27056 26628
rect 27072 26684 27136 26688
rect 27072 26628 27076 26684
rect 27076 26628 27132 26684
rect 27132 26628 27136 26684
rect 27072 26624 27136 26628
rect 27152 26684 27216 26688
rect 27152 26628 27156 26684
rect 27156 26628 27212 26684
rect 27212 26628 27216 26684
rect 27152 26624 27216 26628
rect 27232 26684 27296 26688
rect 27232 26628 27236 26684
rect 27236 26628 27292 26684
rect 27292 26628 27296 26684
rect 27232 26624 27296 26628
rect 3652 26140 3716 26144
rect 3652 26084 3656 26140
rect 3656 26084 3712 26140
rect 3712 26084 3716 26140
rect 3652 26080 3716 26084
rect 3732 26140 3796 26144
rect 3732 26084 3736 26140
rect 3736 26084 3792 26140
rect 3792 26084 3796 26140
rect 3732 26080 3796 26084
rect 3812 26140 3876 26144
rect 3812 26084 3816 26140
rect 3816 26084 3872 26140
rect 3872 26084 3876 26140
rect 3812 26080 3876 26084
rect 3892 26140 3956 26144
rect 3892 26084 3896 26140
rect 3896 26084 3952 26140
rect 3952 26084 3956 26140
rect 3892 26080 3956 26084
rect 3972 26140 4036 26144
rect 3972 26084 3976 26140
rect 3976 26084 4032 26140
rect 4032 26084 4036 26140
rect 3972 26080 4036 26084
rect 11652 26140 11716 26144
rect 11652 26084 11656 26140
rect 11656 26084 11712 26140
rect 11712 26084 11716 26140
rect 11652 26080 11716 26084
rect 11732 26140 11796 26144
rect 11732 26084 11736 26140
rect 11736 26084 11792 26140
rect 11792 26084 11796 26140
rect 11732 26080 11796 26084
rect 11812 26140 11876 26144
rect 11812 26084 11816 26140
rect 11816 26084 11872 26140
rect 11872 26084 11876 26140
rect 11812 26080 11876 26084
rect 11892 26140 11956 26144
rect 11892 26084 11896 26140
rect 11896 26084 11952 26140
rect 11952 26084 11956 26140
rect 11892 26080 11956 26084
rect 11972 26140 12036 26144
rect 11972 26084 11976 26140
rect 11976 26084 12032 26140
rect 12032 26084 12036 26140
rect 11972 26080 12036 26084
rect 19652 26140 19716 26144
rect 19652 26084 19656 26140
rect 19656 26084 19712 26140
rect 19712 26084 19716 26140
rect 19652 26080 19716 26084
rect 19732 26140 19796 26144
rect 19732 26084 19736 26140
rect 19736 26084 19792 26140
rect 19792 26084 19796 26140
rect 19732 26080 19796 26084
rect 19812 26140 19876 26144
rect 19812 26084 19816 26140
rect 19816 26084 19872 26140
rect 19872 26084 19876 26140
rect 19812 26080 19876 26084
rect 19892 26140 19956 26144
rect 19892 26084 19896 26140
rect 19896 26084 19952 26140
rect 19952 26084 19956 26140
rect 19892 26080 19956 26084
rect 19972 26140 20036 26144
rect 19972 26084 19976 26140
rect 19976 26084 20032 26140
rect 20032 26084 20036 26140
rect 19972 26080 20036 26084
rect 27652 26140 27716 26144
rect 27652 26084 27656 26140
rect 27656 26084 27712 26140
rect 27712 26084 27716 26140
rect 27652 26080 27716 26084
rect 27732 26140 27796 26144
rect 27732 26084 27736 26140
rect 27736 26084 27792 26140
rect 27792 26084 27796 26140
rect 27732 26080 27796 26084
rect 27812 26140 27876 26144
rect 27812 26084 27816 26140
rect 27816 26084 27872 26140
rect 27872 26084 27876 26140
rect 27812 26080 27876 26084
rect 27892 26140 27956 26144
rect 27892 26084 27896 26140
rect 27896 26084 27952 26140
rect 27952 26084 27956 26140
rect 27892 26080 27956 26084
rect 27972 26140 28036 26144
rect 27972 26084 27976 26140
rect 27976 26084 28032 26140
rect 28032 26084 28036 26140
rect 27972 26080 28036 26084
rect 2912 25596 2976 25600
rect 2912 25540 2916 25596
rect 2916 25540 2972 25596
rect 2972 25540 2976 25596
rect 2912 25536 2976 25540
rect 2992 25596 3056 25600
rect 2992 25540 2996 25596
rect 2996 25540 3052 25596
rect 3052 25540 3056 25596
rect 2992 25536 3056 25540
rect 3072 25596 3136 25600
rect 3072 25540 3076 25596
rect 3076 25540 3132 25596
rect 3132 25540 3136 25596
rect 3072 25536 3136 25540
rect 3152 25596 3216 25600
rect 3152 25540 3156 25596
rect 3156 25540 3212 25596
rect 3212 25540 3216 25596
rect 3152 25536 3216 25540
rect 3232 25596 3296 25600
rect 3232 25540 3236 25596
rect 3236 25540 3292 25596
rect 3292 25540 3296 25596
rect 3232 25536 3296 25540
rect 10912 25596 10976 25600
rect 10912 25540 10916 25596
rect 10916 25540 10972 25596
rect 10972 25540 10976 25596
rect 10912 25536 10976 25540
rect 10992 25596 11056 25600
rect 10992 25540 10996 25596
rect 10996 25540 11052 25596
rect 11052 25540 11056 25596
rect 10992 25536 11056 25540
rect 11072 25596 11136 25600
rect 11072 25540 11076 25596
rect 11076 25540 11132 25596
rect 11132 25540 11136 25596
rect 11072 25536 11136 25540
rect 11152 25596 11216 25600
rect 11152 25540 11156 25596
rect 11156 25540 11212 25596
rect 11212 25540 11216 25596
rect 11152 25536 11216 25540
rect 11232 25596 11296 25600
rect 11232 25540 11236 25596
rect 11236 25540 11292 25596
rect 11292 25540 11296 25596
rect 11232 25536 11296 25540
rect 18912 25596 18976 25600
rect 18912 25540 18916 25596
rect 18916 25540 18972 25596
rect 18972 25540 18976 25596
rect 18912 25536 18976 25540
rect 18992 25596 19056 25600
rect 18992 25540 18996 25596
rect 18996 25540 19052 25596
rect 19052 25540 19056 25596
rect 18992 25536 19056 25540
rect 19072 25596 19136 25600
rect 19072 25540 19076 25596
rect 19076 25540 19132 25596
rect 19132 25540 19136 25596
rect 19072 25536 19136 25540
rect 19152 25596 19216 25600
rect 19152 25540 19156 25596
rect 19156 25540 19212 25596
rect 19212 25540 19216 25596
rect 19152 25536 19216 25540
rect 19232 25596 19296 25600
rect 19232 25540 19236 25596
rect 19236 25540 19292 25596
rect 19292 25540 19296 25596
rect 19232 25536 19296 25540
rect 26912 25596 26976 25600
rect 26912 25540 26916 25596
rect 26916 25540 26972 25596
rect 26972 25540 26976 25596
rect 26912 25536 26976 25540
rect 26992 25596 27056 25600
rect 26992 25540 26996 25596
rect 26996 25540 27052 25596
rect 27052 25540 27056 25596
rect 26992 25536 27056 25540
rect 27072 25596 27136 25600
rect 27072 25540 27076 25596
rect 27076 25540 27132 25596
rect 27132 25540 27136 25596
rect 27072 25536 27136 25540
rect 27152 25596 27216 25600
rect 27152 25540 27156 25596
rect 27156 25540 27212 25596
rect 27212 25540 27216 25596
rect 27152 25536 27216 25540
rect 27232 25596 27296 25600
rect 27232 25540 27236 25596
rect 27236 25540 27292 25596
rect 27292 25540 27296 25596
rect 27232 25536 27296 25540
rect 3652 25052 3716 25056
rect 3652 24996 3656 25052
rect 3656 24996 3712 25052
rect 3712 24996 3716 25052
rect 3652 24992 3716 24996
rect 3732 25052 3796 25056
rect 3732 24996 3736 25052
rect 3736 24996 3792 25052
rect 3792 24996 3796 25052
rect 3732 24992 3796 24996
rect 3812 25052 3876 25056
rect 3812 24996 3816 25052
rect 3816 24996 3872 25052
rect 3872 24996 3876 25052
rect 3812 24992 3876 24996
rect 3892 25052 3956 25056
rect 3892 24996 3896 25052
rect 3896 24996 3952 25052
rect 3952 24996 3956 25052
rect 3892 24992 3956 24996
rect 3972 25052 4036 25056
rect 3972 24996 3976 25052
rect 3976 24996 4032 25052
rect 4032 24996 4036 25052
rect 3972 24992 4036 24996
rect 11652 25052 11716 25056
rect 11652 24996 11656 25052
rect 11656 24996 11712 25052
rect 11712 24996 11716 25052
rect 11652 24992 11716 24996
rect 11732 25052 11796 25056
rect 11732 24996 11736 25052
rect 11736 24996 11792 25052
rect 11792 24996 11796 25052
rect 11732 24992 11796 24996
rect 11812 25052 11876 25056
rect 11812 24996 11816 25052
rect 11816 24996 11872 25052
rect 11872 24996 11876 25052
rect 11812 24992 11876 24996
rect 11892 25052 11956 25056
rect 11892 24996 11896 25052
rect 11896 24996 11952 25052
rect 11952 24996 11956 25052
rect 11892 24992 11956 24996
rect 11972 25052 12036 25056
rect 11972 24996 11976 25052
rect 11976 24996 12032 25052
rect 12032 24996 12036 25052
rect 11972 24992 12036 24996
rect 19652 25052 19716 25056
rect 19652 24996 19656 25052
rect 19656 24996 19712 25052
rect 19712 24996 19716 25052
rect 19652 24992 19716 24996
rect 19732 25052 19796 25056
rect 19732 24996 19736 25052
rect 19736 24996 19792 25052
rect 19792 24996 19796 25052
rect 19732 24992 19796 24996
rect 19812 25052 19876 25056
rect 19812 24996 19816 25052
rect 19816 24996 19872 25052
rect 19872 24996 19876 25052
rect 19812 24992 19876 24996
rect 19892 25052 19956 25056
rect 19892 24996 19896 25052
rect 19896 24996 19952 25052
rect 19952 24996 19956 25052
rect 19892 24992 19956 24996
rect 19972 25052 20036 25056
rect 19972 24996 19976 25052
rect 19976 24996 20032 25052
rect 20032 24996 20036 25052
rect 19972 24992 20036 24996
rect 27652 25052 27716 25056
rect 27652 24996 27656 25052
rect 27656 24996 27712 25052
rect 27712 24996 27716 25052
rect 27652 24992 27716 24996
rect 27732 25052 27796 25056
rect 27732 24996 27736 25052
rect 27736 24996 27792 25052
rect 27792 24996 27796 25052
rect 27732 24992 27796 24996
rect 27812 25052 27876 25056
rect 27812 24996 27816 25052
rect 27816 24996 27872 25052
rect 27872 24996 27876 25052
rect 27812 24992 27876 24996
rect 27892 25052 27956 25056
rect 27892 24996 27896 25052
rect 27896 24996 27952 25052
rect 27952 24996 27956 25052
rect 27892 24992 27956 24996
rect 27972 25052 28036 25056
rect 27972 24996 27976 25052
rect 27976 24996 28032 25052
rect 28032 24996 28036 25052
rect 27972 24992 28036 24996
rect 2912 24508 2976 24512
rect 2912 24452 2916 24508
rect 2916 24452 2972 24508
rect 2972 24452 2976 24508
rect 2912 24448 2976 24452
rect 2992 24508 3056 24512
rect 2992 24452 2996 24508
rect 2996 24452 3052 24508
rect 3052 24452 3056 24508
rect 2992 24448 3056 24452
rect 3072 24508 3136 24512
rect 3072 24452 3076 24508
rect 3076 24452 3132 24508
rect 3132 24452 3136 24508
rect 3072 24448 3136 24452
rect 3152 24508 3216 24512
rect 3152 24452 3156 24508
rect 3156 24452 3212 24508
rect 3212 24452 3216 24508
rect 3152 24448 3216 24452
rect 3232 24508 3296 24512
rect 3232 24452 3236 24508
rect 3236 24452 3292 24508
rect 3292 24452 3296 24508
rect 3232 24448 3296 24452
rect 10912 24508 10976 24512
rect 10912 24452 10916 24508
rect 10916 24452 10972 24508
rect 10972 24452 10976 24508
rect 10912 24448 10976 24452
rect 10992 24508 11056 24512
rect 10992 24452 10996 24508
rect 10996 24452 11052 24508
rect 11052 24452 11056 24508
rect 10992 24448 11056 24452
rect 11072 24508 11136 24512
rect 11072 24452 11076 24508
rect 11076 24452 11132 24508
rect 11132 24452 11136 24508
rect 11072 24448 11136 24452
rect 11152 24508 11216 24512
rect 11152 24452 11156 24508
rect 11156 24452 11212 24508
rect 11212 24452 11216 24508
rect 11152 24448 11216 24452
rect 11232 24508 11296 24512
rect 11232 24452 11236 24508
rect 11236 24452 11292 24508
rect 11292 24452 11296 24508
rect 11232 24448 11296 24452
rect 18912 24508 18976 24512
rect 18912 24452 18916 24508
rect 18916 24452 18972 24508
rect 18972 24452 18976 24508
rect 18912 24448 18976 24452
rect 18992 24508 19056 24512
rect 18992 24452 18996 24508
rect 18996 24452 19052 24508
rect 19052 24452 19056 24508
rect 18992 24448 19056 24452
rect 19072 24508 19136 24512
rect 19072 24452 19076 24508
rect 19076 24452 19132 24508
rect 19132 24452 19136 24508
rect 19072 24448 19136 24452
rect 19152 24508 19216 24512
rect 19152 24452 19156 24508
rect 19156 24452 19212 24508
rect 19212 24452 19216 24508
rect 19152 24448 19216 24452
rect 19232 24508 19296 24512
rect 19232 24452 19236 24508
rect 19236 24452 19292 24508
rect 19292 24452 19296 24508
rect 19232 24448 19296 24452
rect 26912 24508 26976 24512
rect 26912 24452 26916 24508
rect 26916 24452 26972 24508
rect 26972 24452 26976 24508
rect 26912 24448 26976 24452
rect 26992 24508 27056 24512
rect 26992 24452 26996 24508
rect 26996 24452 27052 24508
rect 27052 24452 27056 24508
rect 26992 24448 27056 24452
rect 27072 24508 27136 24512
rect 27072 24452 27076 24508
rect 27076 24452 27132 24508
rect 27132 24452 27136 24508
rect 27072 24448 27136 24452
rect 27152 24508 27216 24512
rect 27152 24452 27156 24508
rect 27156 24452 27212 24508
rect 27212 24452 27216 24508
rect 27152 24448 27216 24452
rect 27232 24508 27296 24512
rect 27232 24452 27236 24508
rect 27236 24452 27292 24508
rect 27292 24452 27296 24508
rect 27232 24448 27296 24452
rect 3652 23964 3716 23968
rect 3652 23908 3656 23964
rect 3656 23908 3712 23964
rect 3712 23908 3716 23964
rect 3652 23904 3716 23908
rect 3732 23964 3796 23968
rect 3732 23908 3736 23964
rect 3736 23908 3792 23964
rect 3792 23908 3796 23964
rect 3732 23904 3796 23908
rect 3812 23964 3876 23968
rect 3812 23908 3816 23964
rect 3816 23908 3872 23964
rect 3872 23908 3876 23964
rect 3812 23904 3876 23908
rect 3892 23964 3956 23968
rect 3892 23908 3896 23964
rect 3896 23908 3952 23964
rect 3952 23908 3956 23964
rect 3892 23904 3956 23908
rect 3972 23964 4036 23968
rect 3972 23908 3976 23964
rect 3976 23908 4032 23964
rect 4032 23908 4036 23964
rect 3972 23904 4036 23908
rect 11652 23964 11716 23968
rect 11652 23908 11656 23964
rect 11656 23908 11712 23964
rect 11712 23908 11716 23964
rect 11652 23904 11716 23908
rect 11732 23964 11796 23968
rect 11732 23908 11736 23964
rect 11736 23908 11792 23964
rect 11792 23908 11796 23964
rect 11732 23904 11796 23908
rect 11812 23964 11876 23968
rect 11812 23908 11816 23964
rect 11816 23908 11872 23964
rect 11872 23908 11876 23964
rect 11812 23904 11876 23908
rect 11892 23964 11956 23968
rect 11892 23908 11896 23964
rect 11896 23908 11952 23964
rect 11952 23908 11956 23964
rect 11892 23904 11956 23908
rect 11972 23964 12036 23968
rect 11972 23908 11976 23964
rect 11976 23908 12032 23964
rect 12032 23908 12036 23964
rect 11972 23904 12036 23908
rect 19652 23964 19716 23968
rect 19652 23908 19656 23964
rect 19656 23908 19712 23964
rect 19712 23908 19716 23964
rect 19652 23904 19716 23908
rect 19732 23964 19796 23968
rect 19732 23908 19736 23964
rect 19736 23908 19792 23964
rect 19792 23908 19796 23964
rect 19732 23904 19796 23908
rect 19812 23964 19876 23968
rect 19812 23908 19816 23964
rect 19816 23908 19872 23964
rect 19872 23908 19876 23964
rect 19812 23904 19876 23908
rect 19892 23964 19956 23968
rect 19892 23908 19896 23964
rect 19896 23908 19952 23964
rect 19952 23908 19956 23964
rect 19892 23904 19956 23908
rect 19972 23964 20036 23968
rect 19972 23908 19976 23964
rect 19976 23908 20032 23964
rect 20032 23908 20036 23964
rect 19972 23904 20036 23908
rect 27652 23964 27716 23968
rect 27652 23908 27656 23964
rect 27656 23908 27712 23964
rect 27712 23908 27716 23964
rect 27652 23904 27716 23908
rect 27732 23964 27796 23968
rect 27732 23908 27736 23964
rect 27736 23908 27792 23964
rect 27792 23908 27796 23964
rect 27732 23904 27796 23908
rect 27812 23964 27876 23968
rect 27812 23908 27816 23964
rect 27816 23908 27872 23964
rect 27872 23908 27876 23964
rect 27812 23904 27876 23908
rect 27892 23964 27956 23968
rect 27892 23908 27896 23964
rect 27896 23908 27952 23964
rect 27952 23908 27956 23964
rect 27892 23904 27956 23908
rect 27972 23964 28036 23968
rect 27972 23908 27976 23964
rect 27976 23908 28032 23964
rect 28032 23908 28036 23964
rect 27972 23904 28036 23908
rect 2912 23420 2976 23424
rect 2912 23364 2916 23420
rect 2916 23364 2972 23420
rect 2972 23364 2976 23420
rect 2912 23360 2976 23364
rect 2992 23420 3056 23424
rect 2992 23364 2996 23420
rect 2996 23364 3052 23420
rect 3052 23364 3056 23420
rect 2992 23360 3056 23364
rect 3072 23420 3136 23424
rect 3072 23364 3076 23420
rect 3076 23364 3132 23420
rect 3132 23364 3136 23420
rect 3072 23360 3136 23364
rect 3152 23420 3216 23424
rect 3152 23364 3156 23420
rect 3156 23364 3212 23420
rect 3212 23364 3216 23420
rect 3152 23360 3216 23364
rect 3232 23420 3296 23424
rect 3232 23364 3236 23420
rect 3236 23364 3292 23420
rect 3292 23364 3296 23420
rect 3232 23360 3296 23364
rect 10912 23420 10976 23424
rect 10912 23364 10916 23420
rect 10916 23364 10972 23420
rect 10972 23364 10976 23420
rect 10912 23360 10976 23364
rect 10992 23420 11056 23424
rect 10992 23364 10996 23420
rect 10996 23364 11052 23420
rect 11052 23364 11056 23420
rect 10992 23360 11056 23364
rect 11072 23420 11136 23424
rect 11072 23364 11076 23420
rect 11076 23364 11132 23420
rect 11132 23364 11136 23420
rect 11072 23360 11136 23364
rect 11152 23420 11216 23424
rect 11152 23364 11156 23420
rect 11156 23364 11212 23420
rect 11212 23364 11216 23420
rect 11152 23360 11216 23364
rect 11232 23420 11296 23424
rect 11232 23364 11236 23420
rect 11236 23364 11292 23420
rect 11292 23364 11296 23420
rect 11232 23360 11296 23364
rect 18912 23420 18976 23424
rect 18912 23364 18916 23420
rect 18916 23364 18972 23420
rect 18972 23364 18976 23420
rect 18912 23360 18976 23364
rect 18992 23420 19056 23424
rect 18992 23364 18996 23420
rect 18996 23364 19052 23420
rect 19052 23364 19056 23420
rect 18992 23360 19056 23364
rect 19072 23420 19136 23424
rect 19072 23364 19076 23420
rect 19076 23364 19132 23420
rect 19132 23364 19136 23420
rect 19072 23360 19136 23364
rect 19152 23420 19216 23424
rect 19152 23364 19156 23420
rect 19156 23364 19212 23420
rect 19212 23364 19216 23420
rect 19152 23360 19216 23364
rect 19232 23420 19296 23424
rect 19232 23364 19236 23420
rect 19236 23364 19292 23420
rect 19292 23364 19296 23420
rect 19232 23360 19296 23364
rect 26912 23420 26976 23424
rect 26912 23364 26916 23420
rect 26916 23364 26972 23420
rect 26972 23364 26976 23420
rect 26912 23360 26976 23364
rect 26992 23420 27056 23424
rect 26992 23364 26996 23420
rect 26996 23364 27052 23420
rect 27052 23364 27056 23420
rect 26992 23360 27056 23364
rect 27072 23420 27136 23424
rect 27072 23364 27076 23420
rect 27076 23364 27132 23420
rect 27132 23364 27136 23420
rect 27072 23360 27136 23364
rect 27152 23420 27216 23424
rect 27152 23364 27156 23420
rect 27156 23364 27212 23420
rect 27212 23364 27216 23420
rect 27152 23360 27216 23364
rect 27232 23420 27296 23424
rect 27232 23364 27236 23420
rect 27236 23364 27292 23420
rect 27292 23364 27296 23420
rect 27232 23360 27296 23364
rect 3652 22876 3716 22880
rect 3652 22820 3656 22876
rect 3656 22820 3712 22876
rect 3712 22820 3716 22876
rect 3652 22816 3716 22820
rect 3732 22876 3796 22880
rect 3732 22820 3736 22876
rect 3736 22820 3792 22876
rect 3792 22820 3796 22876
rect 3732 22816 3796 22820
rect 3812 22876 3876 22880
rect 3812 22820 3816 22876
rect 3816 22820 3872 22876
rect 3872 22820 3876 22876
rect 3812 22816 3876 22820
rect 3892 22876 3956 22880
rect 3892 22820 3896 22876
rect 3896 22820 3952 22876
rect 3952 22820 3956 22876
rect 3892 22816 3956 22820
rect 3972 22876 4036 22880
rect 3972 22820 3976 22876
rect 3976 22820 4032 22876
rect 4032 22820 4036 22876
rect 3972 22816 4036 22820
rect 11652 22876 11716 22880
rect 11652 22820 11656 22876
rect 11656 22820 11712 22876
rect 11712 22820 11716 22876
rect 11652 22816 11716 22820
rect 11732 22876 11796 22880
rect 11732 22820 11736 22876
rect 11736 22820 11792 22876
rect 11792 22820 11796 22876
rect 11732 22816 11796 22820
rect 11812 22876 11876 22880
rect 11812 22820 11816 22876
rect 11816 22820 11872 22876
rect 11872 22820 11876 22876
rect 11812 22816 11876 22820
rect 11892 22876 11956 22880
rect 11892 22820 11896 22876
rect 11896 22820 11952 22876
rect 11952 22820 11956 22876
rect 11892 22816 11956 22820
rect 11972 22876 12036 22880
rect 11972 22820 11976 22876
rect 11976 22820 12032 22876
rect 12032 22820 12036 22876
rect 11972 22816 12036 22820
rect 19652 22876 19716 22880
rect 19652 22820 19656 22876
rect 19656 22820 19712 22876
rect 19712 22820 19716 22876
rect 19652 22816 19716 22820
rect 19732 22876 19796 22880
rect 19732 22820 19736 22876
rect 19736 22820 19792 22876
rect 19792 22820 19796 22876
rect 19732 22816 19796 22820
rect 19812 22876 19876 22880
rect 19812 22820 19816 22876
rect 19816 22820 19872 22876
rect 19872 22820 19876 22876
rect 19812 22816 19876 22820
rect 19892 22876 19956 22880
rect 19892 22820 19896 22876
rect 19896 22820 19952 22876
rect 19952 22820 19956 22876
rect 19892 22816 19956 22820
rect 19972 22876 20036 22880
rect 19972 22820 19976 22876
rect 19976 22820 20032 22876
rect 20032 22820 20036 22876
rect 19972 22816 20036 22820
rect 27652 22876 27716 22880
rect 27652 22820 27656 22876
rect 27656 22820 27712 22876
rect 27712 22820 27716 22876
rect 27652 22816 27716 22820
rect 27732 22876 27796 22880
rect 27732 22820 27736 22876
rect 27736 22820 27792 22876
rect 27792 22820 27796 22876
rect 27732 22816 27796 22820
rect 27812 22876 27876 22880
rect 27812 22820 27816 22876
rect 27816 22820 27872 22876
rect 27872 22820 27876 22876
rect 27812 22816 27876 22820
rect 27892 22876 27956 22880
rect 27892 22820 27896 22876
rect 27896 22820 27952 22876
rect 27952 22820 27956 22876
rect 27892 22816 27956 22820
rect 27972 22876 28036 22880
rect 27972 22820 27976 22876
rect 27976 22820 28032 22876
rect 28032 22820 28036 22876
rect 27972 22816 28036 22820
rect 2912 22332 2976 22336
rect 2912 22276 2916 22332
rect 2916 22276 2972 22332
rect 2972 22276 2976 22332
rect 2912 22272 2976 22276
rect 2992 22332 3056 22336
rect 2992 22276 2996 22332
rect 2996 22276 3052 22332
rect 3052 22276 3056 22332
rect 2992 22272 3056 22276
rect 3072 22332 3136 22336
rect 3072 22276 3076 22332
rect 3076 22276 3132 22332
rect 3132 22276 3136 22332
rect 3072 22272 3136 22276
rect 3152 22332 3216 22336
rect 3152 22276 3156 22332
rect 3156 22276 3212 22332
rect 3212 22276 3216 22332
rect 3152 22272 3216 22276
rect 3232 22332 3296 22336
rect 3232 22276 3236 22332
rect 3236 22276 3292 22332
rect 3292 22276 3296 22332
rect 3232 22272 3296 22276
rect 10912 22332 10976 22336
rect 10912 22276 10916 22332
rect 10916 22276 10972 22332
rect 10972 22276 10976 22332
rect 10912 22272 10976 22276
rect 10992 22332 11056 22336
rect 10992 22276 10996 22332
rect 10996 22276 11052 22332
rect 11052 22276 11056 22332
rect 10992 22272 11056 22276
rect 11072 22332 11136 22336
rect 11072 22276 11076 22332
rect 11076 22276 11132 22332
rect 11132 22276 11136 22332
rect 11072 22272 11136 22276
rect 11152 22332 11216 22336
rect 11152 22276 11156 22332
rect 11156 22276 11212 22332
rect 11212 22276 11216 22332
rect 11152 22272 11216 22276
rect 11232 22332 11296 22336
rect 11232 22276 11236 22332
rect 11236 22276 11292 22332
rect 11292 22276 11296 22332
rect 11232 22272 11296 22276
rect 18912 22332 18976 22336
rect 18912 22276 18916 22332
rect 18916 22276 18972 22332
rect 18972 22276 18976 22332
rect 18912 22272 18976 22276
rect 18992 22332 19056 22336
rect 18992 22276 18996 22332
rect 18996 22276 19052 22332
rect 19052 22276 19056 22332
rect 18992 22272 19056 22276
rect 19072 22332 19136 22336
rect 19072 22276 19076 22332
rect 19076 22276 19132 22332
rect 19132 22276 19136 22332
rect 19072 22272 19136 22276
rect 19152 22332 19216 22336
rect 19152 22276 19156 22332
rect 19156 22276 19212 22332
rect 19212 22276 19216 22332
rect 19152 22272 19216 22276
rect 19232 22332 19296 22336
rect 19232 22276 19236 22332
rect 19236 22276 19292 22332
rect 19292 22276 19296 22332
rect 19232 22272 19296 22276
rect 26912 22332 26976 22336
rect 26912 22276 26916 22332
rect 26916 22276 26972 22332
rect 26972 22276 26976 22332
rect 26912 22272 26976 22276
rect 26992 22332 27056 22336
rect 26992 22276 26996 22332
rect 26996 22276 27052 22332
rect 27052 22276 27056 22332
rect 26992 22272 27056 22276
rect 27072 22332 27136 22336
rect 27072 22276 27076 22332
rect 27076 22276 27132 22332
rect 27132 22276 27136 22332
rect 27072 22272 27136 22276
rect 27152 22332 27216 22336
rect 27152 22276 27156 22332
rect 27156 22276 27212 22332
rect 27212 22276 27216 22332
rect 27152 22272 27216 22276
rect 27232 22332 27296 22336
rect 27232 22276 27236 22332
rect 27236 22276 27292 22332
rect 27292 22276 27296 22332
rect 27232 22272 27296 22276
rect 3372 21932 3436 21996
rect 3652 21788 3716 21792
rect 3652 21732 3656 21788
rect 3656 21732 3712 21788
rect 3712 21732 3716 21788
rect 3652 21728 3716 21732
rect 3732 21788 3796 21792
rect 3732 21732 3736 21788
rect 3736 21732 3792 21788
rect 3792 21732 3796 21788
rect 3732 21728 3796 21732
rect 3812 21788 3876 21792
rect 3812 21732 3816 21788
rect 3816 21732 3872 21788
rect 3872 21732 3876 21788
rect 3812 21728 3876 21732
rect 3892 21788 3956 21792
rect 3892 21732 3896 21788
rect 3896 21732 3952 21788
rect 3952 21732 3956 21788
rect 3892 21728 3956 21732
rect 3972 21788 4036 21792
rect 3972 21732 3976 21788
rect 3976 21732 4032 21788
rect 4032 21732 4036 21788
rect 3972 21728 4036 21732
rect 11652 21788 11716 21792
rect 11652 21732 11656 21788
rect 11656 21732 11712 21788
rect 11712 21732 11716 21788
rect 11652 21728 11716 21732
rect 11732 21788 11796 21792
rect 11732 21732 11736 21788
rect 11736 21732 11792 21788
rect 11792 21732 11796 21788
rect 11732 21728 11796 21732
rect 11812 21788 11876 21792
rect 11812 21732 11816 21788
rect 11816 21732 11872 21788
rect 11872 21732 11876 21788
rect 11812 21728 11876 21732
rect 11892 21788 11956 21792
rect 11892 21732 11896 21788
rect 11896 21732 11952 21788
rect 11952 21732 11956 21788
rect 11892 21728 11956 21732
rect 11972 21788 12036 21792
rect 11972 21732 11976 21788
rect 11976 21732 12032 21788
rect 12032 21732 12036 21788
rect 11972 21728 12036 21732
rect 19652 21788 19716 21792
rect 19652 21732 19656 21788
rect 19656 21732 19712 21788
rect 19712 21732 19716 21788
rect 19652 21728 19716 21732
rect 19732 21788 19796 21792
rect 19732 21732 19736 21788
rect 19736 21732 19792 21788
rect 19792 21732 19796 21788
rect 19732 21728 19796 21732
rect 19812 21788 19876 21792
rect 19812 21732 19816 21788
rect 19816 21732 19872 21788
rect 19872 21732 19876 21788
rect 19812 21728 19876 21732
rect 19892 21788 19956 21792
rect 19892 21732 19896 21788
rect 19896 21732 19952 21788
rect 19952 21732 19956 21788
rect 19892 21728 19956 21732
rect 19972 21788 20036 21792
rect 19972 21732 19976 21788
rect 19976 21732 20032 21788
rect 20032 21732 20036 21788
rect 19972 21728 20036 21732
rect 27652 21788 27716 21792
rect 27652 21732 27656 21788
rect 27656 21732 27712 21788
rect 27712 21732 27716 21788
rect 27652 21728 27716 21732
rect 27732 21788 27796 21792
rect 27732 21732 27736 21788
rect 27736 21732 27792 21788
rect 27792 21732 27796 21788
rect 27732 21728 27796 21732
rect 27812 21788 27876 21792
rect 27812 21732 27816 21788
rect 27816 21732 27872 21788
rect 27872 21732 27876 21788
rect 27812 21728 27876 21732
rect 27892 21788 27956 21792
rect 27892 21732 27896 21788
rect 27896 21732 27952 21788
rect 27952 21732 27956 21788
rect 27892 21728 27956 21732
rect 27972 21788 28036 21792
rect 27972 21732 27976 21788
rect 27976 21732 28032 21788
rect 28032 21732 28036 21788
rect 27972 21728 28036 21732
rect 1716 21252 1780 21316
rect 2912 21244 2976 21248
rect 2912 21188 2916 21244
rect 2916 21188 2972 21244
rect 2972 21188 2976 21244
rect 2912 21184 2976 21188
rect 2992 21244 3056 21248
rect 2992 21188 2996 21244
rect 2996 21188 3052 21244
rect 3052 21188 3056 21244
rect 2992 21184 3056 21188
rect 3072 21244 3136 21248
rect 3072 21188 3076 21244
rect 3076 21188 3132 21244
rect 3132 21188 3136 21244
rect 3072 21184 3136 21188
rect 3152 21244 3216 21248
rect 3152 21188 3156 21244
rect 3156 21188 3212 21244
rect 3212 21188 3216 21244
rect 3152 21184 3216 21188
rect 3232 21244 3296 21248
rect 3232 21188 3236 21244
rect 3236 21188 3292 21244
rect 3292 21188 3296 21244
rect 3232 21184 3296 21188
rect 10912 21244 10976 21248
rect 10912 21188 10916 21244
rect 10916 21188 10972 21244
rect 10972 21188 10976 21244
rect 10912 21184 10976 21188
rect 10992 21244 11056 21248
rect 10992 21188 10996 21244
rect 10996 21188 11052 21244
rect 11052 21188 11056 21244
rect 10992 21184 11056 21188
rect 11072 21244 11136 21248
rect 11072 21188 11076 21244
rect 11076 21188 11132 21244
rect 11132 21188 11136 21244
rect 11072 21184 11136 21188
rect 11152 21244 11216 21248
rect 11152 21188 11156 21244
rect 11156 21188 11212 21244
rect 11212 21188 11216 21244
rect 11152 21184 11216 21188
rect 11232 21244 11296 21248
rect 11232 21188 11236 21244
rect 11236 21188 11292 21244
rect 11292 21188 11296 21244
rect 11232 21184 11296 21188
rect 18912 21244 18976 21248
rect 18912 21188 18916 21244
rect 18916 21188 18972 21244
rect 18972 21188 18976 21244
rect 18912 21184 18976 21188
rect 18992 21244 19056 21248
rect 18992 21188 18996 21244
rect 18996 21188 19052 21244
rect 19052 21188 19056 21244
rect 18992 21184 19056 21188
rect 19072 21244 19136 21248
rect 19072 21188 19076 21244
rect 19076 21188 19132 21244
rect 19132 21188 19136 21244
rect 19072 21184 19136 21188
rect 19152 21244 19216 21248
rect 19152 21188 19156 21244
rect 19156 21188 19212 21244
rect 19212 21188 19216 21244
rect 19152 21184 19216 21188
rect 19232 21244 19296 21248
rect 19232 21188 19236 21244
rect 19236 21188 19292 21244
rect 19292 21188 19296 21244
rect 19232 21184 19296 21188
rect 26912 21244 26976 21248
rect 26912 21188 26916 21244
rect 26916 21188 26972 21244
rect 26972 21188 26976 21244
rect 26912 21184 26976 21188
rect 26992 21244 27056 21248
rect 26992 21188 26996 21244
rect 26996 21188 27052 21244
rect 27052 21188 27056 21244
rect 26992 21184 27056 21188
rect 27072 21244 27136 21248
rect 27072 21188 27076 21244
rect 27076 21188 27132 21244
rect 27132 21188 27136 21244
rect 27072 21184 27136 21188
rect 27152 21244 27216 21248
rect 27152 21188 27156 21244
rect 27156 21188 27212 21244
rect 27212 21188 27216 21244
rect 27152 21184 27216 21188
rect 27232 21244 27296 21248
rect 27232 21188 27236 21244
rect 27236 21188 27292 21244
rect 27292 21188 27296 21244
rect 27232 21184 27296 21188
rect 2636 20708 2700 20772
rect 3652 20700 3716 20704
rect 3652 20644 3656 20700
rect 3656 20644 3712 20700
rect 3712 20644 3716 20700
rect 3652 20640 3716 20644
rect 3732 20700 3796 20704
rect 3732 20644 3736 20700
rect 3736 20644 3792 20700
rect 3792 20644 3796 20700
rect 3732 20640 3796 20644
rect 3812 20700 3876 20704
rect 3812 20644 3816 20700
rect 3816 20644 3872 20700
rect 3872 20644 3876 20700
rect 3812 20640 3876 20644
rect 3892 20700 3956 20704
rect 3892 20644 3896 20700
rect 3896 20644 3952 20700
rect 3952 20644 3956 20700
rect 3892 20640 3956 20644
rect 3972 20700 4036 20704
rect 3972 20644 3976 20700
rect 3976 20644 4032 20700
rect 4032 20644 4036 20700
rect 3972 20640 4036 20644
rect 11652 20700 11716 20704
rect 11652 20644 11656 20700
rect 11656 20644 11712 20700
rect 11712 20644 11716 20700
rect 11652 20640 11716 20644
rect 11732 20700 11796 20704
rect 11732 20644 11736 20700
rect 11736 20644 11792 20700
rect 11792 20644 11796 20700
rect 11732 20640 11796 20644
rect 11812 20700 11876 20704
rect 11812 20644 11816 20700
rect 11816 20644 11872 20700
rect 11872 20644 11876 20700
rect 11812 20640 11876 20644
rect 11892 20700 11956 20704
rect 11892 20644 11896 20700
rect 11896 20644 11952 20700
rect 11952 20644 11956 20700
rect 11892 20640 11956 20644
rect 11972 20700 12036 20704
rect 11972 20644 11976 20700
rect 11976 20644 12032 20700
rect 12032 20644 12036 20700
rect 11972 20640 12036 20644
rect 19652 20700 19716 20704
rect 19652 20644 19656 20700
rect 19656 20644 19712 20700
rect 19712 20644 19716 20700
rect 19652 20640 19716 20644
rect 19732 20700 19796 20704
rect 19732 20644 19736 20700
rect 19736 20644 19792 20700
rect 19792 20644 19796 20700
rect 19732 20640 19796 20644
rect 19812 20700 19876 20704
rect 19812 20644 19816 20700
rect 19816 20644 19872 20700
rect 19872 20644 19876 20700
rect 19812 20640 19876 20644
rect 19892 20700 19956 20704
rect 19892 20644 19896 20700
rect 19896 20644 19952 20700
rect 19952 20644 19956 20700
rect 19892 20640 19956 20644
rect 19972 20700 20036 20704
rect 19972 20644 19976 20700
rect 19976 20644 20032 20700
rect 20032 20644 20036 20700
rect 19972 20640 20036 20644
rect 27652 20700 27716 20704
rect 27652 20644 27656 20700
rect 27656 20644 27712 20700
rect 27712 20644 27716 20700
rect 27652 20640 27716 20644
rect 27732 20700 27796 20704
rect 27732 20644 27736 20700
rect 27736 20644 27792 20700
rect 27792 20644 27796 20700
rect 27732 20640 27796 20644
rect 27812 20700 27876 20704
rect 27812 20644 27816 20700
rect 27816 20644 27872 20700
rect 27872 20644 27876 20700
rect 27812 20640 27876 20644
rect 27892 20700 27956 20704
rect 27892 20644 27896 20700
rect 27896 20644 27952 20700
rect 27952 20644 27956 20700
rect 27892 20640 27956 20644
rect 27972 20700 28036 20704
rect 27972 20644 27976 20700
rect 27976 20644 28032 20700
rect 28032 20644 28036 20700
rect 27972 20640 28036 20644
rect 2912 20156 2976 20160
rect 2912 20100 2916 20156
rect 2916 20100 2972 20156
rect 2972 20100 2976 20156
rect 2912 20096 2976 20100
rect 2992 20156 3056 20160
rect 2992 20100 2996 20156
rect 2996 20100 3052 20156
rect 3052 20100 3056 20156
rect 2992 20096 3056 20100
rect 3072 20156 3136 20160
rect 3072 20100 3076 20156
rect 3076 20100 3132 20156
rect 3132 20100 3136 20156
rect 3072 20096 3136 20100
rect 3152 20156 3216 20160
rect 3152 20100 3156 20156
rect 3156 20100 3212 20156
rect 3212 20100 3216 20156
rect 3152 20096 3216 20100
rect 3232 20156 3296 20160
rect 3232 20100 3236 20156
rect 3236 20100 3292 20156
rect 3292 20100 3296 20156
rect 3232 20096 3296 20100
rect 10912 20156 10976 20160
rect 10912 20100 10916 20156
rect 10916 20100 10972 20156
rect 10972 20100 10976 20156
rect 10912 20096 10976 20100
rect 10992 20156 11056 20160
rect 10992 20100 10996 20156
rect 10996 20100 11052 20156
rect 11052 20100 11056 20156
rect 10992 20096 11056 20100
rect 11072 20156 11136 20160
rect 11072 20100 11076 20156
rect 11076 20100 11132 20156
rect 11132 20100 11136 20156
rect 11072 20096 11136 20100
rect 11152 20156 11216 20160
rect 11152 20100 11156 20156
rect 11156 20100 11212 20156
rect 11212 20100 11216 20156
rect 11152 20096 11216 20100
rect 11232 20156 11296 20160
rect 11232 20100 11236 20156
rect 11236 20100 11292 20156
rect 11292 20100 11296 20156
rect 11232 20096 11296 20100
rect 18912 20156 18976 20160
rect 18912 20100 18916 20156
rect 18916 20100 18972 20156
rect 18972 20100 18976 20156
rect 18912 20096 18976 20100
rect 18992 20156 19056 20160
rect 18992 20100 18996 20156
rect 18996 20100 19052 20156
rect 19052 20100 19056 20156
rect 18992 20096 19056 20100
rect 19072 20156 19136 20160
rect 19072 20100 19076 20156
rect 19076 20100 19132 20156
rect 19132 20100 19136 20156
rect 19072 20096 19136 20100
rect 19152 20156 19216 20160
rect 19152 20100 19156 20156
rect 19156 20100 19212 20156
rect 19212 20100 19216 20156
rect 19152 20096 19216 20100
rect 19232 20156 19296 20160
rect 19232 20100 19236 20156
rect 19236 20100 19292 20156
rect 19292 20100 19296 20156
rect 19232 20096 19296 20100
rect 26912 20156 26976 20160
rect 26912 20100 26916 20156
rect 26916 20100 26972 20156
rect 26972 20100 26976 20156
rect 26912 20096 26976 20100
rect 26992 20156 27056 20160
rect 26992 20100 26996 20156
rect 26996 20100 27052 20156
rect 27052 20100 27056 20156
rect 26992 20096 27056 20100
rect 27072 20156 27136 20160
rect 27072 20100 27076 20156
rect 27076 20100 27132 20156
rect 27132 20100 27136 20156
rect 27072 20096 27136 20100
rect 27152 20156 27216 20160
rect 27152 20100 27156 20156
rect 27156 20100 27212 20156
rect 27212 20100 27216 20156
rect 27152 20096 27216 20100
rect 27232 20156 27296 20160
rect 27232 20100 27236 20156
rect 27236 20100 27292 20156
rect 27292 20100 27296 20156
rect 27232 20096 27296 20100
rect 3652 19612 3716 19616
rect 3652 19556 3656 19612
rect 3656 19556 3712 19612
rect 3712 19556 3716 19612
rect 3652 19552 3716 19556
rect 3732 19612 3796 19616
rect 3732 19556 3736 19612
rect 3736 19556 3792 19612
rect 3792 19556 3796 19612
rect 3732 19552 3796 19556
rect 3812 19612 3876 19616
rect 3812 19556 3816 19612
rect 3816 19556 3872 19612
rect 3872 19556 3876 19612
rect 3812 19552 3876 19556
rect 3892 19612 3956 19616
rect 3892 19556 3896 19612
rect 3896 19556 3952 19612
rect 3952 19556 3956 19612
rect 3892 19552 3956 19556
rect 3972 19612 4036 19616
rect 3972 19556 3976 19612
rect 3976 19556 4032 19612
rect 4032 19556 4036 19612
rect 3972 19552 4036 19556
rect 11652 19612 11716 19616
rect 11652 19556 11656 19612
rect 11656 19556 11712 19612
rect 11712 19556 11716 19612
rect 11652 19552 11716 19556
rect 11732 19612 11796 19616
rect 11732 19556 11736 19612
rect 11736 19556 11792 19612
rect 11792 19556 11796 19612
rect 11732 19552 11796 19556
rect 11812 19612 11876 19616
rect 11812 19556 11816 19612
rect 11816 19556 11872 19612
rect 11872 19556 11876 19612
rect 11812 19552 11876 19556
rect 11892 19612 11956 19616
rect 11892 19556 11896 19612
rect 11896 19556 11952 19612
rect 11952 19556 11956 19612
rect 11892 19552 11956 19556
rect 11972 19612 12036 19616
rect 11972 19556 11976 19612
rect 11976 19556 12032 19612
rect 12032 19556 12036 19612
rect 11972 19552 12036 19556
rect 19652 19612 19716 19616
rect 19652 19556 19656 19612
rect 19656 19556 19712 19612
rect 19712 19556 19716 19612
rect 19652 19552 19716 19556
rect 19732 19612 19796 19616
rect 19732 19556 19736 19612
rect 19736 19556 19792 19612
rect 19792 19556 19796 19612
rect 19732 19552 19796 19556
rect 19812 19612 19876 19616
rect 19812 19556 19816 19612
rect 19816 19556 19872 19612
rect 19872 19556 19876 19612
rect 19812 19552 19876 19556
rect 19892 19612 19956 19616
rect 19892 19556 19896 19612
rect 19896 19556 19952 19612
rect 19952 19556 19956 19612
rect 19892 19552 19956 19556
rect 19972 19612 20036 19616
rect 19972 19556 19976 19612
rect 19976 19556 20032 19612
rect 20032 19556 20036 19612
rect 19972 19552 20036 19556
rect 27652 19612 27716 19616
rect 27652 19556 27656 19612
rect 27656 19556 27712 19612
rect 27712 19556 27716 19612
rect 27652 19552 27716 19556
rect 27732 19612 27796 19616
rect 27732 19556 27736 19612
rect 27736 19556 27792 19612
rect 27792 19556 27796 19612
rect 27732 19552 27796 19556
rect 27812 19612 27876 19616
rect 27812 19556 27816 19612
rect 27816 19556 27872 19612
rect 27872 19556 27876 19612
rect 27812 19552 27876 19556
rect 27892 19612 27956 19616
rect 27892 19556 27896 19612
rect 27896 19556 27952 19612
rect 27952 19556 27956 19612
rect 27892 19552 27956 19556
rect 27972 19612 28036 19616
rect 27972 19556 27976 19612
rect 27976 19556 28032 19612
rect 28032 19556 28036 19612
rect 27972 19552 28036 19556
rect 2084 19348 2148 19412
rect 3372 19348 3436 19412
rect 2912 19068 2976 19072
rect 2912 19012 2916 19068
rect 2916 19012 2972 19068
rect 2972 19012 2976 19068
rect 2912 19008 2976 19012
rect 2992 19068 3056 19072
rect 2992 19012 2996 19068
rect 2996 19012 3052 19068
rect 3052 19012 3056 19068
rect 2992 19008 3056 19012
rect 3072 19068 3136 19072
rect 3072 19012 3076 19068
rect 3076 19012 3132 19068
rect 3132 19012 3136 19068
rect 3072 19008 3136 19012
rect 3152 19068 3216 19072
rect 3152 19012 3156 19068
rect 3156 19012 3212 19068
rect 3212 19012 3216 19068
rect 3152 19008 3216 19012
rect 3232 19068 3296 19072
rect 3232 19012 3236 19068
rect 3236 19012 3292 19068
rect 3292 19012 3296 19068
rect 3232 19008 3296 19012
rect 10912 19068 10976 19072
rect 10912 19012 10916 19068
rect 10916 19012 10972 19068
rect 10972 19012 10976 19068
rect 10912 19008 10976 19012
rect 10992 19068 11056 19072
rect 10992 19012 10996 19068
rect 10996 19012 11052 19068
rect 11052 19012 11056 19068
rect 10992 19008 11056 19012
rect 11072 19068 11136 19072
rect 11072 19012 11076 19068
rect 11076 19012 11132 19068
rect 11132 19012 11136 19068
rect 11072 19008 11136 19012
rect 11152 19068 11216 19072
rect 11152 19012 11156 19068
rect 11156 19012 11212 19068
rect 11212 19012 11216 19068
rect 11152 19008 11216 19012
rect 11232 19068 11296 19072
rect 11232 19012 11236 19068
rect 11236 19012 11292 19068
rect 11292 19012 11296 19068
rect 11232 19008 11296 19012
rect 18912 19068 18976 19072
rect 18912 19012 18916 19068
rect 18916 19012 18972 19068
rect 18972 19012 18976 19068
rect 18912 19008 18976 19012
rect 18992 19068 19056 19072
rect 18992 19012 18996 19068
rect 18996 19012 19052 19068
rect 19052 19012 19056 19068
rect 18992 19008 19056 19012
rect 19072 19068 19136 19072
rect 19072 19012 19076 19068
rect 19076 19012 19132 19068
rect 19132 19012 19136 19068
rect 19072 19008 19136 19012
rect 19152 19068 19216 19072
rect 19152 19012 19156 19068
rect 19156 19012 19212 19068
rect 19212 19012 19216 19068
rect 19152 19008 19216 19012
rect 19232 19068 19296 19072
rect 19232 19012 19236 19068
rect 19236 19012 19292 19068
rect 19292 19012 19296 19068
rect 19232 19008 19296 19012
rect 26912 19068 26976 19072
rect 26912 19012 26916 19068
rect 26916 19012 26972 19068
rect 26972 19012 26976 19068
rect 26912 19008 26976 19012
rect 26992 19068 27056 19072
rect 26992 19012 26996 19068
rect 26996 19012 27052 19068
rect 27052 19012 27056 19068
rect 26992 19008 27056 19012
rect 27072 19068 27136 19072
rect 27072 19012 27076 19068
rect 27076 19012 27132 19068
rect 27132 19012 27136 19068
rect 27072 19008 27136 19012
rect 27152 19068 27216 19072
rect 27152 19012 27156 19068
rect 27156 19012 27212 19068
rect 27212 19012 27216 19068
rect 27152 19008 27216 19012
rect 27232 19068 27296 19072
rect 27232 19012 27236 19068
rect 27236 19012 27292 19068
rect 27292 19012 27296 19068
rect 27232 19008 27296 19012
rect 3652 18524 3716 18528
rect 3652 18468 3656 18524
rect 3656 18468 3712 18524
rect 3712 18468 3716 18524
rect 3652 18464 3716 18468
rect 3732 18524 3796 18528
rect 3732 18468 3736 18524
rect 3736 18468 3792 18524
rect 3792 18468 3796 18524
rect 3732 18464 3796 18468
rect 3812 18524 3876 18528
rect 3812 18468 3816 18524
rect 3816 18468 3872 18524
rect 3872 18468 3876 18524
rect 3812 18464 3876 18468
rect 3892 18524 3956 18528
rect 3892 18468 3896 18524
rect 3896 18468 3952 18524
rect 3952 18468 3956 18524
rect 3892 18464 3956 18468
rect 3972 18524 4036 18528
rect 3972 18468 3976 18524
rect 3976 18468 4032 18524
rect 4032 18468 4036 18524
rect 3972 18464 4036 18468
rect 11652 18524 11716 18528
rect 11652 18468 11656 18524
rect 11656 18468 11712 18524
rect 11712 18468 11716 18524
rect 11652 18464 11716 18468
rect 11732 18524 11796 18528
rect 11732 18468 11736 18524
rect 11736 18468 11792 18524
rect 11792 18468 11796 18524
rect 11732 18464 11796 18468
rect 11812 18524 11876 18528
rect 11812 18468 11816 18524
rect 11816 18468 11872 18524
rect 11872 18468 11876 18524
rect 11812 18464 11876 18468
rect 11892 18524 11956 18528
rect 11892 18468 11896 18524
rect 11896 18468 11952 18524
rect 11952 18468 11956 18524
rect 11892 18464 11956 18468
rect 11972 18524 12036 18528
rect 11972 18468 11976 18524
rect 11976 18468 12032 18524
rect 12032 18468 12036 18524
rect 11972 18464 12036 18468
rect 19652 18524 19716 18528
rect 19652 18468 19656 18524
rect 19656 18468 19712 18524
rect 19712 18468 19716 18524
rect 19652 18464 19716 18468
rect 19732 18524 19796 18528
rect 19732 18468 19736 18524
rect 19736 18468 19792 18524
rect 19792 18468 19796 18524
rect 19732 18464 19796 18468
rect 19812 18524 19876 18528
rect 19812 18468 19816 18524
rect 19816 18468 19872 18524
rect 19872 18468 19876 18524
rect 19812 18464 19876 18468
rect 19892 18524 19956 18528
rect 19892 18468 19896 18524
rect 19896 18468 19952 18524
rect 19952 18468 19956 18524
rect 19892 18464 19956 18468
rect 19972 18524 20036 18528
rect 19972 18468 19976 18524
rect 19976 18468 20032 18524
rect 20032 18468 20036 18524
rect 19972 18464 20036 18468
rect 27652 18524 27716 18528
rect 27652 18468 27656 18524
rect 27656 18468 27712 18524
rect 27712 18468 27716 18524
rect 27652 18464 27716 18468
rect 27732 18524 27796 18528
rect 27732 18468 27736 18524
rect 27736 18468 27792 18524
rect 27792 18468 27796 18524
rect 27732 18464 27796 18468
rect 27812 18524 27876 18528
rect 27812 18468 27816 18524
rect 27816 18468 27872 18524
rect 27872 18468 27876 18524
rect 27812 18464 27876 18468
rect 27892 18524 27956 18528
rect 27892 18468 27896 18524
rect 27896 18468 27952 18524
rect 27952 18468 27956 18524
rect 27892 18464 27956 18468
rect 27972 18524 28036 18528
rect 27972 18468 27976 18524
rect 27976 18468 28032 18524
rect 28032 18468 28036 18524
rect 27972 18464 28036 18468
rect 2912 17980 2976 17984
rect 2912 17924 2916 17980
rect 2916 17924 2972 17980
rect 2972 17924 2976 17980
rect 2912 17920 2976 17924
rect 2992 17980 3056 17984
rect 2992 17924 2996 17980
rect 2996 17924 3052 17980
rect 3052 17924 3056 17980
rect 2992 17920 3056 17924
rect 3072 17980 3136 17984
rect 3072 17924 3076 17980
rect 3076 17924 3132 17980
rect 3132 17924 3136 17980
rect 3072 17920 3136 17924
rect 3152 17980 3216 17984
rect 3152 17924 3156 17980
rect 3156 17924 3212 17980
rect 3212 17924 3216 17980
rect 3152 17920 3216 17924
rect 3232 17980 3296 17984
rect 3232 17924 3236 17980
rect 3236 17924 3292 17980
rect 3292 17924 3296 17980
rect 3232 17920 3296 17924
rect 10912 17980 10976 17984
rect 10912 17924 10916 17980
rect 10916 17924 10972 17980
rect 10972 17924 10976 17980
rect 10912 17920 10976 17924
rect 10992 17980 11056 17984
rect 10992 17924 10996 17980
rect 10996 17924 11052 17980
rect 11052 17924 11056 17980
rect 10992 17920 11056 17924
rect 11072 17980 11136 17984
rect 11072 17924 11076 17980
rect 11076 17924 11132 17980
rect 11132 17924 11136 17980
rect 11072 17920 11136 17924
rect 11152 17980 11216 17984
rect 11152 17924 11156 17980
rect 11156 17924 11212 17980
rect 11212 17924 11216 17980
rect 11152 17920 11216 17924
rect 11232 17980 11296 17984
rect 11232 17924 11236 17980
rect 11236 17924 11292 17980
rect 11292 17924 11296 17980
rect 11232 17920 11296 17924
rect 18912 17980 18976 17984
rect 18912 17924 18916 17980
rect 18916 17924 18972 17980
rect 18972 17924 18976 17980
rect 18912 17920 18976 17924
rect 18992 17980 19056 17984
rect 18992 17924 18996 17980
rect 18996 17924 19052 17980
rect 19052 17924 19056 17980
rect 18992 17920 19056 17924
rect 19072 17980 19136 17984
rect 19072 17924 19076 17980
rect 19076 17924 19132 17980
rect 19132 17924 19136 17980
rect 19072 17920 19136 17924
rect 19152 17980 19216 17984
rect 19152 17924 19156 17980
rect 19156 17924 19212 17980
rect 19212 17924 19216 17980
rect 19152 17920 19216 17924
rect 19232 17980 19296 17984
rect 19232 17924 19236 17980
rect 19236 17924 19292 17980
rect 19292 17924 19296 17980
rect 19232 17920 19296 17924
rect 26912 17980 26976 17984
rect 26912 17924 26916 17980
rect 26916 17924 26972 17980
rect 26972 17924 26976 17980
rect 26912 17920 26976 17924
rect 26992 17980 27056 17984
rect 26992 17924 26996 17980
rect 26996 17924 27052 17980
rect 27052 17924 27056 17980
rect 26992 17920 27056 17924
rect 27072 17980 27136 17984
rect 27072 17924 27076 17980
rect 27076 17924 27132 17980
rect 27132 17924 27136 17980
rect 27072 17920 27136 17924
rect 27152 17980 27216 17984
rect 27152 17924 27156 17980
rect 27156 17924 27212 17980
rect 27212 17924 27216 17980
rect 27152 17920 27216 17924
rect 27232 17980 27296 17984
rect 27232 17924 27236 17980
rect 27236 17924 27292 17980
rect 27292 17924 27296 17980
rect 27232 17920 27296 17924
rect 3652 17436 3716 17440
rect 3652 17380 3656 17436
rect 3656 17380 3712 17436
rect 3712 17380 3716 17436
rect 3652 17376 3716 17380
rect 3732 17436 3796 17440
rect 3732 17380 3736 17436
rect 3736 17380 3792 17436
rect 3792 17380 3796 17436
rect 3732 17376 3796 17380
rect 3812 17436 3876 17440
rect 3812 17380 3816 17436
rect 3816 17380 3872 17436
rect 3872 17380 3876 17436
rect 3812 17376 3876 17380
rect 3892 17436 3956 17440
rect 3892 17380 3896 17436
rect 3896 17380 3952 17436
rect 3952 17380 3956 17436
rect 3892 17376 3956 17380
rect 3972 17436 4036 17440
rect 3972 17380 3976 17436
rect 3976 17380 4032 17436
rect 4032 17380 4036 17436
rect 3972 17376 4036 17380
rect 11652 17436 11716 17440
rect 11652 17380 11656 17436
rect 11656 17380 11712 17436
rect 11712 17380 11716 17436
rect 11652 17376 11716 17380
rect 11732 17436 11796 17440
rect 11732 17380 11736 17436
rect 11736 17380 11792 17436
rect 11792 17380 11796 17436
rect 11732 17376 11796 17380
rect 11812 17436 11876 17440
rect 11812 17380 11816 17436
rect 11816 17380 11872 17436
rect 11872 17380 11876 17436
rect 11812 17376 11876 17380
rect 11892 17436 11956 17440
rect 11892 17380 11896 17436
rect 11896 17380 11952 17436
rect 11952 17380 11956 17436
rect 11892 17376 11956 17380
rect 11972 17436 12036 17440
rect 11972 17380 11976 17436
rect 11976 17380 12032 17436
rect 12032 17380 12036 17436
rect 11972 17376 12036 17380
rect 19652 17436 19716 17440
rect 19652 17380 19656 17436
rect 19656 17380 19712 17436
rect 19712 17380 19716 17436
rect 19652 17376 19716 17380
rect 19732 17436 19796 17440
rect 19732 17380 19736 17436
rect 19736 17380 19792 17436
rect 19792 17380 19796 17436
rect 19732 17376 19796 17380
rect 19812 17436 19876 17440
rect 19812 17380 19816 17436
rect 19816 17380 19872 17436
rect 19872 17380 19876 17436
rect 19812 17376 19876 17380
rect 19892 17436 19956 17440
rect 19892 17380 19896 17436
rect 19896 17380 19952 17436
rect 19952 17380 19956 17436
rect 19892 17376 19956 17380
rect 19972 17436 20036 17440
rect 19972 17380 19976 17436
rect 19976 17380 20032 17436
rect 20032 17380 20036 17436
rect 19972 17376 20036 17380
rect 27652 17436 27716 17440
rect 27652 17380 27656 17436
rect 27656 17380 27712 17436
rect 27712 17380 27716 17436
rect 27652 17376 27716 17380
rect 27732 17436 27796 17440
rect 27732 17380 27736 17436
rect 27736 17380 27792 17436
rect 27792 17380 27796 17436
rect 27732 17376 27796 17380
rect 27812 17436 27876 17440
rect 27812 17380 27816 17436
rect 27816 17380 27872 17436
rect 27872 17380 27876 17436
rect 27812 17376 27876 17380
rect 27892 17436 27956 17440
rect 27892 17380 27896 17436
rect 27896 17380 27952 17436
rect 27952 17380 27956 17436
rect 27892 17376 27956 17380
rect 27972 17436 28036 17440
rect 27972 17380 27976 17436
rect 27976 17380 28032 17436
rect 28032 17380 28036 17436
rect 27972 17376 28036 17380
rect 3372 17036 3436 17100
rect 2912 16892 2976 16896
rect 2912 16836 2916 16892
rect 2916 16836 2972 16892
rect 2972 16836 2976 16892
rect 2912 16832 2976 16836
rect 2992 16892 3056 16896
rect 2992 16836 2996 16892
rect 2996 16836 3052 16892
rect 3052 16836 3056 16892
rect 2992 16832 3056 16836
rect 3072 16892 3136 16896
rect 3072 16836 3076 16892
rect 3076 16836 3132 16892
rect 3132 16836 3136 16892
rect 3072 16832 3136 16836
rect 3152 16892 3216 16896
rect 3152 16836 3156 16892
rect 3156 16836 3212 16892
rect 3212 16836 3216 16892
rect 3152 16832 3216 16836
rect 3232 16892 3296 16896
rect 3232 16836 3236 16892
rect 3236 16836 3292 16892
rect 3292 16836 3296 16892
rect 3232 16832 3296 16836
rect 10912 16892 10976 16896
rect 10912 16836 10916 16892
rect 10916 16836 10972 16892
rect 10972 16836 10976 16892
rect 10912 16832 10976 16836
rect 10992 16892 11056 16896
rect 10992 16836 10996 16892
rect 10996 16836 11052 16892
rect 11052 16836 11056 16892
rect 10992 16832 11056 16836
rect 11072 16892 11136 16896
rect 11072 16836 11076 16892
rect 11076 16836 11132 16892
rect 11132 16836 11136 16892
rect 11072 16832 11136 16836
rect 11152 16892 11216 16896
rect 11152 16836 11156 16892
rect 11156 16836 11212 16892
rect 11212 16836 11216 16892
rect 11152 16832 11216 16836
rect 11232 16892 11296 16896
rect 11232 16836 11236 16892
rect 11236 16836 11292 16892
rect 11292 16836 11296 16892
rect 11232 16832 11296 16836
rect 18912 16892 18976 16896
rect 18912 16836 18916 16892
rect 18916 16836 18972 16892
rect 18972 16836 18976 16892
rect 18912 16832 18976 16836
rect 18992 16892 19056 16896
rect 18992 16836 18996 16892
rect 18996 16836 19052 16892
rect 19052 16836 19056 16892
rect 18992 16832 19056 16836
rect 19072 16892 19136 16896
rect 19072 16836 19076 16892
rect 19076 16836 19132 16892
rect 19132 16836 19136 16892
rect 19072 16832 19136 16836
rect 19152 16892 19216 16896
rect 19152 16836 19156 16892
rect 19156 16836 19212 16892
rect 19212 16836 19216 16892
rect 19152 16832 19216 16836
rect 19232 16892 19296 16896
rect 19232 16836 19236 16892
rect 19236 16836 19292 16892
rect 19292 16836 19296 16892
rect 19232 16832 19296 16836
rect 26912 16892 26976 16896
rect 26912 16836 26916 16892
rect 26916 16836 26972 16892
rect 26972 16836 26976 16892
rect 26912 16832 26976 16836
rect 26992 16892 27056 16896
rect 26992 16836 26996 16892
rect 26996 16836 27052 16892
rect 27052 16836 27056 16892
rect 26992 16832 27056 16836
rect 27072 16892 27136 16896
rect 27072 16836 27076 16892
rect 27076 16836 27132 16892
rect 27132 16836 27136 16892
rect 27072 16832 27136 16836
rect 27152 16892 27216 16896
rect 27152 16836 27156 16892
rect 27156 16836 27212 16892
rect 27212 16836 27216 16892
rect 27152 16832 27216 16836
rect 27232 16892 27296 16896
rect 27232 16836 27236 16892
rect 27236 16836 27292 16892
rect 27292 16836 27296 16892
rect 27232 16832 27296 16836
rect 2636 16492 2700 16556
rect 3652 16348 3716 16352
rect 3652 16292 3656 16348
rect 3656 16292 3712 16348
rect 3712 16292 3716 16348
rect 3652 16288 3716 16292
rect 3732 16348 3796 16352
rect 3732 16292 3736 16348
rect 3736 16292 3792 16348
rect 3792 16292 3796 16348
rect 3732 16288 3796 16292
rect 3812 16348 3876 16352
rect 3812 16292 3816 16348
rect 3816 16292 3872 16348
rect 3872 16292 3876 16348
rect 3812 16288 3876 16292
rect 3892 16348 3956 16352
rect 3892 16292 3896 16348
rect 3896 16292 3952 16348
rect 3952 16292 3956 16348
rect 3892 16288 3956 16292
rect 3972 16348 4036 16352
rect 3972 16292 3976 16348
rect 3976 16292 4032 16348
rect 4032 16292 4036 16348
rect 3972 16288 4036 16292
rect 11652 16348 11716 16352
rect 11652 16292 11656 16348
rect 11656 16292 11712 16348
rect 11712 16292 11716 16348
rect 11652 16288 11716 16292
rect 11732 16348 11796 16352
rect 11732 16292 11736 16348
rect 11736 16292 11792 16348
rect 11792 16292 11796 16348
rect 11732 16288 11796 16292
rect 11812 16348 11876 16352
rect 11812 16292 11816 16348
rect 11816 16292 11872 16348
rect 11872 16292 11876 16348
rect 11812 16288 11876 16292
rect 11892 16348 11956 16352
rect 11892 16292 11896 16348
rect 11896 16292 11952 16348
rect 11952 16292 11956 16348
rect 11892 16288 11956 16292
rect 11972 16348 12036 16352
rect 11972 16292 11976 16348
rect 11976 16292 12032 16348
rect 12032 16292 12036 16348
rect 11972 16288 12036 16292
rect 19652 16348 19716 16352
rect 19652 16292 19656 16348
rect 19656 16292 19712 16348
rect 19712 16292 19716 16348
rect 19652 16288 19716 16292
rect 19732 16348 19796 16352
rect 19732 16292 19736 16348
rect 19736 16292 19792 16348
rect 19792 16292 19796 16348
rect 19732 16288 19796 16292
rect 19812 16348 19876 16352
rect 19812 16292 19816 16348
rect 19816 16292 19872 16348
rect 19872 16292 19876 16348
rect 19812 16288 19876 16292
rect 19892 16348 19956 16352
rect 19892 16292 19896 16348
rect 19896 16292 19952 16348
rect 19952 16292 19956 16348
rect 19892 16288 19956 16292
rect 19972 16348 20036 16352
rect 19972 16292 19976 16348
rect 19976 16292 20032 16348
rect 20032 16292 20036 16348
rect 19972 16288 20036 16292
rect 27652 16348 27716 16352
rect 27652 16292 27656 16348
rect 27656 16292 27712 16348
rect 27712 16292 27716 16348
rect 27652 16288 27716 16292
rect 27732 16348 27796 16352
rect 27732 16292 27736 16348
rect 27736 16292 27792 16348
rect 27792 16292 27796 16348
rect 27732 16288 27796 16292
rect 27812 16348 27876 16352
rect 27812 16292 27816 16348
rect 27816 16292 27872 16348
rect 27872 16292 27876 16348
rect 27812 16288 27876 16292
rect 27892 16348 27956 16352
rect 27892 16292 27896 16348
rect 27896 16292 27952 16348
rect 27952 16292 27956 16348
rect 27892 16288 27956 16292
rect 27972 16348 28036 16352
rect 27972 16292 27976 16348
rect 27976 16292 28032 16348
rect 28032 16292 28036 16348
rect 27972 16288 28036 16292
rect 1716 16220 1780 16284
rect 2912 15804 2976 15808
rect 2912 15748 2916 15804
rect 2916 15748 2972 15804
rect 2972 15748 2976 15804
rect 2912 15744 2976 15748
rect 2992 15804 3056 15808
rect 2992 15748 2996 15804
rect 2996 15748 3052 15804
rect 3052 15748 3056 15804
rect 2992 15744 3056 15748
rect 3072 15804 3136 15808
rect 3072 15748 3076 15804
rect 3076 15748 3132 15804
rect 3132 15748 3136 15804
rect 3072 15744 3136 15748
rect 3152 15804 3216 15808
rect 3152 15748 3156 15804
rect 3156 15748 3212 15804
rect 3212 15748 3216 15804
rect 3152 15744 3216 15748
rect 3232 15804 3296 15808
rect 3232 15748 3236 15804
rect 3236 15748 3292 15804
rect 3292 15748 3296 15804
rect 3232 15744 3296 15748
rect 10912 15804 10976 15808
rect 10912 15748 10916 15804
rect 10916 15748 10972 15804
rect 10972 15748 10976 15804
rect 10912 15744 10976 15748
rect 10992 15804 11056 15808
rect 10992 15748 10996 15804
rect 10996 15748 11052 15804
rect 11052 15748 11056 15804
rect 10992 15744 11056 15748
rect 11072 15804 11136 15808
rect 11072 15748 11076 15804
rect 11076 15748 11132 15804
rect 11132 15748 11136 15804
rect 11072 15744 11136 15748
rect 11152 15804 11216 15808
rect 11152 15748 11156 15804
rect 11156 15748 11212 15804
rect 11212 15748 11216 15804
rect 11152 15744 11216 15748
rect 11232 15804 11296 15808
rect 11232 15748 11236 15804
rect 11236 15748 11292 15804
rect 11292 15748 11296 15804
rect 11232 15744 11296 15748
rect 18912 15804 18976 15808
rect 18912 15748 18916 15804
rect 18916 15748 18972 15804
rect 18972 15748 18976 15804
rect 18912 15744 18976 15748
rect 18992 15804 19056 15808
rect 18992 15748 18996 15804
rect 18996 15748 19052 15804
rect 19052 15748 19056 15804
rect 18992 15744 19056 15748
rect 19072 15804 19136 15808
rect 19072 15748 19076 15804
rect 19076 15748 19132 15804
rect 19132 15748 19136 15804
rect 19072 15744 19136 15748
rect 19152 15804 19216 15808
rect 19152 15748 19156 15804
rect 19156 15748 19212 15804
rect 19212 15748 19216 15804
rect 19152 15744 19216 15748
rect 19232 15804 19296 15808
rect 19232 15748 19236 15804
rect 19236 15748 19292 15804
rect 19292 15748 19296 15804
rect 19232 15744 19296 15748
rect 26912 15804 26976 15808
rect 26912 15748 26916 15804
rect 26916 15748 26972 15804
rect 26972 15748 26976 15804
rect 26912 15744 26976 15748
rect 26992 15804 27056 15808
rect 26992 15748 26996 15804
rect 26996 15748 27052 15804
rect 27052 15748 27056 15804
rect 26992 15744 27056 15748
rect 27072 15804 27136 15808
rect 27072 15748 27076 15804
rect 27076 15748 27132 15804
rect 27132 15748 27136 15804
rect 27072 15744 27136 15748
rect 27152 15804 27216 15808
rect 27152 15748 27156 15804
rect 27156 15748 27212 15804
rect 27212 15748 27216 15804
rect 27152 15744 27216 15748
rect 27232 15804 27296 15808
rect 27232 15748 27236 15804
rect 27236 15748 27292 15804
rect 27292 15748 27296 15804
rect 27232 15744 27296 15748
rect 3652 15260 3716 15264
rect 3652 15204 3656 15260
rect 3656 15204 3712 15260
rect 3712 15204 3716 15260
rect 3652 15200 3716 15204
rect 3732 15260 3796 15264
rect 3732 15204 3736 15260
rect 3736 15204 3792 15260
rect 3792 15204 3796 15260
rect 3732 15200 3796 15204
rect 3812 15260 3876 15264
rect 3812 15204 3816 15260
rect 3816 15204 3872 15260
rect 3872 15204 3876 15260
rect 3812 15200 3876 15204
rect 3892 15260 3956 15264
rect 3892 15204 3896 15260
rect 3896 15204 3952 15260
rect 3952 15204 3956 15260
rect 3892 15200 3956 15204
rect 3972 15260 4036 15264
rect 3972 15204 3976 15260
rect 3976 15204 4032 15260
rect 4032 15204 4036 15260
rect 3972 15200 4036 15204
rect 11652 15260 11716 15264
rect 11652 15204 11656 15260
rect 11656 15204 11712 15260
rect 11712 15204 11716 15260
rect 11652 15200 11716 15204
rect 11732 15260 11796 15264
rect 11732 15204 11736 15260
rect 11736 15204 11792 15260
rect 11792 15204 11796 15260
rect 11732 15200 11796 15204
rect 11812 15260 11876 15264
rect 11812 15204 11816 15260
rect 11816 15204 11872 15260
rect 11872 15204 11876 15260
rect 11812 15200 11876 15204
rect 11892 15260 11956 15264
rect 11892 15204 11896 15260
rect 11896 15204 11952 15260
rect 11952 15204 11956 15260
rect 11892 15200 11956 15204
rect 11972 15260 12036 15264
rect 11972 15204 11976 15260
rect 11976 15204 12032 15260
rect 12032 15204 12036 15260
rect 11972 15200 12036 15204
rect 19652 15260 19716 15264
rect 19652 15204 19656 15260
rect 19656 15204 19712 15260
rect 19712 15204 19716 15260
rect 19652 15200 19716 15204
rect 19732 15260 19796 15264
rect 19732 15204 19736 15260
rect 19736 15204 19792 15260
rect 19792 15204 19796 15260
rect 19732 15200 19796 15204
rect 19812 15260 19876 15264
rect 19812 15204 19816 15260
rect 19816 15204 19872 15260
rect 19872 15204 19876 15260
rect 19812 15200 19876 15204
rect 19892 15260 19956 15264
rect 19892 15204 19896 15260
rect 19896 15204 19952 15260
rect 19952 15204 19956 15260
rect 19892 15200 19956 15204
rect 19972 15260 20036 15264
rect 19972 15204 19976 15260
rect 19976 15204 20032 15260
rect 20032 15204 20036 15260
rect 19972 15200 20036 15204
rect 27652 15260 27716 15264
rect 27652 15204 27656 15260
rect 27656 15204 27712 15260
rect 27712 15204 27716 15260
rect 27652 15200 27716 15204
rect 27732 15260 27796 15264
rect 27732 15204 27736 15260
rect 27736 15204 27792 15260
rect 27792 15204 27796 15260
rect 27732 15200 27796 15204
rect 27812 15260 27876 15264
rect 27812 15204 27816 15260
rect 27816 15204 27872 15260
rect 27872 15204 27876 15260
rect 27812 15200 27876 15204
rect 27892 15260 27956 15264
rect 27892 15204 27896 15260
rect 27896 15204 27952 15260
rect 27952 15204 27956 15260
rect 27892 15200 27956 15204
rect 27972 15260 28036 15264
rect 27972 15204 27976 15260
rect 27976 15204 28032 15260
rect 28032 15204 28036 15260
rect 27972 15200 28036 15204
rect 2636 14996 2700 15060
rect 2912 14716 2976 14720
rect 2912 14660 2916 14716
rect 2916 14660 2972 14716
rect 2972 14660 2976 14716
rect 2912 14656 2976 14660
rect 2992 14716 3056 14720
rect 2992 14660 2996 14716
rect 2996 14660 3052 14716
rect 3052 14660 3056 14716
rect 2992 14656 3056 14660
rect 3072 14716 3136 14720
rect 3072 14660 3076 14716
rect 3076 14660 3132 14716
rect 3132 14660 3136 14716
rect 3072 14656 3136 14660
rect 3152 14716 3216 14720
rect 3152 14660 3156 14716
rect 3156 14660 3212 14716
rect 3212 14660 3216 14716
rect 3152 14656 3216 14660
rect 3232 14716 3296 14720
rect 3232 14660 3236 14716
rect 3236 14660 3292 14716
rect 3292 14660 3296 14716
rect 3232 14656 3296 14660
rect 10912 14716 10976 14720
rect 10912 14660 10916 14716
rect 10916 14660 10972 14716
rect 10972 14660 10976 14716
rect 10912 14656 10976 14660
rect 10992 14716 11056 14720
rect 10992 14660 10996 14716
rect 10996 14660 11052 14716
rect 11052 14660 11056 14716
rect 10992 14656 11056 14660
rect 11072 14716 11136 14720
rect 11072 14660 11076 14716
rect 11076 14660 11132 14716
rect 11132 14660 11136 14716
rect 11072 14656 11136 14660
rect 11152 14716 11216 14720
rect 11152 14660 11156 14716
rect 11156 14660 11212 14716
rect 11212 14660 11216 14716
rect 11152 14656 11216 14660
rect 11232 14716 11296 14720
rect 11232 14660 11236 14716
rect 11236 14660 11292 14716
rect 11292 14660 11296 14716
rect 11232 14656 11296 14660
rect 18912 14716 18976 14720
rect 18912 14660 18916 14716
rect 18916 14660 18972 14716
rect 18972 14660 18976 14716
rect 18912 14656 18976 14660
rect 18992 14716 19056 14720
rect 18992 14660 18996 14716
rect 18996 14660 19052 14716
rect 19052 14660 19056 14716
rect 18992 14656 19056 14660
rect 19072 14716 19136 14720
rect 19072 14660 19076 14716
rect 19076 14660 19132 14716
rect 19132 14660 19136 14716
rect 19072 14656 19136 14660
rect 19152 14716 19216 14720
rect 19152 14660 19156 14716
rect 19156 14660 19212 14716
rect 19212 14660 19216 14716
rect 19152 14656 19216 14660
rect 19232 14716 19296 14720
rect 19232 14660 19236 14716
rect 19236 14660 19292 14716
rect 19292 14660 19296 14716
rect 19232 14656 19296 14660
rect 26912 14716 26976 14720
rect 26912 14660 26916 14716
rect 26916 14660 26972 14716
rect 26972 14660 26976 14716
rect 26912 14656 26976 14660
rect 26992 14716 27056 14720
rect 26992 14660 26996 14716
rect 26996 14660 27052 14716
rect 27052 14660 27056 14716
rect 26992 14656 27056 14660
rect 27072 14716 27136 14720
rect 27072 14660 27076 14716
rect 27076 14660 27132 14716
rect 27132 14660 27136 14716
rect 27072 14656 27136 14660
rect 27152 14716 27216 14720
rect 27152 14660 27156 14716
rect 27156 14660 27212 14716
rect 27212 14660 27216 14716
rect 27152 14656 27216 14660
rect 27232 14716 27296 14720
rect 27232 14660 27236 14716
rect 27236 14660 27292 14716
rect 27292 14660 27296 14716
rect 27232 14656 27296 14660
rect 3652 14172 3716 14176
rect 3652 14116 3656 14172
rect 3656 14116 3712 14172
rect 3712 14116 3716 14172
rect 3652 14112 3716 14116
rect 3732 14172 3796 14176
rect 3732 14116 3736 14172
rect 3736 14116 3792 14172
rect 3792 14116 3796 14172
rect 3732 14112 3796 14116
rect 3812 14172 3876 14176
rect 3812 14116 3816 14172
rect 3816 14116 3872 14172
rect 3872 14116 3876 14172
rect 3812 14112 3876 14116
rect 3892 14172 3956 14176
rect 3892 14116 3896 14172
rect 3896 14116 3952 14172
rect 3952 14116 3956 14172
rect 3892 14112 3956 14116
rect 3972 14172 4036 14176
rect 3972 14116 3976 14172
rect 3976 14116 4032 14172
rect 4032 14116 4036 14172
rect 3972 14112 4036 14116
rect 11652 14172 11716 14176
rect 11652 14116 11656 14172
rect 11656 14116 11712 14172
rect 11712 14116 11716 14172
rect 11652 14112 11716 14116
rect 11732 14172 11796 14176
rect 11732 14116 11736 14172
rect 11736 14116 11792 14172
rect 11792 14116 11796 14172
rect 11732 14112 11796 14116
rect 11812 14172 11876 14176
rect 11812 14116 11816 14172
rect 11816 14116 11872 14172
rect 11872 14116 11876 14172
rect 11812 14112 11876 14116
rect 11892 14172 11956 14176
rect 11892 14116 11896 14172
rect 11896 14116 11952 14172
rect 11952 14116 11956 14172
rect 11892 14112 11956 14116
rect 11972 14172 12036 14176
rect 11972 14116 11976 14172
rect 11976 14116 12032 14172
rect 12032 14116 12036 14172
rect 11972 14112 12036 14116
rect 19652 14172 19716 14176
rect 19652 14116 19656 14172
rect 19656 14116 19712 14172
rect 19712 14116 19716 14172
rect 19652 14112 19716 14116
rect 19732 14172 19796 14176
rect 19732 14116 19736 14172
rect 19736 14116 19792 14172
rect 19792 14116 19796 14172
rect 19732 14112 19796 14116
rect 19812 14172 19876 14176
rect 19812 14116 19816 14172
rect 19816 14116 19872 14172
rect 19872 14116 19876 14172
rect 19812 14112 19876 14116
rect 19892 14172 19956 14176
rect 19892 14116 19896 14172
rect 19896 14116 19952 14172
rect 19952 14116 19956 14172
rect 19892 14112 19956 14116
rect 19972 14172 20036 14176
rect 19972 14116 19976 14172
rect 19976 14116 20032 14172
rect 20032 14116 20036 14172
rect 19972 14112 20036 14116
rect 27652 14172 27716 14176
rect 27652 14116 27656 14172
rect 27656 14116 27712 14172
rect 27712 14116 27716 14172
rect 27652 14112 27716 14116
rect 27732 14172 27796 14176
rect 27732 14116 27736 14172
rect 27736 14116 27792 14172
rect 27792 14116 27796 14172
rect 27732 14112 27796 14116
rect 27812 14172 27876 14176
rect 27812 14116 27816 14172
rect 27816 14116 27872 14172
rect 27872 14116 27876 14172
rect 27812 14112 27876 14116
rect 27892 14172 27956 14176
rect 27892 14116 27896 14172
rect 27896 14116 27952 14172
rect 27952 14116 27956 14172
rect 27892 14112 27956 14116
rect 27972 14172 28036 14176
rect 27972 14116 27976 14172
rect 27976 14116 28032 14172
rect 28032 14116 28036 14172
rect 27972 14112 28036 14116
rect 2912 13628 2976 13632
rect 2912 13572 2916 13628
rect 2916 13572 2972 13628
rect 2972 13572 2976 13628
rect 2912 13568 2976 13572
rect 2992 13628 3056 13632
rect 2992 13572 2996 13628
rect 2996 13572 3052 13628
rect 3052 13572 3056 13628
rect 2992 13568 3056 13572
rect 3072 13628 3136 13632
rect 3072 13572 3076 13628
rect 3076 13572 3132 13628
rect 3132 13572 3136 13628
rect 3072 13568 3136 13572
rect 3152 13628 3216 13632
rect 3152 13572 3156 13628
rect 3156 13572 3212 13628
rect 3212 13572 3216 13628
rect 3152 13568 3216 13572
rect 3232 13628 3296 13632
rect 3232 13572 3236 13628
rect 3236 13572 3292 13628
rect 3292 13572 3296 13628
rect 3232 13568 3296 13572
rect 10912 13628 10976 13632
rect 10912 13572 10916 13628
rect 10916 13572 10972 13628
rect 10972 13572 10976 13628
rect 10912 13568 10976 13572
rect 10992 13628 11056 13632
rect 10992 13572 10996 13628
rect 10996 13572 11052 13628
rect 11052 13572 11056 13628
rect 10992 13568 11056 13572
rect 11072 13628 11136 13632
rect 11072 13572 11076 13628
rect 11076 13572 11132 13628
rect 11132 13572 11136 13628
rect 11072 13568 11136 13572
rect 11152 13628 11216 13632
rect 11152 13572 11156 13628
rect 11156 13572 11212 13628
rect 11212 13572 11216 13628
rect 11152 13568 11216 13572
rect 11232 13628 11296 13632
rect 11232 13572 11236 13628
rect 11236 13572 11292 13628
rect 11292 13572 11296 13628
rect 11232 13568 11296 13572
rect 18912 13628 18976 13632
rect 18912 13572 18916 13628
rect 18916 13572 18972 13628
rect 18972 13572 18976 13628
rect 18912 13568 18976 13572
rect 18992 13628 19056 13632
rect 18992 13572 18996 13628
rect 18996 13572 19052 13628
rect 19052 13572 19056 13628
rect 18992 13568 19056 13572
rect 19072 13628 19136 13632
rect 19072 13572 19076 13628
rect 19076 13572 19132 13628
rect 19132 13572 19136 13628
rect 19072 13568 19136 13572
rect 19152 13628 19216 13632
rect 19152 13572 19156 13628
rect 19156 13572 19212 13628
rect 19212 13572 19216 13628
rect 19152 13568 19216 13572
rect 19232 13628 19296 13632
rect 19232 13572 19236 13628
rect 19236 13572 19292 13628
rect 19292 13572 19296 13628
rect 19232 13568 19296 13572
rect 26912 13628 26976 13632
rect 26912 13572 26916 13628
rect 26916 13572 26972 13628
rect 26972 13572 26976 13628
rect 26912 13568 26976 13572
rect 26992 13628 27056 13632
rect 26992 13572 26996 13628
rect 26996 13572 27052 13628
rect 27052 13572 27056 13628
rect 26992 13568 27056 13572
rect 27072 13628 27136 13632
rect 27072 13572 27076 13628
rect 27076 13572 27132 13628
rect 27132 13572 27136 13628
rect 27072 13568 27136 13572
rect 27152 13628 27216 13632
rect 27152 13572 27156 13628
rect 27156 13572 27212 13628
rect 27212 13572 27216 13628
rect 27152 13568 27216 13572
rect 27232 13628 27296 13632
rect 27232 13572 27236 13628
rect 27236 13572 27292 13628
rect 27292 13572 27296 13628
rect 27232 13568 27296 13572
rect 3652 13084 3716 13088
rect 3652 13028 3656 13084
rect 3656 13028 3712 13084
rect 3712 13028 3716 13084
rect 3652 13024 3716 13028
rect 3732 13084 3796 13088
rect 3732 13028 3736 13084
rect 3736 13028 3792 13084
rect 3792 13028 3796 13084
rect 3732 13024 3796 13028
rect 3812 13084 3876 13088
rect 3812 13028 3816 13084
rect 3816 13028 3872 13084
rect 3872 13028 3876 13084
rect 3812 13024 3876 13028
rect 3892 13084 3956 13088
rect 3892 13028 3896 13084
rect 3896 13028 3952 13084
rect 3952 13028 3956 13084
rect 3892 13024 3956 13028
rect 3972 13084 4036 13088
rect 3972 13028 3976 13084
rect 3976 13028 4032 13084
rect 4032 13028 4036 13084
rect 3972 13024 4036 13028
rect 11652 13084 11716 13088
rect 11652 13028 11656 13084
rect 11656 13028 11712 13084
rect 11712 13028 11716 13084
rect 11652 13024 11716 13028
rect 11732 13084 11796 13088
rect 11732 13028 11736 13084
rect 11736 13028 11792 13084
rect 11792 13028 11796 13084
rect 11732 13024 11796 13028
rect 11812 13084 11876 13088
rect 11812 13028 11816 13084
rect 11816 13028 11872 13084
rect 11872 13028 11876 13084
rect 11812 13024 11876 13028
rect 11892 13084 11956 13088
rect 11892 13028 11896 13084
rect 11896 13028 11952 13084
rect 11952 13028 11956 13084
rect 11892 13024 11956 13028
rect 11972 13084 12036 13088
rect 11972 13028 11976 13084
rect 11976 13028 12032 13084
rect 12032 13028 12036 13084
rect 11972 13024 12036 13028
rect 19652 13084 19716 13088
rect 19652 13028 19656 13084
rect 19656 13028 19712 13084
rect 19712 13028 19716 13084
rect 19652 13024 19716 13028
rect 19732 13084 19796 13088
rect 19732 13028 19736 13084
rect 19736 13028 19792 13084
rect 19792 13028 19796 13084
rect 19732 13024 19796 13028
rect 19812 13084 19876 13088
rect 19812 13028 19816 13084
rect 19816 13028 19872 13084
rect 19872 13028 19876 13084
rect 19812 13024 19876 13028
rect 19892 13084 19956 13088
rect 19892 13028 19896 13084
rect 19896 13028 19952 13084
rect 19952 13028 19956 13084
rect 19892 13024 19956 13028
rect 19972 13084 20036 13088
rect 19972 13028 19976 13084
rect 19976 13028 20032 13084
rect 20032 13028 20036 13084
rect 19972 13024 20036 13028
rect 27652 13084 27716 13088
rect 27652 13028 27656 13084
rect 27656 13028 27712 13084
rect 27712 13028 27716 13084
rect 27652 13024 27716 13028
rect 27732 13084 27796 13088
rect 27732 13028 27736 13084
rect 27736 13028 27792 13084
rect 27792 13028 27796 13084
rect 27732 13024 27796 13028
rect 27812 13084 27876 13088
rect 27812 13028 27816 13084
rect 27816 13028 27872 13084
rect 27872 13028 27876 13084
rect 27812 13024 27876 13028
rect 27892 13084 27956 13088
rect 27892 13028 27896 13084
rect 27896 13028 27952 13084
rect 27952 13028 27956 13084
rect 27892 13024 27956 13028
rect 27972 13084 28036 13088
rect 27972 13028 27976 13084
rect 27976 13028 28032 13084
rect 28032 13028 28036 13084
rect 27972 13024 28036 13028
rect 2912 12540 2976 12544
rect 2912 12484 2916 12540
rect 2916 12484 2972 12540
rect 2972 12484 2976 12540
rect 2912 12480 2976 12484
rect 2992 12540 3056 12544
rect 2992 12484 2996 12540
rect 2996 12484 3052 12540
rect 3052 12484 3056 12540
rect 2992 12480 3056 12484
rect 3072 12540 3136 12544
rect 3072 12484 3076 12540
rect 3076 12484 3132 12540
rect 3132 12484 3136 12540
rect 3072 12480 3136 12484
rect 3152 12540 3216 12544
rect 3152 12484 3156 12540
rect 3156 12484 3212 12540
rect 3212 12484 3216 12540
rect 3152 12480 3216 12484
rect 3232 12540 3296 12544
rect 3232 12484 3236 12540
rect 3236 12484 3292 12540
rect 3292 12484 3296 12540
rect 3232 12480 3296 12484
rect 10912 12540 10976 12544
rect 10912 12484 10916 12540
rect 10916 12484 10972 12540
rect 10972 12484 10976 12540
rect 10912 12480 10976 12484
rect 10992 12540 11056 12544
rect 10992 12484 10996 12540
rect 10996 12484 11052 12540
rect 11052 12484 11056 12540
rect 10992 12480 11056 12484
rect 11072 12540 11136 12544
rect 11072 12484 11076 12540
rect 11076 12484 11132 12540
rect 11132 12484 11136 12540
rect 11072 12480 11136 12484
rect 11152 12540 11216 12544
rect 11152 12484 11156 12540
rect 11156 12484 11212 12540
rect 11212 12484 11216 12540
rect 11152 12480 11216 12484
rect 11232 12540 11296 12544
rect 11232 12484 11236 12540
rect 11236 12484 11292 12540
rect 11292 12484 11296 12540
rect 11232 12480 11296 12484
rect 18912 12540 18976 12544
rect 18912 12484 18916 12540
rect 18916 12484 18972 12540
rect 18972 12484 18976 12540
rect 18912 12480 18976 12484
rect 18992 12540 19056 12544
rect 18992 12484 18996 12540
rect 18996 12484 19052 12540
rect 19052 12484 19056 12540
rect 18992 12480 19056 12484
rect 19072 12540 19136 12544
rect 19072 12484 19076 12540
rect 19076 12484 19132 12540
rect 19132 12484 19136 12540
rect 19072 12480 19136 12484
rect 19152 12540 19216 12544
rect 19152 12484 19156 12540
rect 19156 12484 19212 12540
rect 19212 12484 19216 12540
rect 19152 12480 19216 12484
rect 19232 12540 19296 12544
rect 19232 12484 19236 12540
rect 19236 12484 19292 12540
rect 19292 12484 19296 12540
rect 19232 12480 19296 12484
rect 26912 12540 26976 12544
rect 26912 12484 26916 12540
rect 26916 12484 26972 12540
rect 26972 12484 26976 12540
rect 26912 12480 26976 12484
rect 26992 12540 27056 12544
rect 26992 12484 26996 12540
rect 26996 12484 27052 12540
rect 27052 12484 27056 12540
rect 26992 12480 27056 12484
rect 27072 12540 27136 12544
rect 27072 12484 27076 12540
rect 27076 12484 27132 12540
rect 27132 12484 27136 12540
rect 27072 12480 27136 12484
rect 27152 12540 27216 12544
rect 27152 12484 27156 12540
rect 27156 12484 27212 12540
rect 27212 12484 27216 12540
rect 27152 12480 27216 12484
rect 27232 12540 27296 12544
rect 27232 12484 27236 12540
rect 27236 12484 27292 12540
rect 27292 12484 27296 12540
rect 27232 12480 27296 12484
rect 2084 12004 2148 12068
rect 3652 11996 3716 12000
rect 3652 11940 3656 11996
rect 3656 11940 3712 11996
rect 3712 11940 3716 11996
rect 3652 11936 3716 11940
rect 3732 11996 3796 12000
rect 3732 11940 3736 11996
rect 3736 11940 3792 11996
rect 3792 11940 3796 11996
rect 3732 11936 3796 11940
rect 3812 11996 3876 12000
rect 3812 11940 3816 11996
rect 3816 11940 3872 11996
rect 3872 11940 3876 11996
rect 3812 11936 3876 11940
rect 3892 11996 3956 12000
rect 3892 11940 3896 11996
rect 3896 11940 3952 11996
rect 3952 11940 3956 11996
rect 3892 11936 3956 11940
rect 3972 11996 4036 12000
rect 3972 11940 3976 11996
rect 3976 11940 4032 11996
rect 4032 11940 4036 11996
rect 3972 11936 4036 11940
rect 11652 11996 11716 12000
rect 11652 11940 11656 11996
rect 11656 11940 11712 11996
rect 11712 11940 11716 11996
rect 11652 11936 11716 11940
rect 11732 11996 11796 12000
rect 11732 11940 11736 11996
rect 11736 11940 11792 11996
rect 11792 11940 11796 11996
rect 11732 11936 11796 11940
rect 11812 11996 11876 12000
rect 11812 11940 11816 11996
rect 11816 11940 11872 11996
rect 11872 11940 11876 11996
rect 11812 11936 11876 11940
rect 11892 11996 11956 12000
rect 11892 11940 11896 11996
rect 11896 11940 11952 11996
rect 11952 11940 11956 11996
rect 11892 11936 11956 11940
rect 11972 11996 12036 12000
rect 11972 11940 11976 11996
rect 11976 11940 12032 11996
rect 12032 11940 12036 11996
rect 11972 11936 12036 11940
rect 19652 11996 19716 12000
rect 19652 11940 19656 11996
rect 19656 11940 19712 11996
rect 19712 11940 19716 11996
rect 19652 11936 19716 11940
rect 19732 11996 19796 12000
rect 19732 11940 19736 11996
rect 19736 11940 19792 11996
rect 19792 11940 19796 11996
rect 19732 11936 19796 11940
rect 19812 11996 19876 12000
rect 19812 11940 19816 11996
rect 19816 11940 19872 11996
rect 19872 11940 19876 11996
rect 19812 11936 19876 11940
rect 19892 11996 19956 12000
rect 19892 11940 19896 11996
rect 19896 11940 19952 11996
rect 19952 11940 19956 11996
rect 19892 11936 19956 11940
rect 19972 11996 20036 12000
rect 19972 11940 19976 11996
rect 19976 11940 20032 11996
rect 20032 11940 20036 11996
rect 19972 11936 20036 11940
rect 27652 11996 27716 12000
rect 27652 11940 27656 11996
rect 27656 11940 27712 11996
rect 27712 11940 27716 11996
rect 27652 11936 27716 11940
rect 27732 11996 27796 12000
rect 27732 11940 27736 11996
rect 27736 11940 27792 11996
rect 27792 11940 27796 11996
rect 27732 11936 27796 11940
rect 27812 11996 27876 12000
rect 27812 11940 27816 11996
rect 27816 11940 27872 11996
rect 27872 11940 27876 11996
rect 27812 11936 27876 11940
rect 27892 11996 27956 12000
rect 27892 11940 27896 11996
rect 27896 11940 27952 11996
rect 27952 11940 27956 11996
rect 27892 11936 27956 11940
rect 27972 11996 28036 12000
rect 27972 11940 27976 11996
rect 27976 11940 28032 11996
rect 28032 11940 28036 11996
rect 27972 11936 28036 11940
rect 2912 11452 2976 11456
rect 2912 11396 2916 11452
rect 2916 11396 2972 11452
rect 2972 11396 2976 11452
rect 2912 11392 2976 11396
rect 2992 11452 3056 11456
rect 2992 11396 2996 11452
rect 2996 11396 3052 11452
rect 3052 11396 3056 11452
rect 2992 11392 3056 11396
rect 3072 11452 3136 11456
rect 3072 11396 3076 11452
rect 3076 11396 3132 11452
rect 3132 11396 3136 11452
rect 3072 11392 3136 11396
rect 3152 11452 3216 11456
rect 3152 11396 3156 11452
rect 3156 11396 3212 11452
rect 3212 11396 3216 11452
rect 3152 11392 3216 11396
rect 3232 11452 3296 11456
rect 3232 11396 3236 11452
rect 3236 11396 3292 11452
rect 3292 11396 3296 11452
rect 3232 11392 3296 11396
rect 10912 11452 10976 11456
rect 10912 11396 10916 11452
rect 10916 11396 10972 11452
rect 10972 11396 10976 11452
rect 10912 11392 10976 11396
rect 10992 11452 11056 11456
rect 10992 11396 10996 11452
rect 10996 11396 11052 11452
rect 11052 11396 11056 11452
rect 10992 11392 11056 11396
rect 11072 11452 11136 11456
rect 11072 11396 11076 11452
rect 11076 11396 11132 11452
rect 11132 11396 11136 11452
rect 11072 11392 11136 11396
rect 11152 11452 11216 11456
rect 11152 11396 11156 11452
rect 11156 11396 11212 11452
rect 11212 11396 11216 11452
rect 11152 11392 11216 11396
rect 11232 11452 11296 11456
rect 11232 11396 11236 11452
rect 11236 11396 11292 11452
rect 11292 11396 11296 11452
rect 11232 11392 11296 11396
rect 18912 11452 18976 11456
rect 18912 11396 18916 11452
rect 18916 11396 18972 11452
rect 18972 11396 18976 11452
rect 18912 11392 18976 11396
rect 18992 11452 19056 11456
rect 18992 11396 18996 11452
rect 18996 11396 19052 11452
rect 19052 11396 19056 11452
rect 18992 11392 19056 11396
rect 19072 11452 19136 11456
rect 19072 11396 19076 11452
rect 19076 11396 19132 11452
rect 19132 11396 19136 11452
rect 19072 11392 19136 11396
rect 19152 11452 19216 11456
rect 19152 11396 19156 11452
rect 19156 11396 19212 11452
rect 19212 11396 19216 11452
rect 19152 11392 19216 11396
rect 19232 11452 19296 11456
rect 19232 11396 19236 11452
rect 19236 11396 19292 11452
rect 19292 11396 19296 11452
rect 19232 11392 19296 11396
rect 26912 11452 26976 11456
rect 26912 11396 26916 11452
rect 26916 11396 26972 11452
rect 26972 11396 26976 11452
rect 26912 11392 26976 11396
rect 26992 11452 27056 11456
rect 26992 11396 26996 11452
rect 26996 11396 27052 11452
rect 27052 11396 27056 11452
rect 26992 11392 27056 11396
rect 27072 11452 27136 11456
rect 27072 11396 27076 11452
rect 27076 11396 27132 11452
rect 27132 11396 27136 11452
rect 27072 11392 27136 11396
rect 27152 11452 27216 11456
rect 27152 11396 27156 11452
rect 27156 11396 27212 11452
rect 27212 11396 27216 11452
rect 27152 11392 27216 11396
rect 27232 11452 27296 11456
rect 27232 11396 27236 11452
rect 27236 11396 27292 11452
rect 27292 11396 27296 11452
rect 27232 11392 27296 11396
rect 3372 11324 3436 11388
rect 3652 10908 3716 10912
rect 3652 10852 3656 10908
rect 3656 10852 3712 10908
rect 3712 10852 3716 10908
rect 3652 10848 3716 10852
rect 3732 10908 3796 10912
rect 3732 10852 3736 10908
rect 3736 10852 3792 10908
rect 3792 10852 3796 10908
rect 3732 10848 3796 10852
rect 3812 10908 3876 10912
rect 3812 10852 3816 10908
rect 3816 10852 3872 10908
rect 3872 10852 3876 10908
rect 3812 10848 3876 10852
rect 3892 10908 3956 10912
rect 3892 10852 3896 10908
rect 3896 10852 3952 10908
rect 3952 10852 3956 10908
rect 3892 10848 3956 10852
rect 3972 10908 4036 10912
rect 3972 10852 3976 10908
rect 3976 10852 4032 10908
rect 4032 10852 4036 10908
rect 3972 10848 4036 10852
rect 11652 10908 11716 10912
rect 11652 10852 11656 10908
rect 11656 10852 11712 10908
rect 11712 10852 11716 10908
rect 11652 10848 11716 10852
rect 11732 10908 11796 10912
rect 11732 10852 11736 10908
rect 11736 10852 11792 10908
rect 11792 10852 11796 10908
rect 11732 10848 11796 10852
rect 11812 10908 11876 10912
rect 11812 10852 11816 10908
rect 11816 10852 11872 10908
rect 11872 10852 11876 10908
rect 11812 10848 11876 10852
rect 11892 10908 11956 10912
rect 11892 10852 11896 10908
rect 11896 10852 11952 10908
rect 11952 10852 11956 10908
rect 11892 10848 11956 10852
rect 11972 10908 12036 10912
rect 11972 10852 11976 10908
rect 11976 10852 12032 10908
rect 12032 10852 12036 10908
rect 11972 10848 12036 10852
rect 19652 10908 19716 10912
rect 19652 10852 19656 10908
rect 19656 10852 19712 10908
rect 19712 10852 19716 10908
rect 19652 10848 19716 10852
rect 19732 10908 19796 10912
rect 19732 10852 19736 10908
rect 19736 10852 19792 10908
rect 19792 10852 19796 10908
rect 19732 10848 19796 10852
rect 19812 10908 19876 10912
rect 19812 10852 19816 10908
rect 19816 10852 19872 10908
rect 19872 10852 19876 10908
rect 19812 10848 19876 10852
rect 19892 10908 19956 10912
rect 19892 10852 19896 10908
rect 19896 10852 19952 10908
rect 19952 10852 19956 10908
rect 19892 10848 19956 10852
rect 19972 10908 20036 10912
rect 19972 10852 19976 10908
rect 19976 10852 20032 10908
rect 20032 10852 20036 10908
rect 19972 10848 20036 10852
rect 27652 10908 27716 10912
rect 27652 10852 27656 10908
rect 27656 10852 27712 10908
rect 27712 10852 27716 10908
rect 27652 10848 27716 10852
rect 27732 10908 27796 10912
rect 27732 10852 27736 10908
rect 27736 10852 27792 10908
rect 27792 10852 27796 10908
rect 27732 10848 27796 10852
rect 27812 10908 27876 10912
rect 27812 10852 27816 10908
rect 27816 10852 27872 10908
rect 27872 10852 27876 10908
rect 27812 10848 27876 10852
rect 27892 10908 27956 10912
rect 27892 10852 27896 10908
rect 27896 10852 27952 10908
rect 27952 10852 27956 10908
rect 27892 10848 27956 10852
rect 27972 10908 28036 10912
rect 27972 10852 27976 10908
rect 27976 10852 28032 10908
rect 28032 10852 28036 10908
rect 27972 10848 28036 10852
rect 2912 10364 2976 10368
rect 2912 10308 2916 10364
rect 2916 10308 2972 10364
rect 2972 10308 2976 10364
rect 2912 10304 2976 10308
rect 2992 10364 3056 10368
rect 2992 10308 2996 10364
rect 2996 10308 3052 10364
rect 3052 10308 3056 10364
rect 2992 10304 3056 10308
rect 3072 10364 3136 10368
rect 3072 10308 3076 10364
rect 3076 10308 3132 10364
rect 3132 10308 3136 10364
rect 3072 10304 3136 10308
rect 3152 10364 3216 10368
rect 3152 10308 3156 10364
rect 3156 10308 3212 10364
rect 3212 10308 3216 10364
rect 3152 10304 3216 10308
rect 3232 10364 3296 10368
rect 3232 10308 3236 10364
rect 3236 10308 3292 10364
rect 3292 10308 3296 10364
rect 3232 10304 3296 10308
rect 10912 10364 10976 10368
rect 10912 10308 10916 10364
rect 10916 10308 10972 10364
rect 10972 10308 10976 10364
rect 10912 10304 10976 10308
rect 10992 10364 11056 10368
rect 10992 10308 10996 10364
rect 10996 10308 11052 10364
rect 11052 10308 11056 10364
rect 10992 10304 11056 10308
rect 11072 10364 11136 10368
rect 11072 10308 11076 10364
rect 11076 10308 11132 10364
rect 11132 10308 11136 10364
rect 11072 10304 11136 10308
rect 11152 10364 11216 10368
rect 11152 10308 11156 10364
rect 11156 10308 11212 10364
rect 11212 10308 11216 10364
rect 11152 10304 11216 10308
rect 11232 10364 11296 10368
rect 11232 10308 11236 10364
rect 11236 10308 11292 10364
rect 11292 10308 11296 10364
rect 11232 10304 11296 10308
rect 18912 10364 18976 10368
rect 18912 10308 18916 10364
rect 18916 10308 18972 10364
rect 18972 10308 18976 10364
rect 18912 10304 18976 10308
rect 18992 10364 19056 10368
rect 18992 10308 18996 10364
rect 18996 10308 19052 10364
rect 19052 10308 19056 10364
rect 18992 10304 19056 10308
rect 19072 10364 19136 10368
rect 19072 10308 19076 10364
rect 19076 10308 19132 10364
rect 19132 10308 19136 10364
rect 19072 10304 19136 10308
rect 19152 10364 19216 10368
rect 19152 10308 19156 10364
rect 19156 10308 19212 10364
rect 19212 10308 19216 10364
rect 19152 10304 19216 10308
rect 19232 10364 19296 10368
rect 19232 10308 19236 10364
rect 19236 10308 19292 10364
rect 19292 10308 19296 10364
rect 19232 10304 19296 10308
rect 26912 10364 26976 10368
rect 26912 10308 26916 10364
rect 26916 10308 26972 10364
rect 26972 10308 26976 10364
rect 26912 10304 26976 10308
rect 26992 10364 27056 10368
rect 26992 10308 26996 10364
rect 26996 10308 27052 10364
rect 27052 10308 27056 10364
rect 26992 10304 27056 10308
rect 27072 10364 27136 10368
rect 27072 10308 27076 10364
rect 27076 10308 27132 10364
rect 27132 10308 27136 10364
rect 27072 10304 27136 10308
rect 27152 10364 27216 10368
rect 27152 10308 27156 10364
rect 27156 10308 27212 10364
rect 27212 10308 27216 10364
rect 27152 10304 27216 10308
rect 27232 10364 27296 10368
rect 27232 10308 27236 10364
rect 27236 10308 27292 10364
rect 27292 10308 27296 10364
rect 27232 10304 27296 10308
rect 3652 9820 3716 9824
rect 3652 9764 3656 9820
rect 3656 9764 3712 9820
rect 3712 9764 3716 9820
rect 3652 9760 3716 9764
rect 3732 9820 3796 9824
rect 3732 9764 3736 9820
rect 3736 9764 3792 9820
rect 3792 9764 3796 9820
rect 3732 9760 3796 9764
rect 3812 9820 3876 9824
rect 3812 9764 3816 9820
rect 3816 9764 3872 9820
rect 3872 9764 3876 9820
rect 3812 9760 3876 9764
rect 3892 9820 3956 9824
rect 3892 9764 3896 9820
rect 3896 9764 3952 9820
rect 3952 9764 3956 9820
rect 3892 9760 3956 9764
rect 3972 9820 4036 9824
rect 3972 9764 3976 9820
rect 3976 9764 4032 9820
rect 4032 9764 4036 9820
rect 3972 9760 4036 9764
rect 11652 9820 11716 9824
rect 11652 9764 11656 9820
rect 11656 9764 11712 9820
rect 11712 9764 11716 9820
rect 11652 9760 11716 9764
rect 11732 9820 11796 9824
rect 11732 9764 11736 9820
rect 11736 9764 11792 9820
rect 11792 9764 11796 9820
rect 11732 9760 11796 9764
rect 11812 9820 11876 9824
rect 11812 9764 11816 9820
rect 11816 9764 11872 9820
rect 11872 9764 11876 9820
rect 11812 9760 11876 9764
rect 11892 9820 11956 9824
rect 11892 9764 11896 9820
rect 11896 9764 11952 9820
rect 11952 9764 11956 9820
rect 11892 9760 11956 9764
rect 11972 9820 12036 9824
rect 11972 9764 11976 9820
rect 11976 9764 12032 9820
rect 12032 9764 12036 9820
rect 11972 9760 12036 9764
rect 19652 9820 19716 9824
rect 19652 9764 19656 9820
rect 19656 9764 19712 9820
rect 19712 9764 19716 9820
rect 19652 9760 19716 9764
rect 19732 9820 19796 9824
rect 19732 9764 19736 9820
rect 19736 9764 19792 9820
rect 19792 9764 19796 9820
rect 19732 9760 19796 9764
rect 19812 9820 19876 9824
rect 19812 9764 19816 9820
rect 19816 9764 19872 9820
rect 19872 9764 19876 9820
rect 19812 9760 19876 9764
rect 19892 9820 19956 9824
rect 19892 9764 19896 9820
rect 19896 9764 19952 9820
rect 19952 9764 19956 9820
rect 19892 9760 19956 9764
rect 19972 9820 20036 9824
rect 19972 9764 19976 9820
rect 19976 9764 20032 9820
rect 20032 9764 20036 9820
rect 19972 9760 20036 9764
rect 27652 9820 27716 9824
rect 27652 9764 27656 9820
rect 27656 9764 27712 9820
rect 27712 9764 27716 9820
rect 27652 9760 27716 9764
rect 27732 9820 27796 9824
rect 27732 9764 27736 9820
rect 27736 9764 27792 9820
rect 27792 9764 27796 9820
rect 27732 9760 27796 9764
rect 27812 9820 27876 9824
rect 27812 9764 27816 9820
rect 27816 9764 27872 9820
rect 27872 9764 27876 9820
rect 27812 9760 27876 9764
rect 27892 9820 27956 9824
rect 27892 9764 27896 9820
rect 27896 9764 27952 9820
rect 27952 9764 27956 9820
rect 27892 9760 27956 9764
rect 27972 9820 28036 9824
rect 27972 9764 27976 9820
rect 27976 9764 28032 9820
rect 28032 9764 28036 9820
rect 27972 9760 28036 9764
rect 2912 9276 2976 9280
rect 2912 9220 2916 9276
rect 2916 9220 2972 9276
rect 2972 9220 2976 9276
rect 2912 9216 2976 9220
rect 2992 9276 3056 9280
rect 2992 9220 2996 9276
rect 2996 9220 3052 9276
rect 3052 9220 3056 9276
rect 2992 9216 3056 9220
rect 3072 9276 3136 9280
rect 3072 9220 3076 9276
rect 3076 9220 3132 9276
rect 3132 9220 3136 9276
rect 3072 9216 3136 9220
rect 3152 9276 3216 9280
rect 3152 9220 3156 9276
rect 3156 9220 3212 9276
rect 3212 9220 3216 9276
rect 3152 9216 3216 9220
rect 3232 9276 3296 9280
rect 3232 9220 3236 9276
rect 3236 9220 3292 9276
rect 3292 9220 3296 9276
rect 3232 9216 3296 9220
rect 10912 9276 10976 9280
rect 10912 9220 10916 9276
rect 10916 9220 10972 9276
rect 10972 9220 10976 9276
rect 10912 9216 10976 9220
rect 10992 9276 11056 9280
rect 10992 9220 10996 9276
rect 10996 9220 11052 9276
rect 11052 9220 11056 9276
rect 10992 9216 11056 9220
rect 11072 9276 11136 9280
rect 11072 9220 11076 9276
rect 11076 9220 11132 9276
rect 11132 9220 11136 9276
rect 11072 9216 11136 9220
rect 11152 9276 11216 9280
rect 11152 9220 11156 9276
rect 11156 9220 11212 9276
rect 11212 9220 11216 9276
rect 11152 9216 11216 9220
rect 11232 9276 11296 9280
rect 11232 9220 11236 9276
rect 11236 9220 11292 9276
rect 11292 9220 11296 9276
rect 11232 9216 11296 9220
rect 18912 9276 18976 9280
rect 18912 9220 18916 9276
rect 18916 9220 18972 9276
rect 18972 9220 18976 9276
rect 18912 9216 18976 9220
rect 18992 9276 19056 9280
rect 18992 9220 18996 9276
rect 18996 9220 19052 9276
rect 19052 9220 19056 9276
rect 18992 9216 19056 9220
rect 19072 9276 19136 9280
rect 19072 9220 19076 9276
rect 19076 9220 19132 9276
rect 19132 9220 19136 9276
rect 19072 9216 19136 9220
rect 19152 9276 19216 9280
rect 19152 9220 19156 9276
rect 19156 9220 19212 9276
rect 19212 9220 19216 9276
rect 19152 9216 19216 9220
rect 19232 9276 19296 9280
rect 19232 9220 19236 9276
rect 19236 9220 19292 9276
rect 19292 9220 19296 9276
rect 19232 9216 19296 9220
rect 26912 9276 26976 9280
rect 26912 9220 26916 9276
rect 26916 9220 26972 9276
rect 26972 9220 26976 9276
rect 26912 9216 26976 9220
rect 26992 9276 27056 9280
rect 26992 9220 26996 9276
rect 26996 9220 27052 9276
rect 27052 9220 27056 9276
rect 26992 9216 27056 9220
rect 27072 9276 27136 9280
rect 27072 9220 27076 9276
rect 27076 9220 27132 9276
rect 27132 9220 27136 9276
rect 27072 9216 27136 9220
rect 27152 9276 27216 9280
rect 27152 9220 27156 9276
rect 27156 9220 27212 9276
rect 27212 9220 27216 9276
rect 27152 9216 27216 9220
rect 27232 9276 27296 9280
rect 27232 9220 27236 9276
rect 27236 9220 27292 9276
rect 27292 9220 27296 9276
rect 27232 9216 27296 9220
rect 3652 8732 3716 8736
rect 3652 8676 3656 8732
rect 3656 8676 3712 8732
rect 3712 8676 3716 8732
rect 3652 8672 3716 8676
rect 3732 8732 3796 8736
rect 3732 8676 3736 8732
rect 3736 8676 3792 8732
rect 3792 8676 3796 8732
rect 3732 8672 3796 8676
rect 3812 8732 3876 8736
rect 3812 8676 3816 8732
rect 3816 8676 3872 8732
rect 3872 8676 3876 8732
rect 3812 8672 3876 8676
rect 3892 8732 3956 8736
rect 3892 8676 3896 8732
rect 3896 8676 3952 8732
rect 3952 8676 3956 8732
rect 3892 8672 3956 8676
rect 3972 8732 4036 8736
rect 3972 8676 3976 8732
rect 3976 8676 4032 8732
rect 4032 8676 4036 8732
rect 3972 8672 4036 8676
rect 11652 8732 11716 8736
rect 11652 8676 11656 8732
rect 11656 8676 11712 8732
rect 11712 8676 11716 8732
rect 11652 8672 11716 8676
rect 11732 8732 11796 8736
rect 11732 8676 11736 8732
rect 11736 8676 11792 8732
rect 11792 8676 11796 8732
rect 11732 8672 11796 8676
rect 11812 8732 11876 8736
rect 11812 8676 11816 8732
rect 11816 8676 11872 8732
rect 11872 8676 11876 8732
rect 11812 8672 11876 8676
rect 11892 8732 11956 8736
rect 11892 8676 11896 8732
rect 11896 8676 11952 8732
rect 11952 8676 11956 8732
rect 11892 8672 11956 8676
rect 11972 8732 12036 8736
rect 11972 8676 11976 8732
rect 11976 8676 12032 8732
rect 12032 8676 12036 8732
rect 11972 8672 12036 8676
rect 19652 8732 19716 8736
rect 19652 8676 19656 8732
rect 19656 8676 19712 8732
rect 19712 8676 19716 8732
rect 19652 8672 19716 8676
rect 19732 8732 19796 8736
rect 19732 8676 19736 8732
rect 19736 8676 19792 8732
rect 19792 8676 19796 8732
rect 19732 8672 19796 8676
rect 19812 8732 19876 8736
rect 19812 8676 19816 8732
rect 19816 8676 19872 8732
rect 19872 8676 19876 8732
rect 19812 8672 19876 8676
rect 19892 8732 19956 8736
rect 19892 8676 19896 8732
rect 19896 8676 19952 8732
rect 19952 8676 19956 8732
rect 19892 8672 19956 8676
rect 19972 8732 20036 8736
rect 19972 8676 19976 8732
rect 19976 8676 20032 8732
rect 20032 8676 20036 8732
rect 19972 8672 20036 8676
rect 27652 8732 27716 8736
rect 27652 8676 27656 8732
rect 27656 8676 27712 8732
rect 27712 8676 27716 8732
rect 27652 8672 27716 8676
rect 27732 8732 27796 8736
rect 27732 8676 27736 8732
rect 27736 8676 27792 8732
rect 27792 8676 27796 8732
rect 27732 8672 27796 8676
rect 27812 8732 27876 8736
rect 27812 8676 27816 8732
rect 27816 8676 27872 8732
rect 27872 8676 27876 8732
rect 27812 8672 27876 8676
rect 27892 8732 27956 8736
rect 27892 8676 27896 8732
rect 27896 8676 27952 8732
rect 27952 8676 27956 8732
rect 27892 8672 27956 8676
rect 27972 8732 28036 8736
rect 27972 8676 27976 8732
rect 27976 8676 28032 8732
rect 28032 8676 28036 8732
rect 27972 8672 28036 8676
rect 2912 8188 2976 8192
rect 2912 8132 2916 8188
rect 2916 8132 2972 8188
rect 2972 8132 2976 8188
rect 2912 8128 2976 8132
rect 2992 8188 3056 8192
rect 2992 8132 2996 8188
rect 2996 8132 3052 8188
rect 3052 8132 3056 8188
rect 2992 8128 3056 8132
rect 3072 8188 3136 8192
rect 3072 8132 3076 8188
rect 3076 8132 3132 8188
rect 3132 8132 3136 8188
rect 3072 8128 3136 8132
rect 3152 8188 3216 8192
rect 3152 8132 3156 8188
rect 3156 8132 3212 8188
rect 3212 8132 3216 8188
rect 3152 8128 3216 8132
rect 3232 8188 3296 8192
rect 3232 8132 3236 8188
rect 3236 8132 3292 8188
rect 3292 8132 3296 8188
rect 3232 8128 3296 8132
rect 10912 8188 10976 8192
rect 10912 8132 10916 8188
rect 10916 8132 10972 8188
rect 10972 8132 10976 8188
rect 10912 8128 10976 8132
rect 10992 8188 11056 8192
rect 10992 8132 10996 8188
rect 10996 8132 11052 8188
rect 11052 8132 11056 8188
rect 10992 8128 11056 8132
rect 11072 8188 11136 8192
rect 11072 8132 11076 8188
rect 11076 8132 11132 8188
rect 11132 8132 11136 8188
rect 11072 8128 11136 8132
rect 11152 8188 11216 8192
rect 11152 8132 11156 8188
rect 11156 8132 11212 8188
rect 11212 8132 11216 8188
rect 11152 8128 11216 8132
rect 11232 8188 11296 8192
rect 11232 8132 11236 8188
rect 11236 8132 11292 8188
rect 11292 8132 11296 8188
rect 11232 8128 11296 8132
rect 18912 8188 18976 8192
rect 18912 8132 18916 8188
rect 18916 8132 18972 8188
rect 18972 8132 18976 8188
rect 18912 8128 18976 8132
rect 18992 8188 19056 8192
rect 18992 8132 18996 8188
rect 18996 8132 19052 8188
rect 19052 8132 19056 8188
rect 18992 8128 19056 8132
rect 19072 8188 19136 8192
rect 19072 8132 19076 8188
rect 19076 8132 19132 8188
rect 19132 8132 19136 8188
rect 19072 8128 19136 8132
rect 19152 8188 19216 8192
rect 19152 8132 19156 8188
rect 19156 8132 19212 8188
rect 19212 8132 19216 8188
rect 19152 8128 19216 8132
rect 19232 8188 19296 8192
rect 19232 8132 19236 8188
rect 19236 8132 19292 8188
rect 19292 8132 19296 8188
rect 19232 8128 19296 8132
rect 26912 8188 26976 8192
rect 26912 8132 26916 8188
rect 26916 8132 26972 8188
rect 26972 8132 26976 8188
rect 26912 8128 26976 8132
rect 26992 8188 27056 8192
rect 26992 8132 26996 8188
rect 26996 8132 27052 8188
rect 27052 8132 27056 8188
rect 26992 8128 27056 8132
rect 27072 8188 27136 8192
rect 27072 8132 27076 8188
rect 27076 8132 27132 8188
rect 27132 8132 27136 8188
rect 27072 8128 27136 8132
rect 27152 8188 27216 8192
rect 27152 8132 27156 8188
rect 27156 8132 27212 8188
rect 27212 8132 27216 8188
rect 27152 8128 27216 8132
rect 27232 8188 27296 8192
rect 27232 8132 27236 8188
rect 27236 8132 27292 8188
rect 27292 8132 27296 8188
rect 27232 8128 27296 8132
rect 3652 7644 3716 7648
rect 3652 7588 3656 7644
rect 3656 7588 3712 7644
rect 3712 7588 3716 7644
rect 3652 7584 3716 7588
rect 3732 7644 3796 7648
rect 3732 7588 3736 7644
rect 3736 7588 3792 7644
rect 3792 7588 3796 7644
rect 3732 7584 3796 7588
rect 3812 7644 3876 7648
rect 3812 7588 3816 7644
rect 3816 7588 3872 7644
rect 3872 7588 3876 7644
rect 3812 7584 3876 7588
rect 3892 7644 3956 7648
rect 3892 7588 3896 7644
rect 3896 7588 3952 7644
rect 3952 7588 3956 7644
rect 3892 7584 3956 7588
rect 3972 7644 4036 7648
rect 3972 7588 3976 7644
rect 3976 7588 4032 7644
rect 4032 7588 4036 7644
rect 3972 7584 4036 7588
rect 11652 7644 11716 7648
rect 11652 7588 11656 7644
rect 11656 7588 11712 7644
rect 11712 7588 11716 7644
rect 11652 7584 11716 7588
rect 11732 7644 11796 7648
rect 11732 7588 11736 7644
rect 11736 7588 11792 7644
rect 11792 7588 11796 7644
rect 11732 7584 11796 7588
rect 11812 7644 11876 7648
rect 11812 7588 11816 7644
rect 11816 7588 11872 7644
rect 11872 7588 11876 7644
rect 11812 7584 11876 7588
rect 11892 7644 11956 7648
rect 11892 7588 11896 7644
rect 11896 7588 11952 7644
rect 11952 7588 11956 7644
rect 11892 7584 11956 7588
rect 11972 7644 12036 7648
rect 11972 7588 11976 7644
rect 11976 7588 12032 7644
rect 12032 7588 12036 7644
rect 11972 7584 12036 7588
rect 19652 7644 19716 7648
rect 19652 7588 19656 7644
rect 19656 7588 19712 7644
rect 19712 7588 19716 7644
rect 19652 7584 19716 7588
rect 19732 7644 19796 7648
rect 19732 7588 19736 7644
rect 19736 7588 19792 7644
rect 19792 7588 19796 7644
rect 19732 7584 19796 7588
rect 19812 7644 19876 7648
rect 19812 7588 19816 7644
rect 19816 7588 19872 7644
rect 19872 7588 19876 7644
rect 19812 7584 19876 7588
rect 19892 7644 19956 7648
rect 19892 7588 19896 7644
rect 19896 7588 19952 7644
rect 19952 7588 19956 7644
rect 19892 7584 19956 7588
rect 19972 7644 20036 7648
rect 19972 7588 19976 7644
rect 19976 7588 20032 7644
rect 20032 7588 20036 7644
rect 19972 7584 20036 7588
rect 27652 7644 27716 7648
rect 27652 7588 27656 7644
rect 27656 7588 27712 7644
rect 27712 7588 27716 7644
rect 27652 7584 27716 7588
rect 27732 7644 27796 7648
rect 27732 7588 27736 7644
rect 27736 7588 27792 7644
rect 27792 7588 27796 7644
rect 27732 7584 27796 7588
rect 27812 7644 27876 7648
rect 27812 7588 27816 7644
rect 27816 7588 27872 7644
rect 27872 7588 27876 7644
rect 27812 7584 27876 7588
rect 27892 7644 27956 7648
rect 27892 7588 27896 7644
rect 27896 7588 27952 7644
rect 27952 7588 27956 7644
rect 27892 7584 27956 7588
rect 27972 7644 28036 7648
rect 27972 7588 27976 7644
rect 27976 7588 28032 7644
rect 28032 7588 28036 7644
rect 27972 7584 28036 7588
rect 2912 7100 2976 7104
rect 2912 7044 2916 7100
rect 2916 7044 2972 7100
rect 2972 7044 2976 7100
rect 2912 7040 2976 7044
rect 2992 7100 3056 7104
rect 2992 7044 2996 7100
rect 2996 7044 3052 7100
rect 3052 7044 3056 7100
rect 2992 7040 3056 7044
rect 3072 7100 3136 7104
rect 3072 7044 3076 7100
rect 3076 7044 3132 7100
rect 3132 7044 3136 7100
rect 3072 7040 3136 7044
rect 3152 7100 3216 7104
rect 3152 7044 3156 7100
rect 3156 7044 3212 7100
rect 3212 7044 3216 7100
rect 3152 7040 3216 7044
rect 3232 7100 3296 7104
rect 3232 7044 3236 7100
rect 3236 7044 3292 7100
rect 3292 7044 3296 7100
rect 3232 7040 3296 7044
rect 10912 7100 10976 7104
rect 10912 7044 10916 7100
rect 10916 7044 10972 7100
rect 10972 7044 10976 7100
rect 10912 7040 10976 7044
rect 10992 7100 11056 7104
rect 10992 7044 10996 7100
rect 10996 7044 11052 7100
rect 11052 7044 11056 7100
rect 10992 7040 11056 7044
rect 11072 7100 11136 7104
rect 11072 7044 11076 7100
rect 11076 7044 11132 7100
rect 11132 7044 11136 7100
rect 11072 7040 11136 7044
rect 11152 7100 11216 7104
rect 11152 7044 11156 7100
rect 11156 7044 11212 7100
rect 11212 7044 11216 7100
rect 11152 7040 11216 7044
rect 11232 7100 11296 7104
rect 11232 7044 11236 7100
rect 11236 7044 11292 7100
rect 11292 7044 11296 7100
rect 11232 7040 11296 7044
rect 18912 7100 18976 7104
rect 18912 7044 18916 7100
rect 18916 7044 18972 7100
rect 18972 7044 18976 7100
rect 18912 7040 18976 7044
rect 18992 7100 19056 7104
rect 18992 7044 18996 7100
rect 18996 7044 19052 7100
rect 19052 7044 19056 7100
rect 18992 7040 19056 7044
rect 19072 7100 19136 7104
rect 19072 7044 19076 7100
rect 19076 7044 19132 7100
rect 19132 7044 19136 7100
rect 19072 7040 19136 7044
rect 19152 7100 19216 7104
rect 19152 7044 19156 7100
rect 19156 7044 19212 7100
rect 19212 7044 19216 7100
rect 19152 7040 19216 7044
rect 19232 7100 19296 7104
rect 19232 7044 19236 7100
rect 19236 7044 19292 7100
rect 19292 7044 19296 7100
rect 19232 7040 19296 7044
rect 26912 7100 26976 7104
rect 26912 7044 26916 7100
rect 26916 7044 26972 7100
rect 26972 7044 26976 7100
rect 26912 7040 26976 7044
rect 26992 7100 27056 7104
rect 26992 7044 26996 7100
rect 26996 7044 27052 7100
rect 27052 7044 27056 7100
rect 26992 7040 27056 7044
rect 27072 7100 27136 7104
rect 27072 7044 27076 7100
rect 27076 7044 27132 7100
rect 27132 7044 27136 7100
rect 27072 7040 27136 7044
rect 27152 7100 27216 7104
rect 27152 7044 27156 7100
rect 27156 7044 27212 7100
rect 27212 7044 27216 7100
rect 27152 7040 27216 7044
rect 27232 7100 27296 7104
rect 27232 7044 27236 7100
rect 27236 7044 27292 7100
rect 27292 7044 27296 7100
rect 27232 7040 27296 7044
rect 3652 6556 3716 6560
rect 3652 6500 3656 6556
rect 3656 6500 3712 6556
rect 3712 6500 3716 6556
rect 3652 6496 3716 6500
rect 3732 6556 3796 6560
rect 3732 6500 3736 6556
rect 3736 6500 3792 6556
rect 3792 6500 3796 6556
rect 3732 6496 3796 6500
rect 3812 6556 3876 6560
rect 3812 6500 3816 6556
rect 3816 6500 3872 6556
rect 3872 6500 3876 6556
rect 3812 6496 3876 6500
rect 3892 6556 3956 6560
rect 3892 6500 3896 6556
rect 3896 6500 3952 6556
rect 3952 6500 3956 6556
rect 3892 6496 3956 6500
rect 3972 6556 4036 6560
rect 3972 6500 3976 6556
rect 3976 6500 4032 6556
rect 4032 6500 4036 6556
rect 3972 6496 4036 6500
rect 11652 6556 11716 6560
rect 11652 6500 11656 6556
rect 11656 6500 11712 6556
rect 11712 6500 11716 6556
rect 11652 6496 11716 6500
rect 11732 6556 11796 6560
rect 11732 6500 11736 6556
rect 11736 6500 11792 6556
rect 11792 6500 11796 6556
rect 11732 6496 11796 6500
rect 11812 6556 11876 6560
rect 11812 6500 11816 6556
rect 11816 6500 11872 6556
rect 11872 6500 11876 6556
rect 11812 6496 11876 6500
rect 11892 6556 11956 6560
rect 11892 6500 11896 6556
rect 11896 6500 11952 6556
rect 11952 6500 11956 6556
rect 11892 6496 11956 6500
rect 11972 6556 12036 6560
rect 11972 6500 11976 6556
rect 11976 6500 12032 6556
rect 12032 6500 12036 6556
rect 11972 6496 12036 6500
rect 19652 6556 19716 6560
rect 19652 6500 19656 6556
rect 19656 6500 19712 6556
rect 19712 6500 19716 6556
rect 19652 6496 19716 6500
rect 19732 6556 19796 6560
rect 19732 6500 19736 6556
rect 19736 6500 19792 6556
rect 19792 6500 19796 6556
rect 19732 6496 19796 6500
rect 19812 6556 19876 6560
rect 19812 6500 19816 6556
rect 19816 6500 19872 6556
rect 19872 6500 19876 6556
rect 19812 6496 19876 6500
rect 19892 6556 19956 6560
rect 19892 6500 19896 6556
rect 19896 6500 19952 6556
rect 19952 6500 19956 6556
rect 19892 6496 19956 6500
rect 19972 6556 20036 6560
rect 19972 6500 19976 6556
rect 19976 6500 20032 6556
rect 20032 6500 20036 6556
rect 19972 6496 20036 6500
rect 27652 6556 27716 6560
rect 27652 6500 27656 6556
rect 27656 6500 27712 6556
rect 27712 6500 27716 6556
rect 27652 6496 27716 6500
rect 27732 6556 27796 6560
rect 27732 6500 27736 6556
rect 27736 6500 27792 6556
rect 27792 6500 27796 6556
rect 27732 6496 27796 6500
rect 27812 6556 27876 6560
rect 27812 6500 27816 6556
rect 27816 6500 27872 6556
rect 27872 6500 27876 6556
rect 27812 6496 27876 6500
rect 27892 6556 27956 6560
rect 27892 6500 27896 6556
rect 27896 6500 27952 6556
rect 27952 6500 27956 6556
rect 27892 6496 27956 6500
rect 27972 6556 28036 6560
rect 27972 6500 27976 6556
rect 27976 6500 28032 6556
rect 28032 6500 28036 6556
rect 27972 6496 28036 6500
rect 2912 6012 2976 6016
rect 2912 5956 2916 6012
rect 2916 5956 2972 6012
rect 2972 5956 2976 6012
rect 2912 5952 2976 5956
rect 2992 6012 3056 6016
rect 2992 5956 2996 6012
rect 2996 5956 3052 6012
rect 3052 5956 3056 6012
rect 2992 5952 3056 5956
rect 3072 6012 3136 6016
rect 3072 5956 3076 6012
rect 3076 5956 3132 6012
rect 3132 5956 3136 6012
rect 3072 5952 3136 5956
rect 3152 6012 3216 6016
rect 3152 5956 3156 6012
rect 3156 5956 3212 6012
rect 3212 5956 3216 6012
rect 3152 5952 3216 5956
rect 3232 6012 3296 6016
rect 3232 5956 3236 6012
rect 3236 5956 3292 6012
rect 3292 5956 3296 6012
rect 3232 5952 3296 5956
rect 10912 6012 10976 6016
rect 10912 5956 10916 6012
rect 10916 5956 10972 6012
rect 10972 5956 10976 6012
rect 10912 5952 10976 5956
rect 10992 6012 11056 6016
rect 10992 5956 10996 6012
rect 10996 5956 11052 6012
rect 11052 5956 11056 6012
rect 10992 5952 11056 5956
rect 11072 6012 11136 6016
rect 11072 5956 11076 6012
rect 11076 5956 11132 6012
rect 11132 5956 11136 6012
rect 11072 5952 11136 5956
rect 11152 6012 11216 6016
rect 11152 5956 11156 6012
rect 11156 5956 11212 6012
rect 11212 5956 11216 6012
rect 11152 5952 11216 5956
rect 11232 6012 11296 6016
rect 11232 5956 11236 6012
rect 11236 5956 11292 6012
rect 11292 5956 11296 6012
rect 11232 5952 11296 5956
rect 18912 6012 18976 6016
rect 18912 5956 18916 6012
rect 18916 5956 18972 6012
rect 18972 5956 18976 6012
rect 18912 5952 18976 5956
rect 18992 6012 19056 6016
rect 18992 5956 18996 6012
rect 18996 5956 19052 6012
rect 19052 5956 19056 6012
rect 18992 5952 19056 5956
rect 19072 6012 19136 6016
rect 19072 5956 19076 6012
rect 19076 5956 19132 6012
rect 19132 5956 19136 6012
rect 19072 5952 19136 5956
rect 19152 6012 19216 6016
rect 19152 5956 19156 6012
rect 19156 5956 19212 6012
rect 19212 5956 19216 6012
rect 19152 5952 19216 5956
rect 19232 6012 19296 6016
rect 19232 5956 19236 6012
rect 19236 5956 19292 6012
rect 19292 5956 19296 6012
rect 19232 5952 19296 5956
rect 26912 6012 26976 6016
rect 26912 5956 26916 6012
rect 26916 5956 26972 6012
rect 26972 5956 26976 6012
rect 26912 5952 26976 5956
rect 26992 6012 27056 6016
rect 26992 5956 26996 6012
rect 26996 5956 27052 6012
rect 27052 5956 27056 6012
rect 26992 5952 27056 5956
rect 27072 6012 27136 6016
rect 27072 5956 27076 6012
rect 27076 5956 27132 6012
rect 27132 5956 27136 6012
rect 27072 5952 27136 5956
rect 27152 6012 27216 6016
rect 27152 5956 27156 6012
rect 27156 5956 27212 6012
rect 27212 5956 27216 6012
rect 27152 5952 27216 5956
rect 27232 6012 27296 6016
rect 27232 5956 27236 6012
rect 27236 5956 27292 6012
rect 27292 5956 27296 6012
rect 27232 5952 27296 5956
rect 3652 5468 3716 5472
rect 3652 5412 3656 5468
rect 3656 5412 3712 5468
rect 3712 5412 3716 5468
rect 3652 5408 3716 5412
rect 3732 5468 3796 5472
rect 3732 5412 3736 5468
rect 3736 5412 3792 5468
rect 3792 5412 3796 5468
rect 3732 5408 3796 5412
rect 3812 5468 3876 5472
rect 3812 5412 3816 5468
rect 3816 5412 3872 5468
rect 3872 5412 3876 5468
rect 3812 5408 3876 5412
rect 3892 5468 3956 5472
rect 3892 5412 3896 5468
rect 3896 5412 3952 5468
rect 3952 5412 3956 5468
rect 3892 5408 3956 5412
rect 3972 5468 4036 5472
rect 3972 5412 3976 5468
rect 3976 5412 4032 5468
rect 4032 5412 4036 5468
rect 3972 5408 4036 5412
rect 11652 5468 11716 5472
rect 11652 5412 11656 5468
rect 11656 5412 11712 5468
rect 11712 5412 11716 5468
rect 11652 5408 11716 5412
rect 11732 5468 11796 5472
rect 11732 5412 11736 5468
rect 11736 5412 11792 5468
rect 11792 5412 11796 5468
rect 11732 5408 11796 5412
rect 11812 5468 11876 5472
rect 11812 5412 11816 5468
rect 11816 5412 11872 5468
rect 11872 5412 11876 5468
rect 11812 5408 11876 5412
rect 11892 5468 11956 5472
rect 11892 5412 11896 5468
rect 11896 5412 11952 5468
rect 11952 5412 11956 5468
rect 11892 5408 11956 5412
rect 11972 5468 12036 5472
rect 11972 5412 11976 5468
rect 11976 5412 12032 5468
rect 12032 5412 12036 5468
rect 11972 5408 12036 5412
rect 19652 5468 19716 5472
rect 19652 5412 19656 5468
rect 19656 5412 19712 5468
rect 19712 5412 19716 5468
rect 19652 5408 19716 5412
rect 19732 5468 19796 5472
rect 19732 5412 19736 5468
rect 19736 5412 19792 5468
rect 19792 5412 19796 5468
rect 19732 5408 19796 5412
rect 19812 5468 19876 5472
rect 19812 5412 19816 5468
rect 19816 5412 19872 5468
rect 19872 5412 19876 5468
rect 19812 5408 19876 5412
rect 19892 5468 19956 5472
rect 19892 5412 19896 5468
rect 19896 5412 19952 5468
rect 19952 5412 19956 5468
rect 19892 5408 19956 5412
rect 19972 5468 20036 5472
rect 19972 5412 19976 5468
rect 19976 5412 20032 5468
rect 20032 5412 20036 5468
rect 19972 5408 20036 5412
rect 27652 5468 27716 5472
rect 27652 5412 27656 5468
rect 27656 5412 27712 5468
rect 27712 5412 27716 5468
rect 27652 5408 27716 5412
rect 27732 5468 27796 5472
rect 27732 5412 27736 5468
rect 27736 5412 27792 5468
rect 27792 5412 27796 5468
rect 27732 5408 27796 5412
rect 27812 5468 27876 5472
rect 27812 5412 27816 5468
rect 27816 5412 27872 5468
rect 27872 5412 27876 5468
rect 27812 5408 27876 5412
rect 27892 5468 27956 5472
rect 27892 5412 27896 5468
rect 27896 5412 27952 5468
rect 27952 5412 27956 5468
rect 27892 5408 27956 5412
rect 27972 5468 28036 5472
rect 27972 5412 27976 5468
rect 27976 5412 28032 5468
rect 28032 5412 28036 5468
rect 27972 5408 28036 5412
rect 2912 4924 2976 4928
rect 2912 4868 2916 4924
rect 2916 4868 2972 4924
rect 2972 4868 2976 4924
rect 2912 4864 2976 4868
rect 2992 4924 3056 4928
rect 2992 4868 2996 4924
rect 2996 4868 3052 4924
rect 3052 4868 3056 4924
rect 2992 4864 3056 4868
rect 3072 4924 3136 4928
rect 3072 4868 3076 4924
rect 3076 4868 3132 4924
rect 3132 4868 3136 4924
rect 3072 4864 3136 4868
rect 3152 4924 3216 4928
rect 3152 4868 3156 4924
rect 3156 4868 3212 4924
rect 3212 4868 3216 4924
rect 3152 4864 3216 4868
rect 3232 4924 3296 4928
rect 3232 4868 3236 4924
rect 3236 4868 3292 4924
rect 3292 4868 3296 4924
rect 3232 4864 3296 4868
rect 10912 4924 10976 4928
rect 10912 4868 10916 4924
rect 10916 4868 10972 4924
rect 10972 4868 10976 4924
rect 10912 4864 10976 4868
rect 10992 4924 11056 4928
rect 10992 4868 10996 4924
rect 10996 4868 11052 4924
rect 11052 4868 11056 4924
rect 10992 4864 11056 4868
rect 11072 4924 11136 4928
rect 11072 4868 11076 4924
rect 11076 4868 11132 4924
rect 11132 4868 11136 4924
rect 11072 4864 11136 4868
rect 11152 4924 11216 4928
rect 11152 4868 11156 4924
rect 11156 4868 11212 4924
rect 11212 4868 11216 4924
rect 11152 4864 11216 4868
rect 11232 4924 11296 4928
rect 11232 4868 11236 4924
rect 11236 4868 11292 4924
rect 11292 4868 11296 4924
rect 11232 4864 11296 4868
rect 18912 4924 18976 4928
rect 18912 4868 18916 4924
rect 18916 4868 18972 4924
rect 18972 4868 18976 4924
rect 18912 4864 18976 4868
rect 18992 4924 19056 4928
rect 18992 4868 18996 4924
rect 18996 4868 19052 4924
rect 19052 4868 19056 4924
rect 18992 4864 19056 4868
rect 19072 4924 19136 4928
rect 19072 4868 19076 4924
rect 19076 4868 19132 4924
rect 19132 4868 19136 4924
rect 19072 4864 19136 4868
rect 19152 4924 19216 4928
rect 19152 4868 19156 4924
rect 19156 4868 19212 4924
rect 19212 4868 19216 4924
rect 19152 4864 19216 4868
rect 19232 4924 19296 4928
rect 19232 4868 19236 4924
rect 19236 4868 19292 4924
rect 19292 4868 19296 4924
rect 19232 4864 19296 4868
rect 26912 4924 26976 4928
rect 26912 4868 26916 4924
rect 26916 4868 26972 4924
rect 26972 4868 26976 4924
rect 26912 4864 26976 4868
rect 26992 4924 27056 4928
rect 26992 4868 26996 4924
rect 26996 4868 27052 4924
rect 27052 4868 27056 4924
rect 26992 4864 27056 4868
rect 27072 4924 27136 4928
rect 27072 4868 27076 4924
rect 27076 4868 27132 4924
rect 27132 4868 27136 4924
rect 27072 4864 27136 4868
rect 27152 4924 27216 4928
rect 27152 4868 27156 4924
rect 27156 4868 27212 4924
rect 27212 4868 27216 4924
rect 27152 4864 27216 4868
rect 27232 4924 27296 4928
rect 27232 4868 27236 4924
rect 27236 4868 27292 4924
rect 27292 4868 27296 4924
rect 27232 4864 27296 4868
rect 3652 4380 3716 4384
rect 3652 4324 3656 4380
rect 3656 4324 3712 4380
rect 3712 4324 3716 4380
rect 3652 4320 3716 4324
rect 3732 4380 3796 4384
rect 3732 4324 3736 4380
rect 3736 4324 3792 4380
rect 3792 4324 3796 4380
rect 3732 4320 3796 4324
rect 3812 4380 3876 4384
rect 3812 4324 3816 4380
rect 3816 4324 3872 4380
rect 3872 4324 3876 4380
rect 3812 4320 3876 4324
rect 3892 4380 3956 4384
rect 3892 4324 3896 4380
rect 3896 4324 3952 4380
rect 3952 4324 3956 4380
rect 3892 4320 3956 4324
rect 3972 4380 4036 4384
rect 3972 4324 3976 4380
rect 3976 4324 4032 4380
rect 4032 4324 4036 4380
rect 3972 4320 4036 4324
rect 11652 4380 11716 4384
rect 11652 4324 11656 4380
rect 11656 4324 11712 4380
rect 11712 4324 11716 4380
rect 11652 4320 11716 4324
rect 11732 4380 11796 4384
rect 11732 4324 11736 4380
rect 11736 4324 11792 4380
rect 11792 4324 11796 4380
rect 11732 4320 11796 4324
rect 11812 4380 11876 4384
rect 11812 4324 11816 4380
rect 11816 4324 11872 4380
rect 11872 4324 11876 4380
rect 11812 4320 11876 4324
rect 11892 4380 11956 4384
rect 11892 4324 11896 4380
rect 11896 4324 11952 4380
rect 11952 4324 11956 4380
rect 11892 4320 11956 4324
rect 11972 4380 12036 4384
rect 11972 4324 11976 4380
rect 11976 4324 12032 4380
rect 12032 4324 12036 4380
rect 11972 4320 12036 4324
rect 19652 4380 19716 4384
rect 19652 4324 19656 4380
rect 19656 4324 19712 4380
rect 19712 4324 19716 4380
rect 19652 4320 19716 4324
rect 19732 4380 19796 4384
rect 19732 4324 19736 4380
rect 19736 4324 19792 4380
rect 19792 4324 19796 4380
rect 19732 4320 19796 4324
rect 19812 4380 19876 4384
rect 19812 4324 19816 4380
rect 19816 4324 19872 4380
rect 19872 4324 19876 4380
rect 19812 4320 19876 4324
rect 19892 4380 19956 4384
rect 19892 4324 19896 4380
rect 19896 4324 19952 4380
rect 19952 4324 19956 4380
rect 19892 4320 19956 4324
rect 19972 4380 20036 4384
rect 19972 4324 19976 4380
rect 19976 4324 20032 4380
rect 20032 4324 20036 4380
rect 19972 4320 20036 4324
rect 27652 4380 27716 4384
rect 27652 4324 27656 4380
rect 27656 4324 27712 4380
rect 27712 4324 27716 4380
rect 27652 4320 27716 4324
rect 27732 4380 27796 4384
rect 27732 4324 27736 4380
rect 27736 4324 27792 4380
rect 27792 4324 27796 4380
rect 27732 4320 27796 4324
rect 27812 4380 27876 4384
rect 27812 4324 27816 4380
rect 27816 4324 27872 4380
rect 27872 4324 27876 4380
rect 27812 4320 27876 4324
rect 27892 4380 27956 4384
rect 27892 4324 27896 4380
rect 27896 4324 27952 4380
rect 27952 4324 27956 4380
rect 27892 4320 27956 4324
rect 27972 4380 28036 4384
rect 27972 4324 27976 4380
rect 27976 4324 28032 4380
rect 28032 4324 28036 4380
rect 27972 4320 28036 4324
rect 2912 3836 2976 3840
rect 2912 3780 2916 3836
rect 2916 3780 2972 3836
rect 2972 3780 2976 3836
rect 2912 3776 2976 3780
rect 2992 3836 3056 3840
rect 2992 3780 2996 3836
rect 2996 3780 3052 3836
rect 3052 3780 3056 3836
rect 2992 3776 3056 3780
rect 3072 3836 3136 3840
rect 3072 3780 3076 3836
rect 3076 3780 3132 3836
rect 3132 3780 3136 3836
rect 3072 3776 3136 3780
rect 3152 3836 3216 3840
rect 3152 3780 3156 3836
rect 3156 3780 3212 3836
rect 3212 3780 3216 3836
rect 3152 3776 3216 3780
rect 3232 3836 3296 3840
rect 3232 3780 3236 3836
rect 3236 3780 3292 3836
rect 3292 3780 3296 3836
rect 3232 3776 3296 3780
rect 10912 3836 10976 3840
rect 10912 3780 10916 3836
rect 10916 3780 10972 3836
rect 10972 3780 10976 3836
rect 10912 3776 10976 3780
rect 10992 3836 11056 3840
rect 10992 3780 10996 3836
rect 10996 3780 11052 3836
rect 11052 3780 11056 3836
rect 10992 3776 11056 3780
rect 11072 3836 11136 3840
rect 11072 3780 11076 3836
rect 11076 3780 11132 3836
rect 11132 3780 11136 3836
rect 11072 3776 11136 3780
rect 11152 3836 11216 3840
rect 11152 3780 11156 3836
rect 11156 3780 11212 3836
rect 11212 3780 11216 3836
rect 11152 3776 11216 3780
rect 11232 3836 11296 3840
rect 11232 3780 11236 3836
rect 11236 3780 11292 3836
rect 11292 3780 11296 3836
rect 11232 3776 11296 3780
rect 18912 3836 18976 3840
rect 18912 3780 18916 3836
rect 18916 3780 18972 3836
rect 18972 3780 18976 3836
rect 18912 3776 18976 3780
rect 18992 3836 19056 3840
rect 18992 3780 18996 3836
rect 18996 3780 19052 3836
rect 19052 3780 19056 3836
rect 18992 3776 19056 3780
rect 19072 3836 19136 3840
rect 19072 3780 19076 3836
rect 19076 3780 19132 3836
rect 19132 3780 19136 3836
rect 19072 3776 19136 3780
rect 19152 3836 19216 3840
rect 19152 3780 19156 3836
rect 19156 3780 19212 3836
rect 19212 3780 19216 3836
rect 19152 3776 19216 3780
rect 19232 3836 19296 3840
rect 19232 3780 19236 3836
rect 19236 3780 19292 3836
rect 19292 3780 19296 3836
rect 19232 3776 19296 3780
rect 26912 3836 26976 3840
rect 26912 3780 26916 3836
rect 26916 3780 26972 3836
rect 26972 3780 26976 3836
rect 26912 3776 26976 3780
rect 26992 3836 27056 3840
rect 26992 3780 26996 3836
rect 26996 3780 27052 3836
rect 27052 3780 27056 3836
rect 26992 3776 27056 3780
rect 27072 3836 27136 3840
rect 27072 3780 27076 3836
rect 27076 3780 27132 3836
rect 27132 3780 27136 3836
rect 27072 3776 27136 3780
rect 27152 3836 27216 3840
rect 27152 3780 27156 3836
rect 27156 3780 27212 3836
rect 27212 3780 27216 3836
rect 27152 3776 27216 3780
rect 27232 3836 27296 3840
rect 27232 3780 27236 3836
rect 27236 3780 27292 3836
rect 27292 3780 27296 3836
rect 27232 3776 27296 3780
rect 3652 3292 3716 3296
rect 3652 3236 3656 3292
rect 3656 3236 3712 3292
rect 3712 3236 3716 3292
rect 3652 3232 3716 3236
rect 3732 3292 3796 3296
rect 3732 3236 3736 3292
rect 3736 3236 3792 3292
rect 3792 3236 3796 3292
rect 3732 3232 3796 3236
rect 3812 3292 3876 3296
rect 3812 3236 3816 3292
rect 3816 3236 3872 3292
rect 3872 3236 3876 3292
rect 3812 3232 3876 3236
rect 3892 3292 3956 3296
rect 3892 3236 3896 3292
rect 3896 3236 3952 3292
rect 3952 3236 3956 3292
rect 3892 3232 3956 3236
rect 3972 3292 4036 3296
rect 3972 3236 3976 3292
rect 3976 3236 4032 3292
rect 4032 3236 4036 3292
rect 3972 3232 4036 3236
rect 11652 3292 11716 3296
rect 11652 3236 11656 3292
rect 11656 3236 11712 3292
rect 11712 3236 11716 3292
rect 11652 3232 11716 3236
rect 11732 3292 11796 3296
rect 11732 3236 11736 3292
rect 11736 3236 11792 3292
rect 11792 3236 11796 3292
rect 11732 3232 11796 3236
rect 11812 3292 11876 3296
rect 11812 3236 11816 3292
rect 11816 3236 11872 3292
rect 11872 3236 11876 3292
rect 11812 3232 11876 3236
rect 11892 3292 11956 3296
rect 11892 3236 11896 3292
rect 11896 3236 11952 3292
rect 11952 3236 11956 3292
rect 11892 3232 11956 3236
rect 11972 3292 12036 3296
rect 11972 3236 11976 3292
rect 11976 3236 12032 3292
rect 12032 3236 12036 3292
rect 11972 3232 12036 3236
rect 19652 3292 19716 3296
rect 19652 3236 19656 3292
rect 19656 3236 19712 3292
rect 19712 3236 19716 3292
rect 19652 3232 19716 3236
rect 19732 3292 19796 3296
rect 19732 3236 19736 3292
rect 19736 3236 19792 3292
rect 19792 3236 19796 3292
rect 19732 3232 19796 3236
rect 19812 3292 19876 3296
rect 19812 3236 19816 3292
rect 19816 3236 19872 3292
rect 19872 3236 19876 3292
rect 19812 3232 19876 3236
rect 19892 3292 19956 3296
rect 19892 3236 19896 3292
rect 19896 3236 19952 3292
rect 19952 3236 19956 3292
rect 19892 3232 19956 3236
rect 19972 3292 20036 3296
rect 19972 3236 19976 3292
rect 19976 3236 20032 3292
rect 20032 3236 20036 3292
rect 19972 3232 20036 3236
rect 27652 3292 27716 3296
rect 27652 3236 27656 3292
rect 27656 3236 27712 3292
rect 27712 3236 27716 3292
rect 27652 3232 27716 3236
rect 27732 3292 27796 3296
rect 27732 3236 27736 3292
rect 27736 3236 27792 3292
rect 27792 3236 27796 3292
rect 27732 3232 27796 3236
rect 27812 3292 27876 3296
rect 27812 3236 27816 3292
rect 27816 3236 27872 3292
rect 27872 3236 27876 3292
rect 27812 3232 27876 3236
rect 27892 3292 27956 3296
rect 27892 3236 27896 3292
rect 27896 3236 27952 3292
rect 27952 3236 27956 3292
rect 27892 3232 27956 3236
rect 27972 3292 28036 3296
rect 27972 3236 27976 3292
rect 27976 3236 28032 3292
rect 28032 3236 28036 3292
rect 27972 3232 28036 3236
rect 2912 2748 2976 2752
rect 2912 2692 2916 2748
rect 2916 2692 2972 2748
rect 2972 2692 2976 2748
rect 2912 2688 2976 2692
rect 2992 2748 3056 2752
rect 2992 2692 2996 2748
rect 2996 2692 3052 2748
rect 3052 2692 3056 2748
rect 2992 2688 3056 2692
rect 3072 2748 3136 2752
rect 3072 2692 3076 2748
rect 3076 2692 3132 2748
rect 3132 2692 3136 2748
rect 3072 2688 3136 2692
rect 3152 2748 3216 2752
rect 3152 2692 3156 2748
rect 3156 2692 3212 2748
rect 3212 2692 3216 2748
rect 3152 2688 3216 2692
rect 3232 2748 3296 2752
rect 3232 2692 3236 2748
rect 3236 2692 3292 2748
rect 3292 2692 3296 2748
rect 3232 2688 3296 2692
rect 10912 2748 10976 2752
rect 10912 2692 10916 2748
rect 10916 2692 10972 2748
rect 10972 2692 10976 2748
rect 10912 2688 10976 2692
rect 10992 2748 11056 2752
rect 10992 2692 10996 2748
rect 10996 2692 11052 2748
rect 11052 2692 11056 2748
rect 10992 2688 11056 2692
rect 11072 2748 11136 2752
rect 11072 2692 11076 2748
rect 11076 2692 11132 2748
rect 11132 2692 11136 2748
rect 11072 2688 11136 2692
rect 11152 2748 11216 2752
rect 11152 2692 11156 2748
rect 11156 2692 11212 2748
rect 11212 2692 11216 2748
rect 11152 2688 11216 2692
rect 11232 2748 11296 2752
rect 11232 2692 11236 2748
rect 11236 2692 11292 2748
rect 11292 2692 11296 2748
rect 11232 2688 11296 2692
rect 18912 2748 18976 2752
rect 18912 2692 18916 2748
rect 18916 2692 18972 2748
rect 18972 2692 18976 2748
rect 18912 2688 18976 2692
rect 18992 2748 19056 2752
rect 18992 2692 18996 2748
rect 18996 2692 19052 2748
rect 19052 2692 19056 2748
rect 18992 2688 19056 2692
rect 19072 2748 19136 2752
rect 19072 2692 19076 2748
rect 19076 2692 19132 2748
rect 19132 2692 19136 2748
rect 19072 2688 19136 2692
rect 19152 2748 19216 2752
rect 19152 2692 19156 2748
rect 19156 2692 19212 2748
rect 19212 2692 19216 2748
rect 19152 2688 19216 2692
rect 19232 2748 19296 2752
rect 19232 2692 19236 2748
rect 19236 2692 19292 2748
rect 19292 2692 19296 2748
rect 19232 2688 19296 2692
rect 26912 2748 26976 2752
rect 26912 2692 26916 2748
rect 26916 2692 26972 2748
rect 26972 2692 26976 2748
rect 26912 2688 26976 2692
rect 26992 2748 27056 2752
rect 26992 2692 26996 2748
rect 26996 2692 27052 2748
rect 27052 2692 27056 2748
rect 26992 2688 27056 2692
rect 27072 2748 27136 2752
rect 27072 2692 27076 2748
rect 27076 2692 27132 2748
rect 27132 2692 27136 2748
rect 27072 2688 27136 2692
rect 27152 2748 27216 2752
rect 27152 2692 27156 2748
rect 27156 2692 27212 2748
rect 27212 2692 27216 2748
rect 27152 2688 27216 2692
rect 27232 2748 27296 2752
rect 27232 2692 27236 2748
rect 27236 2692 27292 2748
rect 27292 2692 27296 2748
rect 27232 2688 27296 2692
rect 3652 2204 3716 2208
rect 3652 2148 3656 2204
rect 3656 2148 3712 2204
rect 3712 2148 3716 2204
rect 3652 2144 3716 2148
rect 3732 2204 3796 2208
rect 3732 2148 3736 2204
rect 3736 2148 3792 2204
rect 3792 2148 3796 2204
rect 3732 2144 3796 2148
rect 3812 2204 3876 2208
rect 3812 2148 3816 2204
rect 3816 2148 3872 2204
rect 3872 2148 3876 2204
rect 3812 2144 3876 2148
rect 3892 2204 3956 2208
rect 3892 2148 3896 2204
rect 3896 2148 3952 2204
rect 3952 2148 3956 2204
rect 3892 2144 3956 2148
rect 3972 2204 4036 2208
rect 3972 2148 3976 2204
rect 3976 2148 4032 2204
rect 4032 2148 4036 2204
rect 3972 2144 4036 2148
rect 11652 2204 11716 2208
rect 11652 2148 11656 2204
rect 11656 2148 11712 2204
rect 11712 2148 11716 2204
rect 11652 2144 11716 2148
rect 11732 2204 11796 2208
rect 11732 2148 11736 2204
rect 11736 2148 11792 2204
rect 11792 2148 11796 2204
rect 11732 2144 11796 2148
rect 11812 2204 11876 2208
rect 11812 2148 11816 2204
rect 11816 2148 11872 2204
rect 11872 2148 11876 2204
rect 11812 2144 11876 2148
rect 11892 2204 11956 2208
rect 11892 2148 11896 2204
rect 11896 2148 11952 2204
rect 11952 2148 11956 2204
rect 11892 2144 11956 2148
rect 11972 2204 12036 2208
rect 11972 2148 11976 2204
rect 11976 2148 12032 2204
rect 12032 2148 12036 2204
rect 11972 2144 12036 2148
rect 19652 2204 19716 2208
rect 19652 2148 19656 2204
rect 19656 2148 19712 2204
rect 19712 2148 19716 2204
rect 19652 2144 19716 2148
rect 19732 2204 19796 2208
rect 19732 2148 19736 2204
rect 19736 2148 19792 2204
rect 19792 2148 19796 2204
rect 19732 2144 19796 2148
rect 19812 2204 19876 2208
rect 19812 2148 19816 2204
rect 19816 2148 19872 2204
rect 19872 2148 19876 2204
rect 19812 2144 19876 2148
rect 19892 2204 19956 2208
rect 19892 2148 19896 2204
rect 19896 2148 19952 2204
rect 19952 2148 19956 2204
rect 19892 2144 19956 2148
rect 19972 2204 20036 2208
rect 19972 2148 19976 2204
rect 19976 2148 20032 2204
rect 20032 2148 20036 2204
rect 19972 2144 20036 2148
rect 27652 2204 27716 2208
rect 27652 2148 27656 2204
rect 27656 2148 27712 2204
rect 27712 2148 27716 2204
rect 27652 2144 27716 2148
rect 27732 2204 27796 2208
rect 27732 2148 27736 2204
rect 27736 2148 27792 2204
rect 27792 2148 27796 2204
rect 27732 2144 27796 2148
rect 27812 2204 27876 2208
rect 27812 2148 27816 2204
rect 27816 2148 27872 2204
rect 27872 2148 27876 2204
rect 27812 2144 27876 2148
rect 27892 2204 27956 2208
rect 27892 2148 27896 2204
rect 27896 2148 27952 2204
rect 27952 2148 27956 2204
rect 27892 2144 27956 2148
rect 27972 2204 28036 2208
rect 27972 2148 27976 2204
rect 27976 2148 28032 2204
rect 28032 2148 28036 2204
rect 27972 2144 28036 2148
<< metal4 >>
rect 2904 27776 3304 27792
rect 2904 27712 2912 27776
rect 2976 27712 2992 27776
rect 3056 27712 3072 27776
rect 3136 27712 3152 27776
rect 3216 27712 3232 27776
rect 3296 27712 3304 27776
rect 2904 26688 3304 27712
rect 2904 26624 2912 26688
rect 2976 26624 2992 26688
rect 3056 26624 3072 26688
rect 3136 26624 3152 26688
rect 3216 26624 3232 26688
rect 3296 26624 3304 26688
rect 2904 25600 3304 26624
rect 2904 25536 2912 25600
rect 2976 25536 2992 25600
rect 3056 25536 3072 25600
rect 3136 25536 3152 25600
rect 3216 25536 3232 25600
rect 3296 25536 3304 25600
rect 2904 24512 3304 25536
rect 2904 24448 2912 24512
rect 2976 24448 2992 24512
rect 3056 24448 3072 24512
rect 3136 24448 3152 24512
rect 3216 24448 3232 24512
rect 3296 24448 3304 24512
rect 2904 23424 3304 24448
rect 2904 23360 2912 23424
rect 2976 23360 2992 23424
rect 3056 23360 3072 23424
rect 3136 23360 3152 23424
rect 3216 23360 3232 23424
rect 3296 23360 3304 23424
rect 2904 22336 3304 23360
rect 2904 22272 2912 22336
rect 2976 22272 2992 22336
rect 3056 22272 3072 22336
rect 3136 22272 3152 22336
rect 3216 22272 3232 22336
rect 3296 22272 3304 22336
rect 1715 21316 1781 21317
rect 1715 21252 1716 21316
rect 1780 21252 1781 21316
rect 1715 21251 1781 21252
rect 1718 16285 1778 21251
rect 2904 21248 3304 22272
rect 3644 27232 4044 27792
rect 3644 27168 3652 27232
rect 3716 27168 3732 27232
rect 3796 27168 3812 27232
rect 3876 27168 3892 27232
rect 3956 27168 3972 27232
rect 4036 27168 4044 27232
rect 3644 26144 4044 27168
rect 3644 26080 3652 26144
rect 3716 26080 3732 26144
rect 3796 26080 3812 26144
rect 3876 26080 3892 26144
rect 3956 26080 3972 26144
rect 4036 26080 4044 26144
rect 3644 25056 4044 26080
rect 3644 24992 3652 25056
rect 3716 24992 3732 25056
rect 3796 24992 3812 25056
rect 3876 24992 3892 25056
rect 3956 24992 3972 25056
rect 4036 24992 4044 25056
rect 3644 23968 4044 24992
rect 3644 23904 3652 23968
rect 3716 23904 3732 23968
rect 3796 23904 3812 23968
rect 3876 23904 3892 23968
rect 3956 23904 3972 23968
rect 4036 23904 4044 23968
rect 3644 22880 4044 23904
rect 3644 22816 3652 22880
rect 3716 22816 3732 22880
rect 3796 22816 3812 22880
rect 3876 22816 3892 22880
rect 3956 22816 3972 22880
rect 4036 22816 4044 22880
rect 3371 21996 3437 21997
rect 3371 21932 3372 21996
rect 3436 21932 3437 21996
rect 3371 21931 3437 21932
rect 2904 21184 2912 21248
rect 2976 21184 2992 21248
rect 3056 21184 3072 21248
rect 3136 21184 3152 21248
rect 3216 21184 3232 21248
rect 3296 21184 3304 21248
rect 2635 20772 2701 20773
rect 2635 20708 2636 20772
rect 2700 20708 2701 20772
rect 2635 20707 2701 20708
rect 2083 19412 2149 19413
rect 2083 19348 2084 19412
rect 2148 19348 2149 19412
rect 2083 19347 2149 19348
rect 1715 16284 1781 16285
rect 1715 16220 1716 16284
rect 1780 16220 1781 16284
rect 1715 16219 1781 16220
rect 2086 12069 2146 19347
rect 2638 16557 2698 20707
rect 2904 20160 3304 21184
rect 2904 20096 2912 20160
rect 2976 20096 2992 20160
rect 3056 20096 3072 20160
rect 3136 20096 3152 20160
rect 3216 20096 3232 20160
rect 3296 20096 3304 20160
rect 2904 19072 3304 20096
rect 3374 19413 3434 21931
rect 3644 21792 4044 22816
rect 3644 21728 3652 21792
rect 3716 21728 3732 21792
rect 3796 21728 3812 21792
rect 3876 21728 3892 21792
rect 3956 21728 3972 21792
rect 4036 21728 4044 21792
rect 3644 20704 4044 21728
rect 3644 20640 3652 20704
rect 3716 20640 3732 20704
rect 3796 20640 3812 20704
rect 3876 20640 3892 20704
rect 3956 20640 3972 20704
rect 4036 20640 4044 20704
rect 3644 19616 4044 20640
rect 3644 19552 3652 19616
rect 3716 19552 3732 19616
rect 3796 19552 3812 19616
rect 3876 19552 3892 19616
rect 3956 19552 3972 19616
rect 4036 19552 4044 19616
rect 3371 19412 3437 19413
rect 3371 19348 3372 19412
rect 3436 19348 3437 19412
rect 3371 19347 3437 19348
rect 2904 19008 2912 19072
rect 2976 19008 2992 19072
rect 3056 19008 3072 19072
rect 3136 19008 3152 19072
rect 3216 19008 3232 19072
rect 3296 19008 3304 19072
rect 2904 17984 3304 19008
rect 2904 17920 2912 17984
rect 2976 17920 2992 17984
rect 3056 17920 3072 17984
rect 3136 17920 3152 17984
rect 3216 17920 3232 17984
rect 3296 17920 3304 17984
rect 2904 16896 3304 17920
rect 3644 18528 4044 19552
rect 3644 18464 3652 18528
rect 3716 18464 3732 18528
rect 3796 18464 3812 18528
rect 3876 18464 3892 18528
rect 3956 18464 3972 18528
rect 4036 18464 4044 18528
rect 3644 17440 4044 18464
rect 3644 17376 3652 17440
rect 3716 17376 3732 17440
rect 3796 17376 3812 17440
rect 3876 17376 3892 17440
rect 3956 17376 3972 17440
rect 4036 17376 4044 17440
rect 3371 17100 3437 17101
rect 3371 17036 3372 17100
rect 3436 17036 3437 17100
rect 3371 17035 3437 17036
rect 2904 16832 2912 16896
rect 2976 16832 2992 16896
rect 3056 16832 3072 16896
rect 3136 16832 3152 16896
rect 3216 16832 3232 16896
rect 3296 16832 3304 16896
rect 2635 16556 2701 16557
rect 2635 16492 2636 16556
rect 2700 16492 2701 16556
rect 2635 16491 2701 16492
rect 2638 15061 2698 16491
rect 2904 15808 3304 16832
rect 2904 15744 2912 15808
rect 2976 15744 2992 15808
rect 3056 15744 3072 15808
rect 3136 15744 3152 15808
rect 3216 15744 3232 15808
rect 3296 15744 3304 15808
rect 2635 15060 2701 15061
rect 2635 14996 2636 15060
rect 2700 14996 2701 15060
rect 2635 14995 2701 14996
rect 2904 14720 3304 15744
rect 2904 14656 2912 14720
rect 2976 14656 2992 14720
rect 3056 14656 3072 14720
rect 3136 14656 3152 14720
rect 3216 14656 3232 14720
rect 3296 14656 3304 14720
rect 2904 13632 3304 14656
rect 2904 13568 2912 13632
rect 2976 13568 2992 13632
rect 3056 13568 3072 13632
rect 3136 13568 3152 13632
rect 3216 13568 3232 13632
rect 3296 13568 3304 13632
rect 2904 12544 3304 13568
rect 2904 12480 2912 12544
rect 2976 12480 2992 12544
rect 3056 12480 3072 12544
rect 3136 12480 3152 12544
rect 3216 12480 3232 12544
rect 3296 12480 3304 12544
rect 2083 12068 2149 12069
rect 2083 12004 2084 12068
rect 2148 12004 2149 12068
rect 2083 12003 2149 12004
rect 2904 11456 3304 12480
rect 2904 11392 2912 11456
rect 2976 11392 2992 11456
rect 3056 11392 3072 11456
rect 3136 11392 3152 11456
rect 3216 11392 3232 11456
rect 3296 11392 3304 11456
rect 2904 10368 3304 11392
rect 3374 11389 3434 17035
rect 3644 16352 4044 17376
rect 3644 16288 3652 16352
rect 3716 16288 3732 16352
rect 3796 16288 3812 16352
rect 3876 16288 3892 16352
rect 3956 16288 3972 16352
rect 4036 16288 4044 16352
rect 3644 15264 4044 16288
rect 3644 15200 3652 15264
rect 3716 15200 3732 15264
rect 3796 15200 3812 15264
rect 3876 15200 3892 15264
rect 3956 15200 3972 15264
rect 4036 15200 4044 15264
rect 3644 14176 4044 15200
rect 3644 14112 3652 14176
rect 3716 14112 3732 14176
rect 3796 14112 3812 14176
rect 3876 14112 3892 14176
rect 3956 14112 3972 14176
rect 4036 14112 4044 14176
rect 3644 13088 4044 14112
rect 3644 13024 3652 13088
rect 3716 13024 3732 13088
rect 3796 13024 3812 13088
rect 3876 13024 3892 13088
rect 3956 13024 3972 13088
rect 4036 13024 4044 13088
rect 3644 12000 4044 13024
rect 3644 11936 3652 12000
rect 3716 11936 3732 12000
rect 3796 11936 3812 12000
rect 3876 11936 3892 12000
rect 3956 11936 3972 12000
rect 4036 11936 4044 12000
rect 3371 11388 3437 11389
rect 3371 11324 3372 11388
rect 3436 11324 3437 11388
rect 3371 11323 3437 11324
rect 2904 10304 2912 10368
rect 2976 10304 2992 10368
rect 3056 10304 3072 10368
rect 3136 10304 3152 10368
rect 3216 10304 3232 10368
rect 3296 10304 3304 10368
rect 2904 9280 3304 10304
rect 2904 9216 2912 9280
rect 2976 9216 2992 9280
rect 3056 9216 3072 9280
rect 3136 9216 3152 9280
rect 3216 9216 3232 9280
rect 3296 9216 3304 9280
rect 2904 8192 3304 9216
rect 2904 8128 2912 8192
rect 2976 8128 2992 8192
rect 3056 8128 3072 8192
rect 3136 8128 3152 8192
rect 3216 8128 3232 8192
rect 3296 8128 3304 8192
rect 2904 7104 3304 8128
rect 2904 7040 2912 7104
rect 2976 7040 2992 7104
rect 3056 7040 3072 7104
rect 3136 7040 3152 7104
rect 3216 7040 3232 7104
rect 3296 7040 3304 7104
rect 2904 6016 3304 7040
rect 2904 5952 2912 6016
rect 2976 5952 2992 6016
rect 3056 5952 3072 6016
rect 3136 5952 3152 6016
rect 3216 5952 3232 6016
rect 3296 5952 3304 6016
rect 2904 4928 3304 5952
rect 2904 4864 2912 4928
rect 2976 4864 2992 4928
rect 3056 4864 3072 4928
rect 3136 4864 3152 4928
rect 3216 4864 3232 4928
rect 3296 4864 3304 4928
rect 2904 3840 3304 4864
rect 2904 3776 2912 3840
rect 2976 3776 2992 3840
rect 3056 3776 3072 3840
rect 3136 3776 3152 3840
rect 3216 3776 3232 3840
rect 3296 3776 3304 3840
rect 2904 2752 3304 3776
rect 2904 2688 2912 2752
rect 2976 2688 2992 2752
rect 3056 2688 3072 2752
rect 3136 2688 3152 2752
rect 3216 2688 3232 2752
rect 3296 2688 3304 2752
rect 2904 2128 3304 2688
rect 3644 10912 4044 11936
rect 3644 10848 3652 10912
rect 3716 10848 3732 10912
rect 3796 10848 3812 10912
rect 3876 10848 3892 10912
rect 3956 10848 3972 10912
rect 4036 10848 4044 10912
rect 3644 9824 4044 10848
rect 3644 9760 3652 9824
rect 3716 9760 3732 9824
rect 3796 9760 3812 9824
rect 3876 9760 3892 9824
rect 3956 9760 3972 9824
rect 4036 9760 4044 9824
rect 3644 8736 4044 9760
rect 3644 8672 3652 8736
rect 3716 8672 3732 8736
rect 3796 8672 3812 8736
rect 3876 8672 3892 8736
rect 3956 8672 3972 8736
rect 4036 8672 4044 8736
rect 3644 7648 4044 8672
rect 3644 7584 3652 7648
rect 3716 7584 3732 7648
rect 3796 7584 3812 7648
rect 3876 7584 3892 7648
rect 3956 7584 3972 7648
rect 4036 7584 4044 7648
rect 3644 6560 4044 7584
rect 3644 6496 3652 6560
rect 3716 6496 3732 6560
rect 3796 6496 3812 6560
rect 3876 6496 3892 6560
rect 3956 6496 3972 6560
rect 4036 6496 4044 6560
rect 3644 5472 4044 6496
rect 3644 5408 3652 5472
rect 3716 5408 3732 5472
rect 3796 5408 3812 5472
rect 3876 5408 3892 5472
rect 3956 5408 3972 5472
rect 4036 5408 4044 5472
rect 3644 4384 4044 5408
rect 3644 4320 3652 4384
rect 3716 4320 3732 4384
rect 3796 4320 3812 4384
rect 3876 4320 3892 4384
rect 3956 4320 3972 4384
rect 4036 4320 4044 4384
rect 3644 3296 4044 4320
rect 3644 3232 3652 3296
rect 3716 3232 3732 3296
rect 3796 3232 3812 3296
rect 3876 3232 3892 3296
rect 3956 3232 3972 3296
rect 4036 3232 4044 3296
rect 3644 2208 4044 3232
rect 3644 2144 3652 2208
rect 3716 2144 3732 2208
rect 3796 2144 3812 2208
rect 3876 2144 3892 2208
rect 3956 2144 3972 2208
rect 4036 2144 4044 2208
rect 3644 2128 4044 2144
rect 10904 27776 11304 27792
rect 10904 27712 10912 27776
rect 10976 27712 10992 27776
rect 11056 27712 11072 27776
rect 11136 27712 11152 27776
rect 11216 27712 11232 27776
rect 11296 27712 11304 27776
rect 10904 26688 11304 27712
rect 10904 26624 10912 26688
rect 10976 26624 10992 26688
rect 11056 26624 11072 26688
rect 11136 26624 11152 26688
rect 11216 26624 11232 26688
rect 11296 26624 11304 26688
rect 10904 25600 11304 26624
rect 10904 25536 10912 25600
rect 10976 25536 10992 25600
rect 11056 25536 11072 25600
rect 11136 25536 11152 25600
rect 11216 25536 11232 25600
rect 11296 25536 11304 25600
rect 10904 24512 11304 25536
rect 10904 24448 10912 24512
rect 10976 24448 10992 24512
rect 11056 24448 11072 24512
rect 11136 24448 11152 24512
rect 11216 24448 11232 24512
rect 11296 24448 11304 24512
rect 10904 23424 11304 24448
rect 10904 23360 10912 23424
rect 10976 23360 10992 23424
rect 11056 23360 11072 23424
rect 11136 23360 11152 23424
rect 11216 23360 11232 23424
rect 11296 23360 11304 23424
rect 10904 22336 11304 23360
rect 10904 22272 10912 22336
rect 10976 22272 10992 22336
rect 11056 22272 11072 22336
rect 11136 22272 11152 22336
rect 11216 22272 11232 22336
rect 11296 22272 11304 22336
rect 10904 21248 11304 22272
rect 10904 21184 10912 21248
rect 10976 21184 10992 21248
rect 11056 21184 11072 21248
rect 11136 21184 11152 21248
rect 11216 21184 11232 21248
rect 11296 21184 11304 21248
rect 10904 20160 11304 21184
rect 10904 20096 10912 20160
rect 10976 20096 10992 20160
rect 11056 20096 11072 20160
rect 11136 20096 11152 20160
rect 11216 20096 11232 20160
rect 11296 20096 11304 20160
rect 10904 19072 11304 20096
rect 10904 19008 10912 19072
rect 10976 19008 10992 19072
rect 11056 19008 11072 19072
rect 11136 19008 11152 19072
rect 11216 19008 11232 19072
rect 11296 19008 11304 19072
rect 10904 17984 11304 19008
rect 10904 17920 10912 17984
rect 10976 17920 10992 17984
rect 11056 17920 11072 17984
rect 11136 17920 11152 17984
rect 11216 17920 11232 17984
rect 11296 17920 11304 17984
rect 10904 16896 11304 17920
rect 10904 16832 10912 16896
rect 10976 16832 10992 16896
rect 11056 16832 11072 16896
rect 11136 16832 11152 16896
rect 11216 16832 11232 16896
rect 11296 16832 11304 16896
rect 10904 15808 11304 16832
rect 10904 15744 10912 15808
rect 10976 15744 10992 15808
rect 11056 15744 11072 15808
rect 11136 15744 11152 15808
rect 11216 15744 11232 15808
rect 11296 15744 11304 15808
rect 10904 14720 11304 15744
rect 10904 14656 10912 14720
rect 10976 14656 10992 14720
rect 11056 14656 11072 14720
rect 11136 14656 11152 14720
rect 11216 14656 11232 14720
rect 11296 14656 11304 14720
rect 10904 13632 11304 14656
rect 10904 13568 10912 13632
rect 10976 13568 10992 13632
rect 11056 13568 11072 13632
rect 11136 13568 11152 13632
rect 11216 13568 11232 13632
rect 11296 13568 11304 13632
rect 10904 12544 11304 13568
rect 10904 12480 10912 12544
rect 10976 12480 10992 12544
rect 11056 12480 11072 12544
rect 11136 12480 11152 12544
rect 11216 12480 11232 12544
rect 11296 12480 11304 12544
rect 10904 11456 11304 12480
rect 10904 11392 10912 11456
rect 10976 11392 10992 11456
rect 11056 11392 11072 11456
rect 11136 11392 11152 11456
rect 11216 11392 11232 11456
rect 11296 11392 11304 11456
rect 10904 10368 11304 11392
rect 10904 10304 10912 10368
rect 10976 10304 10992 10368
rect 11056 10304 11072 10368
rect 11136 10304 11152 10368
rect 11216 10304 11232 10368
rect 11296 10304 11304 10368
rect 10904 9280 11304 10304
rect 10904 9216 10912 9280
rect 10976 9216 10992 9280
rect 11056 9216 11072 9280
rect 11136 9216 11152 9280
rect 11216 9216 11232 9280
rect 11296 9216 11304 9280
rect 10904 8192 11304 9216
rect 10904 8128 10912 8192
rect 10976 8128 10992 8192
rect 11056 8128 11072 8192
rect 11136 8128 11152 8192
rect 11216 8128 11232 8192
rect 11296 8128 11304 8192
rect 10904 7104 11304 8128
rect 10904 7040 10912 7104
rect 10976 7040 10992 7104
rect 11056 7040 11072 7104
rect 11136 7040 11152 7104
rect 11216 7040 11232 7104
rect 11296 7040 11304 7104
rect 10904 6016 11304 7040
rect 10904 5952 10912 6016
rect 10976 5952 10992 6016
rect 11056 5952 11072 6016
rect 11136 5952 11152 6016
rect 11216 5952 11232 6016
rect 11296 5952 11304 6016
rect 10904 4928 11304 5952
rect 10904 4864 10912 4928
rect 10976 4864 10992 4928
rect 11056 4864 11072 4928
rect 11136 4864 11152 4928
rect 11216 4864 11232 4928
rect 11296 4864 11304 4928
rect 10904 3840 11304 4864
rect 10904 3776 10912 3840
rect 10976 3776 10992 3840
rect 11056 3776 11072 3840
rect 11136 3776 11152 3840
rect 11216 3776 11232 3840
rect 11296 3776 11304 3840
rect 10904 2752 11304 3776
rect 10904 2688 10912 2752
rect 10976 2688 10992 2752
rect 11056 2688 11072 2752
rect 11136 2688 11152 2752
rect 11216 2688 11232 2752
rect 11296 2688 11304 2752
rect 10904 2128 11304 2688
rect 11644 27232 12044 27792
rect 11644 27168 11652 27232
rect 11716 27168 11732 27232
rect 11796 27168 11812 27232
rect 11876 27168 11892 27232
rect 11956 27168 11972 27232
rect 12036 27168 12044 27232
rect 11644 26144 12044 27168
rect 11644 26080 11652 26144
rect 11716 26080 11732 26144
rect 11796 26080 11812 26144
rect 11876 26080 11892 26144
rect 11956 26080 11972 26144
rect 12036 26080 12044 26144
rect 11644 25056 12044 26080
rect 11644 24992 11652 25056
rect 11716 24992 11732 25056
rect 11796 24992 11812 25056
rect 11876 24992 11892 25056
rect 11956 24992 11972 25056
rect 12036 24992 12044 25056
rect 11644 23968 12044 24992
rect 11644 23904 11652 23968
rect 11716 23904 11732 23968
rect 11796 23904 11812 23968
rect 11876 23904 11892 23968
rect 11956 23904 11972 23968
rect 12036 23904 12044 23968
rect 11644 22880 12044 23904
rect 11644 22816 11652 22880
rect 11716 22816 11732 22880
rect 11796 22816 11812 22880
rect 11876 22816 11892 22880
rect 11956 22816 11972 22880
rect 12036 22816 12044 22880
rect 11644 21792 12044 22816
rect 11644 21728 11652 21792
rect 11716 21728 11732 21792
rect 11796 21728 11812 21792
rect 11876 21728 11892 21792
rect 11956 21728 11972 21792
rect 12036 21728 12044 21792
rect 11644 20704 12044 21728
rect 11644 20640 11652 20704
rect 11716 20640 11732 20704
rect 11796 20640 11812 20704
rect 11876 20640 11892 20704
rect 11956 20640 11972 20704
rect 12036 20640 12044 20704
rect 11644 19616 12044 20640
rect 11644 19552 11652 19616
rect 11716 19552 11732 19616
rect 11796 19552 11812 19616
rect 11876 19552 11892 19616
rect 11956 19552 11972 19616
rect 12036 19552 12044 19616
rect 11644 18528 12044 19552
rect 11644 18464 11652 18528
rect 11716 18464 11732 18528
rect 11796 18464 11812 18528
rect 11876 18464 11892 18528
rect 11956 18464 11972 18528
rect 12036 18464 12044 18528
rect 11644 17440 12044 18464
rect 11644 17376 11652 17440
rect 11716 17376 11732 17440
rect 11796 17376 11812 17440
rect 11876 17376 11892 17440
rect 11956 17376 11972 17440
rect 12036 17376 12044 17440
rect 11644 16352 12044 17376
rect 11644 16288 11652 16352
rect 11716 16288 11732 16352
rect 11796 16288 11812 16352
rect 11876 16288 11892 16352
rect 11956 16288 11972 16352
rect 12036 16288 12044 16352
rect 11644 15264 12044 16288
rect 11644 15200 11652 15264
rect 11716 15200 11732 15264
rect 11796 15200 11812 15264
rect 11876 15200 11892 15264
rect 11956 15200 11972 15264
rect 12036 15200 12044 15264
rect 11644 14176 12044 15200
rect 11644 14112 11652 14176
rect 11716 14112 11732 14176
rect 11796 14112 11812 14176
rect 11876 14112 11892 14176
rect 11956 14112 11972 14176
rect 12036 14112 12044 14176
rect 11644 13088 12044 14112
rect 11644 13024 11652 13088
rect 11716 13024 11732 13088
rect 11796 13024 11812 13088
rect 11876 13024 11892 13088
rect 11956 13024 11972 13088
rect 12036 13024 12044 13088
rect 11644 12000 12044 13024
rect 11644 11936 11652 12000
rect 11716 11936 11732 12000
rect 11796 11936 11812 12000
rect 11876 11936 11892 12000
rect 11956 11936 11972 12000
rect 12036 11936 12044 12000
rect 11644 10912 12044 11936
rect 11644 10848 11652 10912
rect 11716 10848 11732 10912
rect 11796 10848 11812 10912
rect 11876 10848 11892 10912
rect 11956 10848 11972 10912
rect 12036 10848 12044 10912
rect 11644 9824 12044 10848
rect 11644 9760 11652 9824
rect 11716 9760 11732 9824
rect 11796 9760 11812 9824
rect 11876 9760 11892 9824
rect 11956 9760 11972 9824
rect 12036 9760 12044 9824
rect 11644 8736 12044 9760
rect 11644 8672 11652 8736
rect 11716 8672 11732 8736
rect 11796 8672 11812 8736
rect 11876 8672 11892 8736
rect 11956 8672 11972 8736
rect 12036 8672 12044 8736
rect 11644 7648 12044 8672
rect 11644 7584 11652 7648
rect 11716 7584 11732 7648
rect 11796 7584 11812 7648
rect 11876 7584 11892 7648
rect 11956 7584 11972 7648
rect 12036 7584 12044 7648
rect 11644 6560 12044 7584
rect 11644 6496 11652 6560
rect 11716 6496 11732 6560
rect 11796 6496 11812 6560
rect 11876 6496 11892 6560
rect 11956 6496 11972 6560
rect 12036 6496 12044 6560
rect 11644 5472 12044 6496
rect 11644 5408 11652 5472
rect 11716 5408 11732 5472
rect 11796 5408 11812 5472
rect 11876 5408 11892 5472
rect 11956 5408 11972 5472
rect 12036 5408 12044 5472
rect 11644 4384 12044 5408
rect 11644 4320 11652 4384
rect 11716 4320 11732 4384
rect 11796 4320 11812 4384
rect 11876 4320 11892 4384
rect 11956 4320 11972 4384
rect 12036 4320 12044 4384
rect 11644 3296 12044 4320
rect 11644 3232 11652 3296
rect 11716 3232 11732 3296
rect 11796 3232 11812 3296
rect 11876 3232 11892 3296
rect 11956 3232 11972 3296
rect 12036 3232 12044 3296
rect 11644 2208 12044 3232
rect 11644 2144 11652 2208
rect 11716 2144 11732 2208
rect 11796 2144 11812 2208
rect 11876 2144 11892 2208
rect 11956 2144 11972 2208
rect 12036 2144 12044 2208
rect 11644 2128 12044 2144
rect 18904 27776 19304 27792
rect 18904 27712 18912 27776
rect 18976 27712 18992 27776
rect 19056 27712 19072 27776
rect 19136 27712 19152 27776
rect 19216 27712 19232 27776
rect 19296 27712 19304 27776
rect 18904 26688 19304 27712
rect 18904 26624 18912 26688
rect 18976 26624 18992 26688
rect 19056 26624 19072 26688
rect 19136 26624 19152 26688
rect 19216 26624 19232 26688
rect 19296 26624 19304 26688
rect 18904 25600 19304 26624
rect 18904 25536 18912 25600
rect 18976 25536 18992 25600
rect 19056 25536 19072 25600
rect 19136 25536 19152 25600
rect 19216 25536 19232 25600
rect 19296 25536 19304 25600
rect 18904 24512 19304 25536
rect 18904 24448 18912 24512
rect 18976 24448 18992 24512
rect 19056 24448 19072 24512
rect 19136 24448 19152 24512
rect 19216 24448 19232 24512
rect 19296 24448 19304 24512
rect 18904 23424 19304 24448
rect 18904 23360 18912 23424
rect 18976 23360 18992 23424
rect 19056 23360 19072 23424
rect 19136 23360 19152 23424
rect 19216 23360 19232 23424
rect 19296 23360 19304 23424
rect 18904 22336 19304 23360
rect 18904 22272 18912 22336
rect 18976 22272 18992 22336
rect 19056 22272 19072 22336
rect 19136 22272 19152 22336
rect 19216 22272 19232 22336
rect 19296 22272 19304 22336
rect 18904 21248 19304 22272
rect 18904 21184 18912 21248
rect 18976 21184 18992 21248
rect 19056 21184 19072 21248
rect 19136 21184 19152 21248
rect 19216 21184 19232 21248
rect 19296 21184 19304 21248
rect 18904 20160 19304 21184
rect 18904 20096 18912 20160
rect 18976 20096 18992 20160
rect 19056 20096 19072 20160
rect 19136 20096 19152 20160
rect 19216 20096 19232 20160
rect 19296 20096 19304 20160
rect 18904 19072 19304 20096
rect 18904 19008 18912 19072
rect 18976 19008 18992 19072
rect 19056 19008 19072 19072
rect 19136 19008 19152 19072
rect 19216 19008 19232 19072
rect 19296 19008 19304 19072
rect 18904 17984 19304 19008
rect 18904 17920 18912 17984
rect 18976 17920 18992 17984
rect 19056 17920 19072 17984
rect 19136 17920 19152 17984
rect 19216 17920 19232 17984
rect 19296 17920 19304 17984
rect 18904 16896 19304 17920
rect 18904 16832 18912 16896
rect 18976 16832 18992 16896
rect 19056 16832 19072 16896
rect 19136 16832 19152 16896
rect 19216 16832 19232 16896
rect 19296 16832 19304 16896
rect 18904 15808 19304 16832
rect 18904 15744 18912 15808
rect 18976 15744 18992 15808
rect 19056 15744 19072 15808
rect 19136 15744 19152 15808
rect 19216 15744 19232 15808
rect 19296 15744 19304 15808
rect 18904 14720 19304 15744
rect 18904 14656 18912 14720
rect 18976 14656 18992 14720
rect 19056 14656 19072 14720
rect 19136 14656 19152 14720
rect 19216 14656 19232 14720
rect 19296 14656 19304 14720
rect 18904 13632 19304 14656
rect 18904 13568 18912 13632
rect 18976 13568 18992 13632
rect 19056 13568 19072 13632
rect 19136 13568 19152 13632
rect 19216 13568 19232 13632
rect 19296 13568 19304 13632
rect 18904 12544 19304 13568
rect 18904 12480 18912 12544
rect 18976 12480 18992 12544
rect 19056 12480 19072 12544
rect 19136 12480 19152 12544
rect 19216 12480 19232 12544
rect 19296 12480 19304 12544
rect 18904 11456 19304 12480
rect 18904 11392 18912 11456
rect 18976 11392 18992 11456
rect 19056 11392 19072 11456
rect 19136 11392 19152 11456
rect 19216 11392 19232 11456
rect 19296 11392 19304 11456
rect 18904 10368 19304 11392
rect 18904 10304 18912 10368
rect 18976 10304 18992 10368
rect 19056 10304 19072 10368
rect 19136 10304 19152 10368
rect 19216 10304 19232 10368
rect 19296 10304 19304 10368
rect 18904 9280 19304 10304
rect 18904 9216 18912 9280
rect 18976 9216 18992 9280
rect 19056 9216 19072 9280
rect 19136 9216 19152 9280
rect 19216 9216 19232 9280
rect 19296 9216 19304 9280
rect 18904 8192 19304 9216
rect 18904 8128 18912 8192
rect 18976 8128 18992 8192
rect 19056 8128 19072 8192
rect 19136 8128 19152 8192
rect 19216 8128 19232 8192
rect 19296 8128 19304 8192
rect 18904 7104 19304 8128
rect 18904 7040 18912 7104
rect 18976 7040 18992 7104
rect 19056 7040 19072 7104
rect 19136 7040 19152 7104
rect 19216 7040 19232 7104
rect 19296 7040 19304 7104
rect 18904 6016 19304 7040
rect 18904 5952 18912 6016
rect 18976 5952 18992 6016
rect 19056 5952 19072 6016
rect 19136 5952 19152 6016
rect 19216 5952 19232 6016
rect 19296 5952 19304 6016
rect 18904 4928 19304 5952
rect 18904 4864 18912 4928
rect 18976 4864 18992 4928
rect 19056 4864 19072 4928
rect 19136 4864 19152 4928
rect 19216 4864 19232 4928
rect 19296 4864 19304 4928
rect 18904 3840 19304 4864
rect 18904 3776 18912 3840
rect 18976 3776 18992 3840
rect 19056 3776 19072 3840
rect 19136 3776 19152 3840
rect 19216 3776 19232 3840
rect 19296 3776 19304 3840
rect 18904 2752 19304 3776
rect 18904 2688 18912 2752
rect 18976 2688 18992 2752
rect 19056 2688 19072 2752
rect 19136 2688 19152 2752
rect 19216 2688 19232 2752
rect 19296 2688 19304 2752
rect 18904 2128 19304 2688
rect 19644 27232 20044 27792
rect 19644 27168 19652 27232
rect 19716 27168 19732 27232
rect 19796 27168 19812 27232
rect 19876 27168 19892 27232
rect 19956 27168 19972 27232
rect 20036 27168 20044 27232
rect 19644 26144 20044 27168
rect 19644 26080 19652 26144
rect 19716 26080 19732 26144
rect 19796 26080 19812 26144
rect 19876 26080 19892 26144
rect 19956 26080 19972 26144
rect 20036 26080 20044 26144
rect 19644 25056 20044 26080
rect 19644 24992 19652 25056
rect 19716 24992 19732 25056
rect 19796 24992 19812 25056
rect 19876 24992 19892 25056
rect 19956 24992 19972 25056
rect 20036 24992 20044 25056
rect 19644 23968 20044 24992
rect 19644 23904 19652 23968
rect 19716 23904 19732 23968
rect 19796 23904 19812 23968
rect 19876 23904 19892 23968
rect 19956 23904 19972 23968
rect 20036 23904 20044 23968
rect 19644 22880 20044 23904
rect 19644 22816 19652 22880
rect 19716 22816 19732 22880
rect 19796 22816 19812 22880
rect 19876 22816 19892 22880
rect 19956 22816 19972 22880
rect 20036 22816 20044 22880
rect 19644 21792 20044 22816
rect 19644 21728 19652 21792
rect 19716 21728 19732 21792
rect 19796 21728 19812 21792
rect 19876 21728 19892 21792
rect 19956 21728 19972 21792
rect 20036 21728 20044 21792
rect 19644 20704 20044 21728
rect 19644 20640 19652 20704
rect 19716 20640 19732 20704
rect 19796 20640 19812 20704
rect 19876 20640 19892 20704
rect 19956 20640 19972 20704
rect 20036 20640 20044 20704
rect 19644 19616 20044 20640
rect 19644 19552 19652 19616
rect 19716 19552 19732 19616
rect 19796 19552 19812 19616
rect 19876 19552 19892 19616
rect 19956 19552 19972 19616
rect 20036 19552 20044 19616
rect 19644 18528 20044 19552
rect 19644 18464 19652 18528
rect 19716 18464 19732 18528
rect 19796 18464 19812 18528
rect 19876 18464 19892 18528
rect 19956 18464 19972 18528
rect 20036 18464 20044 18528
rect 19644 17440 20044 18464
rect 19644 17376 19652 17440
rect 19716 17376 19732 17440
rect 19796 17376 19812 17440
rect 19876 17376 19892 17440
rect 19956 17376 19972 17440
rect 20036 17376 20044 17440
rect 19644 16352 20044 17376
rect 19644 16288 19652 16352
rect 19716 16288 19732 16352
rect 19796 16288 19812 16352
rect 19876 16288 19892 16352
rect 19956 16288 19972 16352
rect 20036 16288 20044 16352
rect 19644 15264 20044 16288
rect 19644 15200 19652 15264
rect 19716 15200 19732 15264
rect 19796 15200 19812 15264
rect 19876 15200 19892 15264
rect 19956 15200 19972 15264
rect 20036 15200 20044 15264
rect 19644 14176 20044 15200
rect 19644 14112 19652 14176
rect 19716 14112 19732 14176
rect 19796 14112 19812 14176
rect 19876 14112 19892 14176
rect 19956 14112 19972 14176
rect 20036 14112 20044 14176
rect 19644 13088 20044 14112
rect 19644 13024 19652 13088
rect 19716 13024 19732 13088
rect 19796 13024 19812 13088
rect 19876 13024 19892 13088
rect 19956 13024 19972 13088
rect 20036 13024 20044 13088
rect 19644 12000 20044 13024
rect 19644 11936 19652 12000
rect 19716 11936 19732 12000
rect 19796 11936 19812 12000
rect 19876 11936 19892 12000
rect 19956 11936 19972 12000
rect 20036 11936 20044 12000
rect 19644 10912 20044 11936
rect 19644 10848 19652 10912
rect 19716 10848 19732 10912
rect 19796 10848 19812 10912
rect 19876 10848 19892 10912
rect 19956 10848 19972 10912
rect 20036 10848 20044 10912
rect 19644 9824 20044 10848
rect 19644 9760 19652 9824
rect 19716 9760 19732 9824
rect 19796 9760 19812 9824
rect 19876 9760 19892 9824
rect 19956 9760 19972 9824
rect 20036 9760 20044 9824
rect 19644 8736 20044 9760
rect 19644 8672 19652 8736
rect 19716 8672 19732 8736
rect 19796 8672 19812 8736
rect 19876 8672 19892 8736
rect 19956 8672 19972 8736
rect 20036 8672 20044 8736
rect 19644 7648 20044 8672
rect 19644 7584 19652 7648
rect 19716 7584 19732 7648
rect 19796 7584 19812 7648
rect 19876 7584 19892 7648
rect 19956 7584 19972 7648
rect 20036 7584 20044 7648
rect 19644 6560 20044 7584
rect 19644 6496 19652 6560
rect 19716 6496 19732 6560
rect 19796 6496 19812 6560
rect 19876 6496 19892 6560
rect 19956 6496 19972 6560
rect 20036 6496 20044 6560
rect 19644 5472 20044 6496
rect 19644 5408 19652 5472
rect 19716 5408 19732 5472
rect 19796 5408 19812 5472
rect 19876 5408 19892 5472
rect 19956 5408 19972 5472
rect 20036 5408 20044 5472
rect 19644 4384 20044 5408
rect 19644 4320 19652 4384
rect 19716 4320 19732 4384
rect 19796 4320 19812 4384
rect 19876 4320 19892 4384
rect 19956 4320 19972 4384
rect 20036 4320 20044 4384
rect 19644 3296 20044 4320
rect 19644 3232 19652 3296
rect 19716 3232 19732 3296
rect 19796 3232 19812 3296
rect 19876 3232 19892 3296
rect 19956 3232 19972 3296
rect 20036 3232 20044 3296
rect 19644 2208 20044 3232
rect 19644 2144 19652 2208
rect 19716 2144 19732 2208
rect 19796 2144 19812 2208
rect 19876 2144 19892 2208
rect 19956 2144 19972 2208
rect 20036 2144 20044 2208
rect 19644 2128 20044 2144
rect 26904 27776 27304 27792
rect 26904 27712 26912 27776
rect 26976 27712 26992 27776
rect 27056 27712 27072 27776
rect 27136 27712 27152 27776
rect 27216 27712 27232 27776
rect 27296 27712 27304 27776
rect 26904 26688 27304 27712
rect 26904 26624 26912 26688
rect 26976 26624 26992 26688
rect 27056 26624 27072 26688
rect 27136 26624 27152 26688
rect 27216 26624 27232 26688
rect 27296 26624 27304 26688
rect 26904 25600 27304 26624
rect 26904 25536 26912 25600
rect 26976 25536 26992 25600
rect 27056 25536 27072 25600
rect 27136 25536 27152 25600
rect 27216 25536 27232 25600
rect 27296 25536 27304 25600
rect 26904 24512 27304 25536
rect 26904 24448 26912 24512
rect 26976 24448 26992 24512
rect 27056 24448 27072 24512
rect 27136 24448 27152 24512
rect 27216 24448 27232 24512
rect 27296 24448 27304 24512
rect 26904 23424 27304 24448
rect 26904 23360 26912 23424
rect 26976 23360 26992 23424
rect 27056 23360 27072 23424
rect 27136 23360 27152 23424
rect 27216 23360 27232 23424
rect 27296 23360 27304 23424
rect 26904 22336 27304 23360
rect 26904 22272 26912 22336
rect 26976 22272 26992 22336
rect 27056 22272 27072 22336
rect 27136 22272 27152 22336
rect 27216 22272 27232 22336
rect 27296 22272 27304 22336
rect 26904 21248 27304 22272
rect 26904 21184 26912 21248
rect 26976 21184 26992 21248
rect 27056 21184 27072 21248
rect 27136 21184 27152 21248
rect 27216 21184 27232 21248
rect 27296 21184 27304 21248
rect 26904 20160 27304 21184
rect 26904 20096 26912 20160
rect 26976 20096 26992 20160
rect 27056 20096 27072 20160
rect 27136 20096 27152 20160
rect 27216 20096 27232 20160
rect 27296 20096 27304 20160
rect 26904 19072 27304 20096
rect 26904 19008 26912 19072
rect 26976 19008 26992 19072
rect 27056 19008 27072 19072
rect 27136 19008 27152 19072
rect 27216 19008 27232 19072
rect 27296 19008 27304 19072
rect 26904 17984 27304 19008
rect 26904 17920 26912 17984
rect 26976 17920 26992 17984
rect 27056 17920 27072 17984
rect 27136 17920 27152 17984
rect 27216 17920 27232 17984
rect 27296 17920 27304 17984
rect 26904 16896 27304 17920
rect 26904 16832 26912 16896
rect 26976 16832 26992 16896
rect 27056 16832 27072 16896
rect 27136 16832 27152 16896
rect 27216 16832 27232 16896
rect 27296 16832 27304 16896
rect 26904 15808 27304 16832
rect 26904 15744 26912 15808
rect 26976 15744 26992 15808
rect 27056 15744 27072 15808
rect 27136 15744 27152 15808
rect 27216 15744 27232 15808
rect 27296 15744 27304 15808
rect 26904 14720 27304 15744
rect 26904 14656 26912 14720
rect 26976 14656 26992 14720
rect 27056 14656 27072 14720
rect 27136 14656 27152 14720
rect 27216 14656 27232 14720
rect 27296 14656 27304 14720
rect 26904 13632 27304 14656
rect 26904 13568 26912 13632
rect 26976 13568 26992 13632
rect 27056 13568 27072 13632
rect 27136 13568 27152 13632
rect 27216 13568 27232 13632
rect 27296 13568 27304 13632
rect 26904 12544 27304 13568
rect 26904 12480 26912 12544
rect 26976 12480 26992 12544
rect 27056 12480 27072 12544
rect 27136 12480 27152 12544
rect 27216 12480 27232 12544
rect 27296 12480 27304 12544
rect 26904 11456 27304 12480
rect 26904 11392 26912 11456
rect 26976 11392 26992 11456
rect 27056 11392 27072 11456
rect 27136 11392 27152 11456
rect 27216 11392 27232 11456
rect 27296 11392 27304 11456
rect 26904 10368 27304 11392
rect 26904 10304 26912 10368
rect 26976 10304 26992 10368
rect 27056 10304 27072 10368
rect 27136 10304 27152 10368
rect 27216 10304 27232 10368
rect 27296 10304 27304 10368
rect 26904 9280 27304 10304
rect 26904 9216 26912 9280
rect 26976 9216 26992 9280
rect 27056 9216 27072 9280
rect 27136 9216 27152 9280
rect 27216 9216 27232 9280
rect 27296 9216 27304 9280
rect 26904 8192 27304 9216
rect 26904 8128 26912 8192
rect 26976 8128 26992 8192
rect 27056 8128 27072 8192
rect 27136 8128 27152 8192
rect 27216 8128 27232 8192
rect 27296 8128 27304 8192
rect 26904 7104 27304 8128
rect 26904 7040 26912 7104
rect 26976 7040 26992 7104
rect 27056 7040 27072 7104
rect 27136 7040 27152 7104
rect 27216 7040 27232 7104
rect 27296 7040 27304 7104
rect 26904 6016 27304 7040
rect 26904 5952 26912 6016
rect 26976 5952 26992 6016
rect 27056 5952 27072 6016
rect 27136 5952 27152 6016
rect 27216 5952 27232 6016
rect 27296 5952 27304 6016
rect 26904 4928 27304 5952
rect 26904 4864 26912 4928
rect 26976 4864 26992 4928
rect 27056 4864 27072 4928
rect 27136 4864 27152 4928
rect 27216 4864 27232 4928
rect 27296 4864 27304 4928
rect 26904 3840 27304 4864
rect 26904 3776 26912 3840
rect 26976 3776 26992 3840
rect 27056 3776 27072 3840
rect 27136 3776 27152 3840
rect 27216 3776 27232 3840
rect 27296 3776 27304 3840
rect 26904 2752 27304 3776
rect 26904 2688 26912 2752
rect 26976 2688 26992 2752
rect 27056 2688 27072 2752
rect 27136 2688 27152 2752
rect 27216 2688 27232 2752
rect 27296 2688 27304 2752
rect 26904 2128 27304 2688
rect 27644 27232 28044 27792
rect 27644 27168 27652 27232
rect 27716 27168 27732 27232
rect 27796 27168 27812 27232
rect 27876 27168 27892 27232
rect 27956 27168 27972 27232
rect 28036 27168 28044 27232
rect 27644 26144 28044 27168
rect 27644 26080 27652 26144
rect 27716 26080 27732 26144
rect 27796 26080 27812 26144
rect 27876 26080 27892 26144
rect 27956 26080 27972 26144
rect 28036 26080 28044 26144
rect 27644 25056 28044 26080
rect 27644 24992 27652 25056
rect 27716 24992 27732 25056
rect 27796 24992 27812 25056
rect 27876 24992 27892 25056
rect 27956 24992 27972 25056
rect 28036 24992 28044 25056
rect 27644 23968 28044 24992
rect 27644 23904 27652 23968
rect 27716 23904 27732 23968
rect 27796 23904 27812 23968
rect 27876 23904 27892 23968
rect 27956 23904 27972 23968
rect 28036 23904 28044 23968
rect 27644 22880 28044 23904
rect 27644 22816 27652 22880
rect 27716 22816 27732 22880
rect 27796 22816 27812 22880
rect 27876 22816 27892 22880
rect 27956 22816 27972 22880
rect 28036 22816 28044 22880
rect 27644 21792 28044 22816
rect 27644 21728 27652 21792
rect 27716 21728 27732 21792
rect 27796 21728 27812 21792
rect 27876 21728 27892 21792
rect 27956 21728 27972 21792
rect 28036 21728 28044 21792
rect 27644 20704 28044 21728
rect 27644 20640 27652 20704
rect 27716 20640 27732 20704
rect 27796 20640 27812 20704
rect 27876 20640 27892 20704
rect 27956 20640 27972 20704
rect 28036 20640 28044 20704
rect 27644 19616 28044 20640
rect 27644 19552 27652 19616
rect 27716 19552 27732 19616
rect 27796 19552 27812 19616
rect 27876 19552 27892 19616
rect 27956 19552 27972 19616
rect 28036 19552 28044 19616
rect 27644 18528 28044 19552
rect 27644 18464 27652 18528
rect 27716 18464 27732 18528
rect 27796 18464 27812 18528
rect 27876 18464 27892 18528
rect 27956 18464 27972 18528
rect 28036 18464 28044 18528
rect 27644 17440 28044 18464
rect 27644 17376 27652 17440
rect 27716 17376 27732 17440
rect 27796 17376 27812 17440
rect 27876 17376 27892 17440
rect 27956 17376 27972 17440
rect 28036 17376 28044 17440
rect 27644 16352 28044 17376
rect 27644 16288 27652 16352
rect 27716 16288 27732 16352
rect 27796 16288 27812 16352
rect 27876 16288 27892 16352
rect 27956 16288 27972 16352
rect 28036 16288 28044 16352
rect 27644 15264 28044 16288
rect 27644 15200 27652 15264
rect 27716 15200 27732 15264
rect 27796 15200 27812 15264
rect 27876 15200 27892 15264
rect 27956 15200 27972 15264
rect 28036 15200 28044 15264
rect 27644 14176 28044 15200
rect 27644 14112 27652 14176
rect 27716 14112 27732 14176
rect 27796 14112 27812 14176
rect 27876 14112 27892 14176
rect 27956 14112 27972 14176
rect 28036 14112 28044 14176
rect 27644 13088 28044 14112
rect 27644 13024 27652 13088
rect 27716 13024 27732 13088
rect 27796 13024 27812 13088
rect 27876 13024 27892 13088
rect 27956 13024 27972 13088
rect 28036 13024 28044 13088
rect 27644 12000 28044 13024
rect 27644 11936 27652 12000
rect 27716 11936 27732 12000
rect 27796 11936 27812 12000
rect 27876 11936 27892 12000
rect 27956 11936 27972 12000
rect 28036 11936 28044 12000
rect 27644 10912 28044 11936
rect 27644 10848 27652 10912
rect 27716 10848 27732 10912
rect 27796 10848 27812 10912
rect 27876 10848 27892 10912
rect 27956 10848 27972 10912
rect 28036 10848 28044 10912
rect 27644 9824 28044 10848
rect 27644 9760 27652 9824
rect 27716 9760 27732 9824
rect 27796 9760 27812 9824
rect 27876 9760 27892 9824
rect 27956 9760 27972 9824
rect 28036 9760 28044 9824
rect 27644 8736 28044 9760
rect 27644 8672 27652 8736
rect 27716 8672 27732 8736
rect 27796 8672 27812 8736
rect 27876 8672 27892 8736
rect 27956 8672 27972 8736
rect 28036 8672 28044 8736
rect 27644 7648 28044 8672
rect 27644 7584 27652 7648
rect 27716 7584 27732 7648
rect 27796 7584 27812 7648
rect 27876 7584 27892 7648
rect 27956 7584 27972 7648
rect 28036 7584 28044 7648
rect 27644 6560 28044 7584
rect 27644 6496 27652 6560
rect 27716 6496 27732 6560
rect 27796 6496 27812 6560
rect 27876 6496 27892 6560
rect 27956 6496 27972 6560
rect 28036 6496 28044 6560
rect 27644 5472 28044 6496
rect 27644 5408 27652 5472
rect 27716 5408 27732 5472
rect 27796 5408 27812 5472
rect 27876 5408 27892 5472
rect 27956 5408 27972 5472
rect 28036 5408 28044 5472
rect 27644 4384 28044 5408
rect 27644 4320 27652 4384
rect 27716 4320 27732 4384
rect 27796 4320 27812 4384
rect 27876 4320 27892 4384
rect 27956 4320 27972 4384
rect 28036 4320 28044 4384
rect 27644 3296 28044 4320
rect 27644 3232 27652 3296
rect 27716 3232 27732 3296
rect 27796 3232 27812 3296
rect 27876 3232 27892 3296
rect 27956 3232 27972 3296
rect 28036 3232 28044 3296
rect 27644 2208 28044 3232
rect 27644 2144 27652 2208
rect 27716 2144 27732 2208
rect 27796 2144 27812 2208
rect 27876 2144 27892 2208
rect 27956 2144 27972 2208
rect 28036 2144 28044 2208
rect 27644 2128 28044 2144
use sky130_fd_sc_hd__inv_2  _247_
timestamp -25199
transform -1 0 20056 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp -25199
transform 1 0 4416 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp -25199
transform -1 0 4324 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp -25199
transform -1 0 3680 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp -25199
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp -25199
transform 1 0 7544 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp -25199
transform 1 0 2300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp -25199
transform -1 0 3588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp -25199
transform -1 0 5060 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp -25199
transform -1 0 3772 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp -25199
transform -1 0 5520 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp -25199
transform 1 0 2208 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp -25199
transform 1 0 5336 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp -25199
transform 1 0 2208 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp -25199
transform -1 0 6716 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp -25199
transform 1 0 9844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp -25199
transform -1 0 4784 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp -25199
transform 1 0 6532 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp -25199
transform 1 0 6348 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp -25199
transform 1 0 7360 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp -25199
transform -1 0 4508 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp -25199
transform 1 0 5428 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp -25199
transform 1 0 6440 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _270_
timestamp -25199
transform -1 0 24840 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _271_
timestamp -25199
transform 1 0 21804 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _272_
timestamp -25199
transform 1 0 23000 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _273_
timestamp -25199
transform 1 0 9384 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _274_
timestamp -25199
transform 1 0 9936 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _275_
timestamp -25199
transform -1 0 9844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _276_
timestamp -25199
transform 1 0 9016 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _277_
timestamp -25199
transform 1 0 7360 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _278_
timestamp -25199
transform 1 0 9476 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _279_
timestamp -25199
transform -1 0 10488 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _280_
timestamp -25199
transform -1 0 7360 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _281_
timestamp -25199
transform 1 0 5612 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _282_
timestamp -25199
transform -1 0 8740 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _283_
timestamp -25199
transform 1 0 6440 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _284_
timestamp -25199
transform 1 0 5980 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _285_
timestamp -25199
transform 1 0 6348 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _286_
timestamp -25199
transform 1 0 7084 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _287_
timestamp -25199
transform 1 0 8832 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _288_
timestamp -25199
transform 1 0 8372 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _289_
timestamp -25199
transform -1 0 10120 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _290_
timestamp -25199
transform 1 0 9200 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _291_
timestamp -25199
transform -1 0 9660 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _292_
timestamp -25199
transform 1 0 6440 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _293_
timestamp -25199
transform 1 0 7728 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _294_
timestamp -25199
transform 1 0 9108 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _295_
timestamp -25199
transform 1 0 9752 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _296_
timestamp -25199
transform -1 0 9844 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _297_
timestamp -25199
transform 1 0 8832 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _298_
timestamp -25199
transform 1 0 10396 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _299_
timestamp -25199
transform 1 0 9108 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _300_
timestamp -25199
transform 1 0 9292 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _301_
timestamp -25199
transform -1 0 7452 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _302_
timestamp -25199
transform -1 0 8648 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _303_
timestamp -25199
transform -1 0 8004 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _304_
timestamp -25199
transform -1 0 8096 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _305_
timestamp -25199
transform -1 0 7544 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _306_
timestamp -25199
transform 1 0 6808 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _307_
timestamp -25199
transform 1 0 7636 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _308_
timestamp -25199
transform 1 0 5612 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _309_
timestamp -25199
transform 1 0 5796 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _310_
timestamp -25199
transform 1 0 6532 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _311_
timestamp -25199
transform 1 0 7176 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _312_
timestamp -25199
transform -1 0 8832 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _313_
timestamp -25199
transform 1 0 6716 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _314_
timestamp -25199
transform 1 0 7912 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _315_
timestamp -25199
transform -1 0 9660 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _316_
timestamp -25199
transform -1 0 10396 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _317_
timestamp -25199
transform -1 0 10304 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _318_
timestamp -25199
transform 1 0 8924 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _319_
timestamp -25199
transform 1 0 9108 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _320_
timestamp -25199
transform -1 0 8556 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _321_
timestamp -25199
transform 1 0 5244 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _322_
timestamp -25199
transform 1 0 5980 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _323_
timestamp -25199
transform 1 0 6624 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _324_
timestamp -25199
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _325_
timestamp -25199
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _326_
timestamp -25199
transform 1 0 5888 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _327_
timestamp -25199
transform 1 0 5796 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _328_
timestamp -25199
transform 1 0 6348 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _329_
timestamp -25199
transform 1 0 7176 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _330_
timestamp -25199
transform -1 0 7360 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _331_
timestamp -25199
transform 1 0 7268 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _332_
timestamp -25199
transform 1 0 6440 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _333_
timestamp -25199
transform -1 0 7636 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _334_
timestamp -25199
transform 1 0 12328 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _335_
timestamp -25199
transform 1 0 2668 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _336_
timestamp -25199
transform 1 0 1932 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _337_
timestamp -25199
transform -1 0 2852 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _338_
timestamp -25199
transform -1 0 3496 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _339_
timestamp -25199
transform -1 0 3036 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _340_
timestamp -25199
transform 1 0 2024 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _341_
timestamp -25199
transform 1 0 2300 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _342_
timestamp -25199
transform -1 0 3680 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _343_
timestamp -25199
transform -1 0 3404 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _344_
timestamp -25199
transform -1 0 4324 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _345_
timestamp -25199
transform -1 0 3220 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _346_
timestamp -25199
transform 1 0 2392 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _347_
timestamp -25199
transform 1 0 2668 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _348_
timestamp -25199
transform 1 0 2944 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _349_
timestamp -25199
transform 1 0 2760 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _350_
timestamp -25199
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _351_
timestamp -25199
transform 1 0 2392 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _352_
timestamp -25199
transform -1 0 4416 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _353_
timestamp -25199
transform 1 0 3956 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _354_
timestamp -25199
transform -1 0 3956 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _355_
timestamp -25199
transform -1 0 2852 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _356_
timestamp -25199
transform 1 0 2576 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _357_
timestamp -25199
transform 1 0 1748 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _358_
timestamp -25199
transform 1 0 2852 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _359_
timestamp -25199
transform 1 0 3220 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _360_
timestamp -25199
transform 1 0 3680 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _361_
timestamp -25199
transform 1 0 4416 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _362_
timestamp -25199
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _363_
timestamp -25199
transform 1 0 3036 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _364_
timestamp -25199
transform 1 0 3772 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _365_
timestamp -25199
transform 1 0 3036 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _366_
timestamp -25199
transform 1 0 3404 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _367_
timestamp -25199
transform 1 0 3772 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _368_
timestamp -25199
transform -1 0 3404 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _369_
timestamp -25199
transform -1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _370_
timestamp -25199
transform -1 0 3036 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _371_
timestamp -25199
transform 1 0 2576 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _372_
timestamp -25199
transform 1 0 3588 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _373_
timestamp -25199
transform -1 0 3588 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _374_
timestamp -25199
transform 1 0 2944 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _375_
timestamp -25199
transform -1 0 4324 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _376_
timestamp -25199
transform -1 0 3680 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _377_
timestamp -25199
transform -1 0 3404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _378_
timestamp -25199
transform 1 0 3036 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _379_
timestamp -25199
transform -1 0 4600 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp -25199
transform -1 0 12972 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _381_
timestamp -25199
transform -1 0 13800 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _382_
timestamp -25199
transform 1 0 18124 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _383_
timestamp -25199
transform 1 0 18400 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _384_
timestamp -25199
transform -1 0 19228 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _385_
timestamp -25199
transform 1 0 21896 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _386_
timestamp -25199
transform 1 0 21804 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _387_
timestamp -25199
transform 1 0 23368 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _388_
timestamp -25199
transform 1 0 21988 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _389_
timestamp -25199
transform 1 0 23644 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _390_
timestamp -25199
transform 1 0 22172 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _391_
timestamp -25199
transform 1 0 21896 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _392_
timestamp -25199
transform -1 0 21620 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _393_
timestamp -25199
transform 1 0 17848 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _394_
timestamp -25199
transform -1 0 15916 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _395_
timestamp -25199
transform 1 0 12236 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _396_
timestamp -25199
transform 1 0 11500 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _397_
timestamp -25199
transform 1 0 8280 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _398_
timestamp -25199
transform 1 0 7452 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _399_
timestamp -25199
transform 1 0 4140 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _400_
timestamp -25199
transform 1 0 2576 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _401_
timestamp -25199
transform 1 0 7268 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp -25199
transform 1 0 7084 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _403_
timestamp -25199
transform -1 0 12328 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _404_
timestamp -25199
transform 1 0 11592 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _405_
timestamp -25199
transform 1 0 14444 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _406_
timestamp -25199
transform -1 0 14904 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _407_
timestamp -25199
transform 1 0 16192 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _408_
timestamp -25199
transform 1 0 14720 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _409_
timestamp -25199
transform 1 0 20700 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _410_
timestamp -25199
transform -1 0 23920 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _411_
timestamp -25199
transform 1 0 24380 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp -25199
transform 1 0 24380 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _413_
timestamp -25199
transform -1 0 24840 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _414_
timestamp -25199
transform 1 0 24472 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _415_
timestamp -25199
transform -1 0 25208 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _416_
timestamp -25199
transform 1 0 22632 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _417_
timestamp -25199
transform 1 0 20056 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _418_
timestamp -25199
transform 1 0 18676 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _419_
timestamp -25199
transform -1 0 17940 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _420_
timestamp -25199
transform 1 0 12144 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _421_
timestamp -25199
transform -1 0 11316 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _422_
timestamp -25199
transform 1 0 8924 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _423_
timestamp -25199
transform 1 0 4416 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _424_
timestamp -25199
transform -1 0 5612 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _425_
timestamp -25199
transform 1 0 4784 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _426_
timestamp -25199
transform -1 0 8464 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _427_
timestamp -25199
transform 1 0 10212 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _428_
timestamp -25199
transform -1 0 12512 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _429_
timestamp -25199
transform -1 0 14812 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _430_
timestamp -25199
transform -1 0 16100 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _431_
timestamp -25199
transform 1 0 15272 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _432_
timestamp -25199
transform -1 0 16192 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _433_
timestamp -25199
transform -1 0 16376 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _434_
timestamp -25199
transform 1 0 18676 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _435_
timestamp -25199
transform 1 0 17664 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _436_
timestamp -25199
transform -1 0 19872 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _437_
timestamp -25199
transform 1 0 18676 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _438_
timestamp -25199
transform 1 0 18308 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _439_
timestamp -25199
transform 1 0 19504 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _440_
timestamp -25199
transform 1 0 19228 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _441_
timestamp -25199
transform 1 0 20332 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _442_
timestamp -25199
transform 1 0 19504 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _443_
timestamp -25199
transform 1 0 18400 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _444_
timestamp -25199
transform 1 0 16652 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _445_
timestamp -25199
transform 1 0 16652 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _446_
timestamp -25199
transform 1 0 14352 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _447_
timestamp -25199
transform 1 0 13524 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _448_
timestamp -25199
transform 1 0 12236 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _449_
timestamp -25199
transform 1 0 10580 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _450_
timestamp -25199
transform -1 0 10396 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _451_
timestamp -25199
transform 1 0 7544 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _452_
timestamp -25199
transform 1 0 3404 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _453_
timestamp -25199
transform -1 0 4324 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _454_
timestamp -25199
transform -1 0 7176 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _455_
timestamp -25199
transform -1 0 9476 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _456_
timestamp -25199
transform 1 0 9660 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _457_
timestamp -25199
transform 1 0 12788 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _458_
timestamp -25199
transform 1 0 12052 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _459_
timestamp -25199
transform 1 0 12696 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _460_
timestamp -25199
transform 1 0 12144 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _461_
timestamp -25199
transform 1 0 20976 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _462_
timestamp -25199
transform -1 0 20332 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _463_
timestamp -25199
transform 1 0 23184 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _464_
timestamp -25199
transform -1 0 21344 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _465_
timestamp -25199
transform 1 0 24196 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _466_
timestamp -25199
transform -1 0 21988 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _467_
timestamp -25199
transform 1 0 21804 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _468_
timestamp -25199
transform 1 0 19228 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _469_
timestamp -25199
transform 1 0 18032 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _470_
timestamp -25199
transform 1 0 16008 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _471_
timestamp -25199
transform 1 0 14260 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _472_
timestamp -25199
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _473_
timestamp -25199
transform 1 0 7544 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _474_
timestamp -25199
transform 1 0 10856 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _475_
timestamp -25199
transform 1 0 4692 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _476_
timestamp -25199
transform 1 0 7820 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _477_
timestamp -25199
transform 1 0 7176 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _478_
timestamp -25199
transform 1 0 3772 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _479_
timestamp -25199
transform 1 0 2576 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _480_
timestamp -25199
transform -1 0 9752 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _481_
timestamp -25199
transform 1 0 14076 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _482_
timestamp -25199
transform -1 0 12788 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _483_
timestamp -25199
transform 1 0 14444 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _484_
timestamp -25199
transform 1 0 12696 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _485_
timestamp -25199
transform 1 0 12052 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _486_
timestamp -25199
transform -1 0 22448 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _487_
timestamp -25199
transform 1 0 20976 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _488_
timestamp -25199
transform 1 0 20884 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _489_
timestamp -25199
transform 1 0 23276 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _490_
timestamp -25199
transform -1 0 23644 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _491_
timestamp -25199
transform 1 0 23276 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _492_
timestamp -25199
transform -1 0 23000 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _493_
timestamp -25199
transform -1 0 23000 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _494_
timestamp -25199
transform 1 0 22816 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _495_
timestamp -25199
transform 1 0 24380 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _496_
timestamp -25199
transform 1 0 17848 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _497_
timestamp -25199
transform 1 0 17664 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _498_
timestamp -25199
transform -1 0 22448 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _499_
timestamp -25199
transform 1 0 21804 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _500_
timestamp -25199
transform 1 0 21804 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _501_
timestamp -25199
transform -1 0 21712 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _502_
timestamp -25199
transform -1 0 16008 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _503_
timestamp -25199
transform -1 0 12236 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _504_
timestamp -25199
transform 1 0 6900 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _505_
timestamp -25199
transform 1 0 1380 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _506_
timestamp -25199
transform 1 0 6348 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _507_
timestamp -25199
transform 1 0 11500 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _508_
timestamp -25199
transform -1 0 15364 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _509_
timestamp -25199
transform 1 0 14168 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _510_
timestamp -25199
transform 1 0 21344 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _511_
timestamp -25199
transform 1 0 23920 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _512_
timestamp -25199
transform 1 0 24380 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _513_
timestamp -25199
transform -1 0 25116 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _514_
timestamp -25199
transform 1 0 19228 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _515_
timestamp -25199
transform -1 0 18124 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _516_
timestamp -25199
transform -1 0 11316 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _517_
timestamp -25199
transform 1 0 3772 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _518_
timestamp -25199
transform 1 0 4324 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _519_
timestamp -25199
transform 1 0 9844 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _520_
timestamp -25199
transform 1 0 14076 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _521_
timestamp -25199
transform 1 0 14904 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _522_
timestamp -25199
transform -1 0 16284 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _523_
timestamp -25199
transform 1 0 16836 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _524_
timestamp -25199
transform 1 0 16928 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _525_
timestamp -25199
transform 1 0 17296 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _526_
timestamp -25199
transform 1 0 17296 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _527_
timestamp -25199
transform 1 0 17848 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _528_
timestamp -25199
transform -1 0 19504 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _529_
timestamp -25199
transform -1 0 17388 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _530_
timestamp -25199
transform 1 0 14076 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _531_
timestamp -25199
transform -1 0 13156 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _532_
timestamp -25199
transform -1 0 10764 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _533_
timestamp -25199
transform 1 0 1564 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _534_
timestamp -25199
transform -1 0 7084 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _535_
timestamp -25199
transform 1 0 9384 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _536_
timestamp -25199
transform 1 0 11500 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _537_
timestamp -25199
transform 1 0 11408 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _538_
timestamp -25199
transform 1 0 21804 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _539_
timestamp -25199
transform 1 0 23000 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _540_
timestamp -25199
transform 1 0 23368 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _541_
timestamp -25199
transform 1 0 21068 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _542_
timestamp -25199
transform 1 0 17388 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _543_
timestamp -25199
transform 1 0 14076 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _544_
timestamp -25199
transform 1 0 6532 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _545_
timestamp -25199
transform 1 0 3772 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _546_
timestamp -25199
transform 1 0 6440 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _547_
timestamp -25199
transform 1 0 1748 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _548_
timestamp -25199
transform 1 0 13800 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _549_
timestamp -25199
transform 1 0 14168 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _550_
timestamp -25199
transform 1 0 11316 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _551_
timestamp -25199
transform 1 0 19780 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _552_
timestamp -25199
transform 1 0 24380 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _553_
timestamp -25199
transform 1 0 23000 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _554_
timestamp -25199
transform 1 0 20516 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A0
timestamp -25199
transform -1 0 19136 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__S
timestamp -25199
transform 1 0 12328 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__S
timestamp -25199
transform -1 0 8556 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__S
timestamp -25199
transform 1 0 4968 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__S
timestamp -25199
transform 1 0 7084 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__403__S
timestamp -25199
transform -1 0 11408 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__S
timestamp -25199
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__S
timestamp -25199
transform 1 0 16008 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__S
timestamp -25199
transform 1 0 11960 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__S
timestamp -25199
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__S
timestamp -25199
transform 1 0 5612 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__S
timestamp -25199
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__S
timestamp -25199
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__S
timestamp -25199
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__S
timestamp -25199
transform 1 0 15180 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__S
timestamp -25199
transform 1 0 12052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__S
timestamp -25199
transform 1 0 9384 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__456__S
timestamp -25199
transform 1 0 9476 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__458__S
timestamp -25199
transform 1 0 11868 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__S
timestamp -25199
transform -1 0 12144 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__S
timestamp -25199
transform -1 0 10856 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__S
timestamp -25199
transform 1 0 7636 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__S
timestamp -25199
transform 1 0 4600 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__S
timestamp -25199
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__485__S
timestamp -25199
transform -1 0 12052 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__Q
timestamp -25199
transform 1 0 19688 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__532__RESET_B
timestamp -25199
transform 1 0 8740 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__535__RESET_B
timestamp -25199
transform 1 0 9200 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__536__RESET_B
timestamp -25199
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__537__RESET_B
timestamp -25199
transform -1 0 11408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__550__RESET_B
timestamp -25199
transform 1 0 11132 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp -25199
transform 1 0 13064 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp -25199
transform 1 0 15088 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_clk_A
timestamp -25199
transform -1 0 9016 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_clk_A
timestamp -25199
transform -1 0 13524 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_clk_A
timestamp -25199
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_clk_A
timestamp -25199
transform 1 0 13248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_clk_A
timestamp -25199
transform 1 0 19320 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_clk_A
timestamp -25199
transform 1 0 20424 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_clk_A
timestamp -25199
transform -1 0 17020 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_clk_A
timestamp -25199
transform -1 0 20148 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout46_A
timestamp -25199
transform -1 0 3680 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout47_A
timestamp -25199
transform 1 0 4324 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout47_X
timestamp -25199
transform 1 0 4140 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout52_A
timestamp -25199
transform 1 0 15824 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout56_A
timestamp -25199
transform 1 0 16468 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout57_X
timestamp -25199
transform 1 0 3588 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout60_A
timestamp -25199
transform -1 0 3404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout61_A
timestamp -25199
transform -1 0 2300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout61_X
timestamp -25199
transform 1 0 3128 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout66_A
timestamp -25199
transform 1 0 14352 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout71_A
timestamp -25199
transform -1 0 16836 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout72_X
timestamp -25199
transform 1 0 2300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout74_A
timestamp -25199
transform 1 0 18124 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout75_A
timestamp -25199
transform -1 0 4140 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout75_X
timestamp -25199
transform -1 0 4324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout77_A
timestamp -25199
transform -1 0 15732 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout78_A
timestamp -25199
transform -1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout79_X
timestamp -25199
transform 1 0 4508 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout81_A
timestamp -25199
transform 1 0 18216 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout82_A
timestamp -25199
transform -1 0 6256 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout82_X
timestamp -25199
transform 1 0 5888 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp -25199
transform -1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_X
timestamp -25199
transform 1 0 1748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp -25199
transform -1 0 2392 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp -25199
transform -1 0 2576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_X
timestamp -25199
transform 1 0 2024 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp -25199
transform -1 0 2760 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp -25199
transform -1 0 1564 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp -25199
transform -1 0 1564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp -25199
transform -1 0 1840 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp -25199
transform -1 0 1840 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp -25199
transform -1 0 2024 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp -25199
transform -1 0 1840 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp -25199
transform -1 0 2760 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp -25199
transform -1 0 2484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp -25199
transform -1 0 2024 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp -25199
transform -1 0 1840 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp -25199
transform -1 0 1932 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp -25199
transform -1 0 2024 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp -25199
transform -1 0 1840 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp -25199
transform -1 0 1932 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp -25199
transform -1 0 1932 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp -25199
transform -1 0 1932 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp -25199
transform -1 0 1932 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp -25199
transform -1 0 1932 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp -25199
transform -1 0 1932 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp -25199
transform -1 0 1840 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp -25199
transform -1 0 1840 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp -25199
transform -1 0 1840 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp -25199
transform -1 0 1840 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp -25199
transform -1 0 1840 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp -25199
transform -1 0 2024 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp -25199
transform -1 0 1932 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp -25199
transform -1 0 1932 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp -25199
transform -1 0 1932 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp -25199
transform -1 0 2116 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp -25199
transform -1 0 1840 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp -25199
transform -1 0 1932 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp -25199
transform -1 0 1932 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp -25199
transform -1 0 1840 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp -25199
transform -1 0 1840 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output39_A
timestamp -25199
transform 1 0 27876 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -25199
transform 1 0 13248 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp -25199
transform -1 0 8832 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp -25199
transform 1 0 11500 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp -25199
transform -1 0 10764 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp -25199
transform 1 0 11408 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp -25199
transform 1 0 19504 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp -25199
transform 1 0 20608 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp -25199
transform -1 0 18860 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp -25199
transform 1 0 20148 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp -25199
transform 1 0 6992 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload1
timestamp -25199
transform 1 0 10856 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  clkload2
timestamp -25199
transform 1 0 8188 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload3
timestamp -25199
transform -1 0 11408 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload4
timestamp -25199
transform 1 0 18124 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  clkload5
timestamp -25199
transform 1 0 20148 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout41
timestamp -25199
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout42
timestamp -25199
transform 1 0 11684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout43
timestamp -25199
transform 1 0 4324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout44
timestamp -25199
transform 1 0 3496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout45
timestamp -25199
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout46
timestamp -25199
transform -1 0 3496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp -25199
transform -1 0 4140 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout48
timestamp -25199
transform -1 0 15180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout49
timestamp -25199
transform 1 0 17756 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout50
timestamp -25199
transform 1 0 21712 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout51
timestamp -25199
transform 1 0 19228 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout52
timestamp -25199
transform 1 0 15548 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout53
timestamp -25199
transform 1 0 15640 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout54
timestamp -25199
transform 1 0 15272 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout55
timestamp -25199
transform 1 0 21620 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout56
timestamp -25199
transform 1 0 16652 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout57
timestamp -25199
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout58
timestamp -25199
transform 1 0 2024 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout59
timestamp -25199
transform -1 0 2760 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp -25199
transform -1 0 3128 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout61
timestamp -25199
transform 1 0 2760 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout62
timestamp -25199
transform 1 0 15180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout63
timestamp -25199
transform 1 0 17388 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout64
timestamp -25199
transform -1 0 21436 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout65
timestamp -25199
transform -1 0 23184 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout66
timestamp -25199
transform 1 0 14536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout67
timestamp -25199
transform -1 0 16468 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout68
timestamp -25199
transform -1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout69
timestamp -25199
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout70
timestamp -25199
transform 1 0 21620 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout71
timestamp -25199
transform 1 0 16744 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout72
timestamp -25199
transform 1 0 2484 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout73
timestamp -25199
transform 1 0 2576 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout74
timestamp -25199
transform 1 0 18308 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout75
timestamp -25199
transform 1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout76
timestamp -25199
transform -1 0 7084 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout77
timestamp -25199
transform 1 0 15180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout78
timestamp -25199
transform 1 0 13340 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout79
timestamp -25199
transform 1 0 4140 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout80
timestamp -25199
transform 1 0 3404 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout81
timestamp -25199
transform 1 0 18400 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout82
timestamp -25199
transform 1 0 5520 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636943256
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636943256
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -25199
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636943256
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636943256
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -25199
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636943256
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636943256
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -25199
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636943256
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636943256
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -25199
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636943256
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636943256
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -25199
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636943256
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636943256
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -25199
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636943256
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636943256
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -25199
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636943256
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636943256
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -25199
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636943256
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636943256
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -25199
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636943256
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636943256
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -25199
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636943256
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_293
timestamp -25199
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636943256
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636943256
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_27
timestamp -25199
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_35
timestamp -25199
transform 1 0 4324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_45
timestamp -25199
transform 1 0 5244 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp -25199
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636943256
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_69
timestamp -25199
transform 1 0 7452 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_79
timestamp 1636943256
transform 1 0 8372 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -25199
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp -25199
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp -25199
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_129
timestamp 1636943256
transform 1 0 12972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_141
timestamp 1636943256
transform 1 0 14076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_153
timestamp 1636943256
transform 1 0 15180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp -25199
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp -25199
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_173
timestamp -25199
transform 1 0 17020 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_183
timestamp 1636943256
transform 1 0 17940 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_195
timestamp -25199
transform 1 0 19044 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_203
timestamp -25199
transform 1 0 19780 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_215
timestamp -25199
transform 1 0 20884 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp -25199
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636943256
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636943256
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636943256
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636943256
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp -25199
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp -25199
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636943256
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_293
timestamp -25199
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636943256
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636943256
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -25199
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_49
timestamp -25199
transform 1 0 5612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_57
timestamp -25199
transform 1 0 6348 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_81
timestamp -25199
transform 1 0 8556 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_94
timestamp -25199
transform 1 0 9752 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_100
timestamp -25199
transform 1 0 10304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_130
timestamp -25199
transform 1 0 13064 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp -25199
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_161
timestamp -25199
transform 1 0 15916 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_185
timestamp -25199
transform 1 0 18124 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp -25199
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_237
timestamp 1636943256
transform 1 0 22908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp -25199
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636943256
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636943256
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636943256
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_289
timestamp -25199
transform 1 0 27692 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_297
timestamp -25199
transform 1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636943256
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_15
timestamp -25199
transform 1 0 2484 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_25
timestamp -25199
transform 1 0 3404 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_44
timestamp 1636943256
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636943256
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_87
timestamp 1636943256
transform 1 0 9108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_99
timestamp -25199
transform 1 0 10212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -25199
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_124
timestamp 1636943256
transform 1 0 12512 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_136
timestamp -25199
transform 1 0 13616 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp -25199
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636943256
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_181
timestamp -25199
transform 1 0 17756 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_200
timestamp 1636943256
transform 1 0 19504 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_212
timestamp 1636943256
transform 1 0 20608 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_243
timestamp 1636943256
transform 1 0 23460 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_255
timestamp 1636943256
transform 1 0 24564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_267
timestamp 1636943256
transform 1 0 25668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp -25199
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636943256
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp -25199
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_25
timestamp -25199
transform 1 0 3404 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_49
timestamp 1636943256
transform 1 0 5612 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_61
timestamp -25199
transform 1 0 6716 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -25199
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636943256
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636943256
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636943256
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636943256
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp -25199
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp -25199
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp -25199
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_161
timestamp 1636943256
transform 1 0 15916 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_173
timestamp 1636943256
transform 1 0 17020 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_191
timestamp -25199
transform 1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp -25199
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636943256
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636943256
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_221
timestamp -25199
transform 1 0 21436 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_225
timestamp -25199
transform 1 0 21804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_235
timestamp 1636943256
transform 1 0 22724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_247
timestamp -25199
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp -25199
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_262
timestamp 1636943256
transform 1 0 25208 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_274
timestamp 1636943256
transform 1 0 26312 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_286
timestamp 1636943256
transform 1 0 27416 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_298
timestamp -25199
transform 1 0 28520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_8
timestamp -25199
transform 1 0 1840 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_30
timestamp -25199
transform 1 0 3864 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636943256
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636943256
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636943256
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636943256
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp -25199
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -25199
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636943256
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636943256
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636943256
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636943256
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp -25199
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -25199
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp -25199
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_197
timestamp 1636943256
transform 1 0 19228 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_209
timestamp -25199
transform 1 0 20332 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_213
timestamp -25199
transform 1 0 20700 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp -25199
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636943256
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp -25199
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636943256
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp -25199
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp -25199
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636943256
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp -25199
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_6_8
timestamp -25199
transform 1 0 1840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_22
timestamp -25199
transform 1 0 3128 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -25199
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_37
timestamp -25199
transform 1 0 4508 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_51
timestamp 1636943256
transform 1 0 5796 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_63
timestamp -25199
transform 1 0 6900 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_69
timestamp -25199
transform 1 0 7452 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp -25199
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp -25199
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636943256
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_97
timestamp -25199
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_103
timestamp -25199
transform 1 0 10580 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_115
timestamp -25199
transform 1 0 11684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_130
timestamp -25199
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp -25199
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_150
timestamp 1636943256
transform 1 0 14904 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_171
timestamp 1636943256
transform 1 0 16836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_183
timestamp -25199
transform 1 0 17940 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp -25199
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_197
timestamp -25199
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_203
timestamp -25199
transform 1 0 19780 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_228
timestamp 1636943256
transform 1 0 22080 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_240
timestamp 1636943256
transform 1 0 23184 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636943256
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636943256
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1636943256
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_289
timestamp -25199
transform 1 0 27692 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_297
timestamp -25199
transform 1 0 28428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_11
timestamp -25199
transform 1 0 2116 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_19
timestamp -25199
transform 1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_24
timestamp -25199
transform 1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_29
timestamp 1636943256
transform 1 0 3772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_41
timestamp 1636943256
transform 1 0 4876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp -25199
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_57
timestamp -25199
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_63
timestamp -25199
transform 1 0 6900 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_70
timestamp -25199
transform 1 0 7544 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_82
timestamp -25199
transform 1 0 8648 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_86
timestamp -25199
transform 1 0 9016 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp -25199
transform 1 0 10396 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_159
timestamp -25199
transform 1 0 15732 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -25199
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_178
timestamp 1636943256
transform 1 0 17480 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_190
timestamp 1636943256
transform 1 0 18584 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_202
timestamp 1636943256
transform 1 0 19688 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_214
timestamp -25199
transform 1 0 20792 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_221
timestamp -25199
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636943256
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636943256
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636943256
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1636943256
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp -25199
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp -25199
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636943256
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp -25199
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_16
timestamp 1636943256
transform 1 0 2576 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp -25199
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_37
timestamp -25199
transform 1 0 4508 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_49
timestamp 1636943256
transform 1 0 5612 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_61
timestamp -25199
transform 1 0 6716 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_105
timestamp -25199
transform 1 0 10764 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_110
timestamp -25199
transform 1 0 11224 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_131
timestamp -25199
transform 1 0 13156 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_135
timestamp -25199
transform 1 0 13524 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_161
timestamp 1636943256
transform 1 0 15916 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_173
timestamp 1636943256
transform 1 0 17020 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_185
timestamp -25199
transform 1 0 18124 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp -25199
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_206
timestamp 1636943256
transform 1 0 20056 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_218
timestamp -25199
transform 1 0 21160 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_226
timestamp -25199
transform 1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_238
timestamp 1636943256
transform 1 0 23000 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp -25199
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636943256
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1636943256
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1636943256
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_289
timestamp -25199
transform 1 0 27692 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_297
timestamp -25199
transform 1 0 28428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_34
timestamp -25199
transform 1 0 4232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -25199
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp -25199
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_65
timestamp -25199
transform 1 0 7084 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_75
timestamp -25199
transform 1 0 8004 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_85
timestamp 1636943256
transform 1 0 8924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_97
timestamp 1636943256
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp -25199
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636943256
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636943256
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_137
timestamp -25199
transform 1 0 13708 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_143
timestamp -25199
transform 1 0 14260 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_162
timestamp -25199
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_178
timestamp -25199
transform 1 0 17480 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_186
timestamp -25199
transform 1 0 18216 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_197
timestamp 1636943256
transform 1 0 19228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_209
timestamp 1636943256
transform 1 0 20332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp -25199
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_263
timestamp 1636943256
transform 1 0 25300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp -25199
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp -25199
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636943256
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp -25199
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_18
timestamp -25199
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp -25199
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_40
timestamp 1636943256
transform 1 0 4784 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_52
timestamp -25199
transform 1 0 5888 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_78
timestamp -25199
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636943256
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1636943256
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1636943256
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1636943256
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp -25199
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp -25199
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636943256
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp -25199
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_184
timestamp -25199
transform 1 0 18032 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp -25199
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp -25199
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_197
timestamp -25199
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_227
timestamp 1636943256
transform 1 0 21988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_239
timestamp 1636943256
transform 1 0 23092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp -25199
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_273
timestamp 1636943256
transform 1 0 26220 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_285
timestamp -25199
transform 1 0 27324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_13
timestamp -25199
transform 1 0 2300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_25
timestamp -25199
transform 1 0 3404 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1636943256
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp -25199
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp -25199
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636943256
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_80
timestamp 1636943256
transform 1 0 8464 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_92
timestamp -25199
transform 1 0 9568 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_98
timestamp -25199
transform 1 0 10120 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp -25199
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_115
timestamp 1636943256
transform 1 0 11684 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_127
timestamp 1636943256
transform 1 0 12788 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_139
timestamp 1636943256
transform 1 0 13892 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_151
timestamp 1636943256
transform 1 0 14996 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_163
timestamp -25199
transform 1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp -25199
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_169
timestamp -25199
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_177
timestamp -25199
transform 1 0 17388 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp -25199
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_245
timestamp -25199
transform 1 0 23644 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_258
timestamp 1636943256
transform 1 0 24840 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_270
timestamp -25199
transform 1 0 25944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp -25199
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1636943256
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp -25199
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_5
timestamp -25199
transform 1 0 1564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp -25199
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_39
timestamp 1636943256
transform 1 0 4692 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_51
timestamp 1636943256
transform 1 0 5796 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_63
timestamp -25199
transform 1 0 6900 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_76
timestamp -25199
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp -25199
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp -25199
transform 1 0 9660 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_124
timestamp 1636943256
transform 1 0 12512 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp -25199
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_161
timestamp 1636943256
transform 1 0 15916 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_173
timestamp 1636943256
transform 1 0 17020 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_185
timestamp -25199
transform 1 0 18124 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp -25199
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1636943256
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_209
timestamp -25199
transform 1 0 20332 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_232
timestamp -25199
transform 1 0 22448 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_236
timestamp -25199
transform 1 0 22816 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_240
timestamp 1636943256
transform 1 0 23184 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1636943256
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1636943256
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1636943256
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_289
timestamp -25199
transform 1 0 27692 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_297
timestamp -25199
transform 1 0 28428 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_8
timestamp 1636943256
transform 1 0 1840 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_20
timestamp 1636943256
transform 1 0 2944 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_32
timestamp 1636943256
transform 1 0 4048 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_44
timestamp 1636943256
transform 1 0 5152 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_66
timestamp 1636943256
transform 1 0 7176 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_78
timestamp 1636943256
transform 1 0 8280 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_90
timestamp 1636943256
transform 1 0 9384 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_102
timestamp -25199
transform 1 0 10488 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_122
timestamp 1636943256
transform 1 0 12328 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_134
timestamp -25199
transform 1 0 13432 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1636943256
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp -25199
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp -25199
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1636943256
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_181
timestamp -25199
transform 1 0 17756 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_202
timestamp 1636943256
transform 1 0 19688 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_214
timestamp -25199
transform 1 0 20792 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp -25199
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp -25199
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_236
timestamp -25199
transform 1 0 22816 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_262
timestamp 1636943256
transform 1 0 25208 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_274
timestamp -25199
transform 1 0 26312 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1636943256
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_293
timestamp -25199
transform 1 0 28060 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_8
timestamp 1636943256
transform 1 0 1840 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp -25199
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636943256
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp -25199
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_74
timestamp -25199
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_94
timestamp 1636943256
transform 1 0 9752 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_106
timestamp -25199
transform 1 0 10856 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_123
timestamp 1636943256
transform 1 0 12420 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp -25199
transform 1 0 13524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp -25199
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_150
timestamp 1636943256
transform 1 0 14904 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_162
timestamp 1636943256
transform 1 0 16008 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_174
timestamp 1636943256
transform 1 0 17112 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_186
timestamp -25199
transform 1 0 18216 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp -25199
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_206
timestamp 1636943256
transform 1 0 20056 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_218
timestamp 1636943256
transform 1 0 21160 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_230
timestamp 1636943256
transform 1 0 22264 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_242
timestamp -25199
transform 1 0 23368 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp -25199
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1636943256
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1636943256
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1636943256
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_289
timestamp -25199
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp -25199
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_10
timestamp 1636943256
transform 1 0 2024 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_22
timestamp -25199
transform 1 0 3128 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_33
timestamp 1636943256
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp -25199
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp -25199
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_77
timestamp -25199
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_81
timestamp -25199
transform 1 0 8556 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_102
timestamp -25199
transform 1 0 10488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp -25199
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_133
timestamp -25199
transform 1 0 13340 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_137
timestamp -25199
transform 1 0 13708 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_158
timestamp -25199
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp -25199
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1636943256
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1636943256
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_193
timestamp -25199
transform 1 0 18860 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_200
timestamp -25199
transform 1 0 19504 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_208
timestamp -25199
transform 1 0 20240 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp -25199
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1636943256
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp -25199
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_241
timestamp -25199
transform 1 0 23276 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_260
timestamp 1636943256
transform 1 0 25024 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_272
timestamp -25199
transform 1 0 26128 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1636943256
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp -25199
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_6
timestamp -25199
transform 1 0 1656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_14
timestamp -25199
transform 1 0 2392 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_42
timestamp 1636943256
transform 1 0 4968 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_54
timestamp 1636943256
transform 1 0 6072 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_66
timestamp -25199
transform 1 0 7176 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_74
timestamp -25199
transform 1 0 7912 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_107
timestamp 1636943256
transform 1 0 10948 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_119
timestamp 1636943256
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_131
timestamp -25199
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp -25199
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp -25199
transform 1 0 16100 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_169
timestamp -25199
transform 1 0 16652 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_175
timestamp -25199
transform 1 0 17204 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp -25199
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_209
timestamp -25199
transform 1 0 20332 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_232
timestamp 1636943256
transform 1 0 22448 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp -25199
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_262
timestamp 1636943256
transform 1 0 25208 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_274
timestamp 1636943256
transform 1 0 26312 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_286
timestamp 1636943256
transform 1 0 27416 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_298
timestamp -25199
transform 1 0 28520 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_18
timestamp -25199
transform 1 0 2760 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_26
timestamp 1636943256
transform 1 0 3496 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_38
timestamp 1636943256
transform 1 0 4600 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_50
timestamp -25199
transform 1 0 5704 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636943256
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1636943256
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_81
timestamp -25199
transform 1 0 8556 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_87
timestamp -25199
transform 1 0 9108 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp -25199
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1636943256
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_125
timestamp -25199
transform 1 0 12604 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_129
timestamp -25199
transform 1 0 12972 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp -25199
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_179
timestamp -25199
transform 1 0 17572 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_196
timestamp 1636943256
transform 1 0 19136 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_208
timestamp 1636943256
transform 1 0 20240 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp -25199
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_234
timestamp -25199
transform 1 0 22632 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_258
timestamp 1636943256
transform 1 0 24840 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_270
timestamp -25199
transform 1 0 25944 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp -25199
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1636943256
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_293
timestamp -25199
transform 1 0 28060 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_15
timestamp -25199
transform 1 0 2484 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_22
timestamp -25199
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_29
timestamp -25199
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_35
timestamp 1636943256
transform 1 0 4324 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_47
timestamp 1636943256
transform 1 0 5428 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_59
timestamp 1636943256
transform 1 0 6532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_71
timestamp 1636943256
transform 1 0 7636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp -25199
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1636943256
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1636943256
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_109
timestamp -25199
transform 1 0 11132 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp -25199
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_141
timestamp -25199
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_149
timestamp -25199
transform 1 0 14812 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_180
timestamp 1636943256
transform 1 0 17664 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp -25199
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1636943256
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1636943256
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp -25199
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_227
timestamp 1636943256
transform 1 0 21988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_239
timestamp -25199
transform 1 0 23092 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_249
timestamp -25199
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_257
timestamp 1636943256
transform 1 0 24748 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_269
timestamp 1636943256
transform 1 0 25852 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_281
timestamp 1636943256
transform 1 0 26956 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_293
timestamp -25199
transform 1 0 28060 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_10
timestamp -25199
transform 1 0 2024 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_19
timestamp -25199
transform 1 0 2852 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_26
timestamp 1636943256
transform 1 0 3496 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_38
timestamp 1636943256
transform 1 0 4600 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp -25199
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_64
timestamp 1636943256
transform 1 0 6992 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_76
timestamp -25199
transform 1 0 8096 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_89
timestamp 1636943256
transform 1 0 9292 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_101
timestamp -25199
transform 1 0 10396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_109
timestamp -25199
transform 1 0 11132 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_143
timestamp 1636943256
transform 1 0 14260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_155
timestamp -25199
transform 1 0 15364 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp -25199
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_171
timestamp 1636943256
transform 1 0 16836 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_183
timestamp -25199
transform 1 0 17940 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_209
timestamp 1636943256
transform 1 0 20332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_221
timestamp -25199
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1636943256
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1636943256
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1636943256
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1636943256
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp -25199
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp -25199
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1636943256
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp -25199
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_13
timestamp 1636943256
transform 1 0 2300 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_39
timestamp 1636943256
transform 1 0 4692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_51
timestamp -25199
transform 1 0 5796 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_73
timestamp -25199
transform 1 0 7820 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_98
timestamp -25199
transform 1 0 10120 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp -25199
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp -25199
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_154
timestamp 1636943256
transform 1 0 15272 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_166
timestamp 1636943256
transform 1 0 16376 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_178
timestamp 1636943256
transform 1 0 17480 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp -25199
transform 1 0 18584 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1636943256
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1636943256
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1636943256
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1636943256
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp -25199
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp -25199
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_262
timestamp 1636943256
transform 1 0 25208 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_274
timestamp 1636943256
transform 1 0 26312 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_286
timestamp 1636943256
transform 1 0 27416 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_298
timestamp -25199
transform 1 0 28520 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_9
timestamp -25199
transform 1 0 1932 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_17
timestamp -25199
transform 1 0 2668 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_34
timestamp 1636943256
transform 1 0 4232 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_46
timestamp -25199
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp -25199
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_57
timestamp -25199
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_63
timestamp -25199
transform 1 0 6900 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_71
timestamp -25199
transform 1 0 7636 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_80
timestamp -25199
transform 1 0 8464 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1636943256
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp -25199
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp -25199
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_113
timestamp -25199
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_128
timestamp 1636943256
transform 1 0 12880 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_140
timestamp -25199
transform 1 0 13984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp -25199
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_169
timestamp -25199
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_177
timestamp -25199
transform 1 0 17388 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_200
timestamp 1636943256
transform 1 0 19504 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_212
timestamp 1636943256
transform 1 0 20608 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_225
timestamp -25199
transform 1 0 21804 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_235
timestamp -25199
transform 1 0 22724 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_268
timestamp 1636943256
transform 1 0 25760 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1636943256
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_293
timestamp -25199
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_10
timestamp -25199
transform 1 0 2024 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_18
timestamp -25199
transform 1 0 2760 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp -25199
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_35
timestamp 1636943256
transform 1 0 4324 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_47
timestamp 1636943256
transform 1 0 5428 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_59
timestamp 1636943256
transform 1 0 6532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_71
timestamp 1636943256
transform 1 0 7636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp -25199
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1636943256
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1636943256
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1636943256
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1636943256
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp -25199
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp -25199
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1636943256
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_173
timestamp -25199
transform 1 0 17020 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_204
timestamp -25199
transform 1 0 19872 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_212
timestamp -25199
transform 1 0 20608 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_240
timestamp 1636943256
transform 1 0 23184 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1636943256
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1636943256
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1636943256
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_289
timestamp -25199
transform 1 0 27692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_297
timestamp -25199
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_9
timestamp -25199
transform 1 0 1932 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_21
timestamp -25199
transform 1 0 3036 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_35
timestamp 1636943256
transform 1 0 4324 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp -25199
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp -25199
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1636943256
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1636943256
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_81
timestamp -25199
transform 1 0 8556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_85
timestamp -25199
transform 1 0 8924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_98
timestamp 1636943256
transform 1 0 10120 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp -25199
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1636943256
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_125
timestamp -25199
transform 1 0 12604 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_135
timestamp 1636943256
transform 1 0 13524 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_147
timestamp 1636943256
transform 1 0 14628 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_159
timestamp -25199
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp -25199
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1636943256
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_181
timestamp -25199
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_189
timestamp -25199
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_197
timestamp -25199
transform 1 0 19228 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_205
timestamp -25199
transform 1 0 19964 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_213
timestamp -25199
transform 1 0 20700 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp -25199
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_245
timestamp 1636943256
transform 1 0 23644 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_257
timestamp 1636943256
transform 1 0 24748 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_269
timestamp -25199
transform 1 0 25852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp -25199
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1636943256
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_293
timestamp -25199
transform 1 0 28060 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp -25199
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_32
timestamp 1636943256
transform 1 0 4048 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_44
timestamp -25199
transform 1 0 5152 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_48
timestamp -25199
transform 1 0 5520 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_56
timestamp -25199
transform 1 0 6256 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_64
timestamp 1636943256
transform 1 0 6992 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_76
timestamp -25199
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp -25199
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_106
timestamp 1636943256
transform 1 0 10856 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_118
timestamp -25199
transform 1 0 11960 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp -25199
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp -25199
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_150
timestamp 1636943256
transform 1 0 14904 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_162
timestamp -25199
transform 1 0 16008 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_170
timestamp -25199
transform 1 0 16744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp -25199
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_197
timestamp -25199
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_227
timestamp 1636943256
transform 1 0 21988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_239
timestamp 1636943256
transform 1 0 23092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp -25199
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1636943256
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1636943256
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1636943256
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_289
timestamp -25199
transform 1 0 27692 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp -25199
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_9
timestamp -25199
transform 1 0 1932 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_28
timestamp 1636943256
transform 1 0 3680 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_40
timestamp -25199
transform 1 0 4784 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_48
timestamp -25199
transform 1 0 5520 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp -25199
transform 1 0 6348 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_71
timestamp 1636943256
transform 1 0 7636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_83
timestamp -25199
transform 1 0 8740 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_100
timestamp 1636943256
transform 1 0 10304 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp -25199
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_128
timestamp -25199
transform 1 0 12880 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_134
timestamp -25199
transform 1 0 13432 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_155
timestamp 1636943256
transform 1 0 15364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp -25199
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1636943256
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_181
timestamp -25199
transform 1 0 17756 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_187
timestamp -25199
transform 1 0 18308 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1636943256
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1636943256
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp -25199
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp -25199
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1636943256
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1636943256
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1636943256
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1636943256
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp -25199
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp -25199
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1636943256
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_293
timestamp -25199
transform 1 0 28060 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_9
timestamp -25199
transform 1 0 1932 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636943256
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_41
timestamp -25199
transform 1 0 4876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_49
timestamp -25199
transform 1 0 5612 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_65
timestamp -25199
transform 1 0 7084 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_73
timestamp -25199
transform 1 0 7820 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp -25199
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1636943256
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1636943256
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_131
timestamp -25199
transform 1 0 13156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp -25199
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1636943256
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1636943256
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_165
timestamp -25199
transform 1 0 16284 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_171
timestamp -25199
transform 1 0 16836 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp -25199
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197
timestamp -25199
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_206
timestamp 1636943256
transform 1 0 20056 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_218
timestamp 1636943256
transform 1 0 21160 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_230
timestamp -25199
transform 1 0 22264 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_238
timestamp -25199
transform 1 0 23000 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp -25199
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_273
timestamp 1636943256
transform 1 0 26220 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_285
timestamp 1636943256
transform 1 0 27324 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_297
timestamp -25199
transform 1 0 28428 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_9
timestamp 1636943256
transform 1 0 1932 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_21
timestamp 1636943256
transform 1 0 3036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_33
timestamp 1636943256
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_45
timestamp -25199
transform 1 0 5244 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_73
timestamp 1636943256
transform 1 0 7820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_90
timestamp 1636943256
transform 1 0 9384 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_102
timestamp -25199
transform 1 0 10488 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp -25199
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1636943256
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1636943256
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1636943256
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1636943256
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp -25199
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp -25199
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp -25199
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_196
timestamp 1636943256
transform 1 0 19136 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_208
timestamp -25199
transform 1 0 20240 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_232
timestamp -25199
transform 1 0 22448 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_256
timestamp 1636943256
transform 1 0 24656 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_268
timestamp 1636943256
transform 1 0 25760 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1636943256
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_293
timestamp -25199
transform 1 0 28060 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_28_9
timestamp -25199
transform 1 0 1932 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_15
timestamp -25199
transform 1 0 2484 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_25
timestamp -25199
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636943256
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_41
timestamp -25199
transform 1 0 4876 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_49
timestamp -25199
transform 1 0 5612 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_56
timestamp -25199
transform 1 0 6256 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_60
timestamp -25199
transform 1 0 6624 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_68
timestamp 1636943256
transform 1 0 7360 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp -25199
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1636943256
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1636943256
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1636943256
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1636943256
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp -25199
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp -25199
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp -25199
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_147
timestamp -25199
transform 1 0 14628 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_166
timestamp 1636943256
transform 1 0 16376 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_178
timestamp -25199
transform 1 0 17480 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp -25199
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp -25199
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp -25199
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1636943256
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp -25199
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp -25199
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1636943256
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1636943256
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1636943256
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_289
timestamp -25199
transform 1 0 27692 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_297
timestamp -25199
transform 1 0 28428 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_9
timestamp -25199
transform 1 0 1932 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_23
timestamp -25199
transform 1 0 3220 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_34
timestamp 1636943256
transform 1 0 4232 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_46
timestamp -25199
transform 1 0 5336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp -25199
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636943256
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1636943256
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_81
timestamp -25199
transform 1 0 8556 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_98
timestamp 1636943256
transform 1 0 10120 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp -25199
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp -25199
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_117
timestamp -25199
transform 1 0 11868 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_129
timestamp 1636943256
transform 1 0 12972 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_141
timestamp -25199
transform 1 0 14076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp -25199
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1636943256
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1636943256
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1636943256
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_205
timestamp -25199
transform 1 0 19964 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_213
timestamp -25199
transform 1 0 20700 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_218
timestamp -25199
transform 1 0 21160 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1636943256
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_237
timestamp -25199
transform 1 0 22908 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_245
timestamp 1636943256
transform 1 0 23644 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_257
timestamp 1636943256
transform 1 0 24748 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp -25199
transform 1 0 25852 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_277
timestamp -25199
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1636943256
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_293
timestamp -25199
transform 1 0 28060 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_8
timestamp -25199
transform 1 0 1840 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_38
timestamp 1636943256
transform 1 0 4600 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_50
timestamp 1636943256
transform 1 0 5704 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_62
timestamp 1636943256
transform 1 0 6808 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_74
timestamp -25199
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp -25199
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1636943256
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1636943256
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_109
timestamp -25199
transform 1 0 11132 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_132
timestamp -25199
transform 1 0 13248 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp -25199
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1636943256
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1636943256
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp -25199
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp -25199
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1636943256
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1636943256
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_221
timestamp -25199
transform 1 0 21436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_232
timestamp -25199
transform 1 0 22448 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp -25199
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp -25199
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_258
timestamp 1636943256
transform 1 0 24840 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_270
timestamp 1636943256
transform 1 0 25944 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_282
timestamp 1636943256
transform 1 0 27048 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_294
timestamp -25199
transform 1 0 28152 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_298
timestamp -25199
transform 1 0 28520 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_8
timestamp -25199
transform 1 0 1840 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_15
timestamp -25199
transform 1 0 2484 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_19
timestamp -25199
transform 1 0 2852 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_31
timestamp 1636943256
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_43
timestamp -25199
transform 1 0 5060 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_57
timestamp -25199
transform 1 0 6348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_71
timestamp -25199
transform 1 0 7636 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_83
timestamp -25199
transform 1 0 8740 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_91
timestamp -25199
transform 1 0 9476 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_95
timestamp 1636943256
transform 1 0 9844 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_107
timestamp -25199
transform 1 0 10948 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp -25199
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp -25199
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_121
timestamp -25199
transform 1 0 12236 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_131
timestamp 1636943256
transform 1 0 13156 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_143
timestamp -25199
transform 1 0 14260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_151
timestamp -25199
transform 1 0 14996 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_157
timestamp -25199
transform 1 0 15548 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp -25199
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1636943256
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_181
timestamp -25199
transform 1 0 17756 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_204
timestamp 1636943256
transform 1 0 19872 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_216
timestamp -25199
transform 1 0 20976 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_225
timestamp -25199
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_233
timestamp -25199
transform 1 0 22540 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_258
timestamp 1636943256
transform 1 0 24840 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_270
timestamp -25199
transform 1 0 25944 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp -25199
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1636943256
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp -25199
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_8
timestamp -25199
transform 1 0 1840 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_16
timestamp -25199
transform 1 0 2576 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp -25199
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636943256
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1636943256
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_53
timestamp -25199
transform 1 0 5980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_60
timestamp -25199
transform 1 0 6624 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_71
timestamp 1636943256
transform 1 0 7636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp -25199
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp -25199
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_102
timestamp 1636943256
transform 1 0 10488 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_114
timestamp -25199
transform 1 0 11592 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp -25199
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1636943256
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1636943256
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1636943256
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_177
timestamp -25199
transform 1 0 17388 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1636943256
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp -25199
transform 1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_238
timestamp -25199
transform 1 0 23000 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp -25199
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp -25199
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_273
timestamp 1636943256
transform 1 0 26220 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_285
timestamp 1636943256
transform 1 0 27324 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp -25199
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_8
timestamp -25199
transform 1 0 1840 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_23
timestamp 1636943256
transform 1 0 3220 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_35
timestamp 1636943256
transform 1 0 4324 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_47
timestamp -25199
transform 1 0 5428 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp -25199
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1636943256
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1636943256
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_81
timestamp -25199
transform 1 0 8556 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_85
timestamp -25199
transform 1 0 8924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_101
timestamp -25199
transform 1 0 10396 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp -25199
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1636943256
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1636943256
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1636943256
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1636943256
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp -25199
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp -25199
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1636943256
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1636943256
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1636943256
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1636943256
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp -25199
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp -25199
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1636943256
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1636943256
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1636943256
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1636943256
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp -25199
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp -25199
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1636943256
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_293
timestamp -25199
transform 1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_13
timestamp -25199
transform 1 0 2300 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_34_25
timestamp -25199
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_38
timestamp -25199
transform 1 0 4600 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_44
timestamp -25199
transform 1 0 5152 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_48
timestamp 1636943256
transform 1 0 5520 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_60
timestamp -25199
transform 1 0 6624 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_71
timestamp 1636943256
transform 1 0 7636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp -25199
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp -25199
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_89
timestamp -25199
transform 1 0 9292 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_95
timestamp 1636943256
transform 1 0 9844 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_107
timestamp 1636943256
transform 1 0 10948 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_119
timestamp 1636943256
transform 1 0 12052 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_131
timestamp -25199
transform 1 0 13156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp -25199
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1636943256
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1636943256
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1636943256
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1636943256
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp -25199
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp -25199
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1636943256
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1636943256
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1636943256
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1636943256
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp -25199
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp -25199
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1636943256
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1636943256
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1636943256
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_289
timestamp -25199
transform 1 0 27692 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_297
timestamp -25199
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_10
timestamp -25199
transform 1 0 2024 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1636943256
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_33
timestamp -25199
transform 1 0 4140 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_39
timestamp -25199
transform 1 0 4692 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_43
timestamp -25199
transform 1 0 5060 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_51
timestamp -25199
transform 1 0 5796 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_57
timestamp -25199
transform 1 0 6348 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1636943256
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1636943256
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp -25199
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp -25199
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1636943256
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1636943256
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1636943256
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1636943256
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp -25199
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp -25199
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1636943256
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1636943256
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1636943256
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1636943256
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp -25199
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp -25199
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1636943256
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1636943256
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1636943256
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1636943256
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp -25199
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp -25199
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1636943256
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_293
timestamp -25199
transform 1 0 28060 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_9
timestamp -25199
transform 1 0 1932 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_23
timestamp -25199
transform 1 0 3220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp -25199
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_36
timestamp -25199
transform 1 0 4416 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_44
timestamp -25199
transform 1 0 5152 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_52
timestamp -25199
transform 1 0 5888 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_67
timestamp 1636943256
transform 1 0 7268 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_79
timestamp -25199
transform 1 0 8372 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp -25199
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_93
timestamp 1636943256
transform 1 0 9660 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_105
timestamp 1636943256
transform 1 0 10764 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_117
timestamp 1636943256
transform 1 0 11868 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_129
timestamp -25199
transform 1 0 12972 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_137
timestamp -25199
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1636943256
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1636943256
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1636943256
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1636943256
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp -25199
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp -25199
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1636943256
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1636943256
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1636943256
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1636943256
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp -25199
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp -25199
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1636943256
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1636943256
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1636943256
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_289
timestamp -25199
transform 1 0 27692 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_297
timestamp -25199
transform 1 0 28428 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_29
timestamp 1636943256
transform 1 0 3772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_41
timestamp 1636943256
transform 1 0 4876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp -25199
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1636943256
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_69
timestamp -25199
transform 1 0 7452 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_75
timestamp 1636943256
transform 1 0 8004 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_87
timestamp 1636943256
transform 1 0 9108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_99
timestamp 1636943256
transform 1 0 10212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp -25199
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1636943256
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1636943256
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1636943256
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1636943256
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp -25199
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp -25199
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1636943256
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1636943256
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1636943256
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1636943256
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp -25199
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp -25199
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1636943256
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1636943256
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1636943256
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1636943256
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp -25199
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp -25199
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1636943256
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_13
timestamp -25199
transform 1 0 2300 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_35
timestamp -25199
transform 1 0 4324 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_40
timestamp 1636943256
transform 1 0 4784 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_52
timestamp -25199
transform 1 0 5888 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_60
timestamp -25199
transform 1 0 6624 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp -25199
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1636943256
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1636943256
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1636943256
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1636943256
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp -25199
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp -25199
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1636943256
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1636943256
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1636943256
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1636943256
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp -25199
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp -25199
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1636943256
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1636943256
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1636943256
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1636943256
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp -25199
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp -25199
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1636943256
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1636943256
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1636943256
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_289
timestamp -25199
transform 1 0 27692 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_297
timestamp -25199
transform 1 0 28428 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_11
timestamp -25199
transform 1 0 2116 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_27
timestamp -25199
transform 1 0 3588 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_33
timestamp -25199
transform 1 0 4140 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_37
timestamp 1636943256
transform 1 0 4508 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_49
timestamp -25199
transform 1 0 5612 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp -25199
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp -25199
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_70
timestamp -25199
transform 1 0 7544 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_84
timestamp 1636943256
transform 1 0 8832 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_96
timestamp 1636943256
transform 1 0 9936 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp -25199
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1636943256
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1636943256
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1636943256
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1636943256
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp -25199
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp -25199
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1636943256
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1636943256
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1636943256
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1636943256
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp -25199
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp -25199
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1636943256
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1636943256
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1636943256
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1636943256
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp -25199
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp -25199
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1636943256
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_293
timestamp -25199
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_8
timestamp 1636943256
transform 1 0 1840 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp -25199
transform 1 0 2944 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636943256
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1636943256
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_53
timestamp -25199
transform 1 0 5980 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_61
timestamp -25199
transform 1 0 6716 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_69
timestamp 1636943256
transform 1 0 7452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_81
timestamp -25199
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1636943256
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1636943256
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1636943256
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1636943256
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp -25199
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp -25199
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1636943256
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1636943256
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1636943256
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1636943256
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp -25199
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp -25199
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1636943256
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1636943256
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1636943256
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1636943256
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp -25199
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp -25199
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1636943256
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1636943256
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1636943256
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_289
timestamp -25199
transform 1 0 27692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_297
timestamp -25199
transform 1 0 28428 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_9
timestamp 1636943256
transform 1 0 1932 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_21
timestamp 1636943256
transform 1 0 3036 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_33
timestamp 1636943256
transform 1 0 4140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_45
timestamp -25199
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp -25199
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1636943256
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1636943256
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1636943256
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1636943256
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp -25199
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp -25199
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1636943256
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1636943256
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1636943256
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1636943256
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp -25199
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp -25199
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1636943256
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1636943256
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1636943256
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1636943256
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp -25199
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp -25199
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1636943256
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1636943256
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1636943256
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1636943256
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp -25199
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp -25199
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1636943256
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp -25199
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_9
timestamp 1636943256
transform 1 0 1932 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp -25199
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp -25199
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636943256
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1636943256
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1636943256
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1636943256
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp -25199
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp -25199
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1636943256
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1636943256
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1636943256
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1636943256
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp -25199
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp -25199
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1636943256
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1636943256
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1636943256
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1636943256
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp -25199
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp -25199
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1636943256
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1636943256
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1636943256
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1636943256
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp -25199
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp -25199
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1636943256
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1636943256
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1636943256
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_289
timestamp -25199
transform 1 0 27692 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_297
timestamp -25199
transform 1 0 28428 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636943256
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636943256
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1636943256
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1636943256
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp -25199
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp -25199
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1636943256
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1636943256
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1636943256
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1636943256
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp -25199
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp -25199
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1636943256
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1636943256
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1636943256
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1636943256
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp -25199
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp -25199
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1636943256
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1636943256
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1636943256
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1636943256
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp -25199
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp -25199
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1636943256
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1636943256
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1636943256
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1636943256
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp -25199
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp -25199
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1636943256
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_293
timestamp -25199
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1636943256
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1636943256
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp -25199
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1636943256
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1636943256
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1636943256
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1636943256
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp -25199
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp -25199
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1636943256
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1636943256
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1636943256
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1636943256
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp -25199
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp -25199
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1636943256
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1636943256
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1636943256
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1636943256
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp -25199
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp -25199
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1636943256
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1636943256
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1636943256
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1636943256
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp -25199
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp -25199
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1636943256
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1636943256
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1636943256
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_289
timestamp -25199
transform 1 0 27692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_297
timestamp -25199
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1636943256
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1636943256
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1636943256
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1636943256
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp -25199
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp -25199
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1636943256
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1636943256
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1636943256
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1636943256
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp -25199
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp -25199
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1636943256
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1636943256
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1636943256
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1636943256
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp -25199
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp -25199
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1636943256
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1636943256
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1636943256
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1636943256
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp -25199
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp -25199
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1636943256
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1636943256
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1636943256
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1636943256
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp -25199
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp -25199
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1636943256
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_293
timestamp -25199
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636943256
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636943256
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp -25199
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1636943256
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1636943256
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_53
timestamp -25199
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_57
timestamp 1636943256
transform 1 0 6348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_69
timestamp 1636943256
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp -25199
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1636943256
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1636943256
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_109
timestamp -25199
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_113
timestamp 1636943256
transform 1 0 11500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_125
timestamp 1636943256
transform 1 0 12604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp -25199
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1636943256
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1636943256
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_165
timestamp -25199
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_169
timestamp 1636943256
transform 1 0 16652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_181
timestamp 1636943256
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_193
timestamp -25199
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1636943256
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1636943256
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_221
timestamp -25199
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_225
timestamp 1636943256
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_237
timestamp 1636943256
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp -25199
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1636943256
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1636943256
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_277
timestamp -25199
transform 1 0 26588 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_281
timestamp 1636943256
transform 1 0 26956 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_293
timestamp -25199
transform 1 0 28060 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp -25199
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp -25199
transform -1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp -25199
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp -25199
transform -1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp -25199
transform 1 0 1380 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp -25199
transform 1 0 1380 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input7
timestamp -25199
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp -25199
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp -25199
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp -25199
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp -25199
transform -1 0 2300 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp -25199
transform -1 0 2300 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input13
timestamp -25199
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp -25199
transform 1 0 1380 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp -25199
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input16
timestamp -25199
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp -25199
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp -25199
transform 1 0 1380 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp -25199
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp -25199
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp -25199
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp -25199
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp -25199
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input24
timestamp -25199
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp -25199
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp -25199
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp -25199
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp -25199
transform 1 0 1380 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input29
timestamp -25199
transform 1 0 1380 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp -25199
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp -25199
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp -25199
transform 1 0 1380 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp -25199
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input34
timestamp -25199
transform 1 0 1380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp -25199
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp -25199
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp -25199
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp -25199
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  output39
timestamp -25199
transform 1 0 28060 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output40
timestamp -25199
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_47
timestamp -25199
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -25199
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_48
timestamp -25199
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -25199
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_49
timestamp -25199
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -25199
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_50
timestamp -25199
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -25199
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_51
timestamp -25199
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -25199
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_52
timestamp -25199
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -25199
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_53
timestamp -25199
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -25199
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_54
timestamp -25199
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -25199
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_55
timestamp -25199
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -25199
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_56
timestamp -25199
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -25199
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_57
timestamp -25199
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -25199
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_58
timestamp -25199
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -25199
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_59
timestamp -25199
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -25199
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_60
timestamp -25199
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -25199
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_61
timestamp -25199
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -25199
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_62
timestamp -25199
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -25199
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_63
timestamp -25199
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -25199
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_64
timestamp -25199
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -25199
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_65
timestamp -25199
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -25199
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_66
timestamp -25199
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -25199
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_67
timestamp -25199
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -25199
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_68
timestamp -25199
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -25199
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_69
timestamp -25199
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -25199
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_70
timestamp -25199
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -25199
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_71
timestamp -25199
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -25199
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_72
timestamp -25199
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp -25199
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_73
timestamp -25199
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp -25199
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_74
timestamp -25199
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp -25199
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_75
timestamp -25199
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp -25199
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_76
timestamp -25199
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp -25199
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_77
timestamp -25199
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp -25199
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_78
timestamp -25199
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp -25199
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_79
timestamp -25199
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp -25199
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_80
timestamp -25199
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp -25199
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_81
timestamp -25199
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp -25199
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_82
timestamp -25199
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp -25199
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_83
timestamp -25199
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp -25199
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_84
timestamp -25199
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp -25199
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_85
timestamp -25199
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp -25199
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_86
timestamp -25199
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp -25199
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_87
timestamp -25199
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp -25199
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_88
timestamp -25199
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp -25199
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_89
timestamp -25199
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp -25199
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_90
timestamp -25199
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp -25199
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_91
timestamp -25199
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp -25199
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_92
timestamp -25199
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp -25199
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_93
timestamp -25199
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp -25199
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_94
timestamp -25199
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_95
timestamp -25199
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_96
timestamp -25199
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_97
timestamp -25199
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_98
timestamp -25199
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_99
timestamp -25199
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_100
timestamp -25199
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_101
timestamp -25199
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_102
timestamp -25199
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_103
timestamp -25199
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_104
timestamp -25199
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_105
timestamp -25199
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_106
timestamp -25199
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_107
timestamp -25199
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_108
timestamp -25199
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_109
timestamp -25199
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_110
timestamp -25199
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_111
timestamp -25199
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_112
timestamp -25199
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_113
timestamp -25199
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_114
timestamp -25199
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_115
timestamp -25199
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_116
timestamp -25199
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_117
timestamp -25199
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_118
timestamp -25199
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_119
timestamp -25199
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_120
timestamp -25199
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_121
timestamp -25199
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_122
timestamp -25199
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_123
timestamp -25199
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_124
timestamp -25199
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_125
timestamp -25199
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_126
timestamp -25199
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_127
timestamp -25199
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_128
timestamp -25199
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_129
timestamp -25199
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_130
timestamp -25199
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_131
timestamp -25199
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_132
timestamp -25199
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_133
timestamp -25199
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_134
timestamp -25199
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_135
timestamp -25199
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_136
timestamp -25199
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_137
timestamp -25199
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_138
timestamp -25199
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_139
timestamp -25199
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_140
timestamp -25199
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_141
timestamp -25199
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_142
timestamp -25199
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_143
timestamp -25199
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_144
timestamp -25199
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_145
timestamp -25199
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_146
timestamp -25199
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_147
timestamp -25199
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_148
timestamp -25199
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_149
timestamp -25199
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_150
timestamp -25199
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_151
timestamp -25199
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_152
timestamp -25199
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_153
timestamp -25199
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_154
timestamp -25199
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_155
timestamp -25199
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_156
timestamp -25199
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_157
timestamp -25199
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_158
timestamp -25199
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_159
timestamp -25199
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_160
timestamp -25199
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_161
timestamp -25199
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_162
timestamp -25199
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_163
timestamp -25199
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_164
timestamp -25199
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_165
timestamp -25199
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_166
timestamp -25199
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_167
timestamp -25199
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_168
timestamp -25199
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_169
timestamp -25199
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_170
timestamp -25199
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_171
timestamp -25199
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_172
timestamp -25199
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_173
timestamp -25199
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_174
timestamp -25199
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_175
timestamp -25199
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_176
timestamp -25199
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_177
timestamp -25199
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_178
timestamp -25199
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_179
timestamp -25199
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_180
timestamp -25199
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_181
timestamp -25199
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_182
timestamp -25199
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_183
timestamp -25199
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_184
timestamp -25199
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_185
timestamp -25199
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_186
timestamp -25199
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_187
timestamp -25199
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_188
timestamp -25199
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_189
timestamp -25199
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_190
timestamp -25199
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_191
timestamp -25199
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_192
timestamp -25199
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_193
timestamp -25199
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_194
timestamp -25199
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_195
timestamp -25199
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_196
timestamp -25199
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_197
timestamp -25199
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_198
timestamp -25199
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_199
timestamp -25199
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_200
timestamp -25199
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_201
timestamp -25199
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_202
timestamp -25199
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_203
timestamp -25199
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_204
timestamp -25199
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_205
timestamp -25199
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_206
timestamp -25199
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_207
timestamp -25199
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_208
timestamp -25199
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_209
timestamp -25199
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_210
timestamp -25199
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_211
timestamp -25199
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_212
timestamp -25199
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_213
timestamp -25199
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_214
timestamp -25199
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_215
timestamp -25199
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_216
timestamp -25199
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_217
timestamp -25199
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_218
timestamp -25199
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_219
timestamp -25199
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_220
timestamp -25199
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_221
timestamp -25199
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_222
timestamp -25199
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_223
timestamp -25199
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_224
timestamp -25199
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_225
timestamp -25199
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_226
timestamp -25199
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_227
timestamp -25199
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_228
timestamp -25199
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_229
timestamp -25199
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_230
timestamp -25199
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_231
timestamp -25199
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_232
timestamp -25199
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_233
timestamp -25199
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_234
timestamp -25199
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_235
timestamp -25199
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_236
timestamp -25199
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_237
timestamp -25199
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_238
timestamp -25199
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_239
timestamp -25199
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_240
timestamp -25199
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_241
timestamp -25199
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_242
timestamp -25199
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_243
timestamp -25199
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_244
timestamp -25199
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_245
timestamp -25199
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_246
timestamp -25199
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_247
timestamp -25199
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_248
timestamp -25199
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_249
timestamp -25199
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_250
timestamp -25199
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_251
timestamp -25199
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_252
timestamp -25199
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp -25199
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_254
timestamp -25199
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_255
timestamp -25199
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_256
timestamp -25199
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_257
timestamp -25199
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp -25199
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_259
timestamp -25199
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_260
timestamp -25199
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_261
timestamp -25199
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_262
timestamp -25199
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp -25199
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_264
timestamp -25199
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp -25199
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_266
timestamp -25199
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_267
timestamp -25199
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp -25199
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_269
timestamp -25199
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_270
timestamp -25199
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_271
timestamp -25199
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_272
timestamp -25199
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp -25199
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_274
timestamp -25199
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_275
timestamp -25199
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_276
timestamp -25199
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_277
timestamp -25199
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp -25199
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_279
timestamp -25199
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_280
timestamp -25199
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_281
timestamp -25199
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_282
timestamp -25199
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp -25199
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_284
timestamp -25199
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_285
timestamp -25199
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_286
timestamp -25199
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_287
timestamp -25199
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp -25199
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_289
timestamp -25199
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_290
timestamp -25199
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_291
timestamp -25199
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_292
timestamp -25199
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp -25199
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_294
timestamp -25199
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_295
timestamp -25199
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_296
timestamp -25199
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_297
timestamp -25199
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_298
timestamp -25199
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_299
timestamp -25199
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_300
timestamp -25199
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_301
timestamp -25199
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_302
timestamp -25199
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_303
timestamp -25199
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_304
timestamp -25199
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_305
timestamp -25199
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_306
timestamp -25199
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_307
timestamp -25199
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_308
timestamp -25199
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_309
timestamp -25199
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_310
timestamp -25199
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_311
timestamp -25199
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_312
timestamp -25199
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_313
timestamp -25199
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_314
timestamp -25199
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_315
timestamp -25199
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_316
timestamp -25199
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_317
timestamp -25199
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_318
timestamp -25199
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_319
timestamp -25199
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_320
timestamp -25199
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_321
timestamp -25199
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_322
timestamp -25199
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_323
timestamp -25199
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_324
timestamp -25199
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_325
timestamp -25199
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_326
timestamp -25199
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_327
timestamp -25199
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_328
timestamp -25199
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_329
timestamp -25199
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_330
timestamp -25199
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_331
timestamp -25199
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_332
timestamp -25199
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_333
timestamp -25199
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_334
timestamp -25199
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_335
timestamp -25199
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_336
timestamp -25199
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_337
timestamp -25199
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_338
timestamp -25199
transform 1 0 26864 0 1 27200
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 dec_bits_i[0]
port 1 nsew signal input
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 dec_bits_i[1]
port 2 nsew signal input
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 dec_bits_i[2]
port 3 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 dec_bits_i[3]
port 4 nsew signal input
flabel metal3 s 29200 7352 30000 7472 0 FreeSans 480 0 0 0 decoded_bit_o
port 5 nsew signal output
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 pm_new_s0_i[0]
port 6 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 pm_new_s0_i[1]
port 7 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 pm_new_s0_i[2]
port 8 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 pm_new_s0_i[3]
port 9 nsew signal input
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 pm_new_s0_i[4]
port 10 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 pm_new_s0_i[5]
port 11 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 pm_new_s0_i[6]
port 12 nsew signal input
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 pm_new_s0_i[7]
port 13 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 pm_new_s1_i[0]
port 14 nsew signal input
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 pm_new_s1_i[1]
port 15 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 pm_new_s1_i[2]
port 16 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 pm_new_s1_i[3]
port 17 nsew signal input
flabel metal3 s 0 14696 800 14816 0 FreeSans 480 0 0 0 pm_new_s1_i[4]
port 18 nsew signal input
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 pm_new_s1_i[5]
port 19 nsew signal input
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 pm_new_s1_i[6]
port 20 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 pm_new_s1_i[7]
port 21 nsew signal input
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 pm_new_s2_i[0]
port 22 nsew signal input
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 pm_new_s2_i[1]
port 23 nsew signal input
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 pm_new_s2_i[2]
port 24 nsew signal input
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 pm_new_s2_i[3]
port 25 nsew signal input
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 pm_new_s2_i[4]
port 26 nsew signal input
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 pm_new_s2_i[5]
port 27 nsew signal input
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 pm_new_s2_i[6]
port 28 nsew signal input
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 pm_new_s2_i[7]
port 29 nsew signal input
flabel metal3 s 0 21224 800 21344 0 FreeSans 480 0 0 0 pm_new_s3_i[0]
port 30 nsew signal input
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 pm_new_s3_i[1]
port 31 nsew signal input
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 pm_new_s3_i[2]
port 32 nsew signal input
flabel metal3 s 0 22856 800 22976 0 FreeSans 480 0 0 0 pm_new_s3_i[3]
port 33 nsew signal input
flabel metal3 s 0 23400 800 23520 0 FreeSans 480 0 0 0 pm_new_s3_i[4]
port 34 nsew signal input
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 pm_new_s3_i[5]
port 35 nsew signal input
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 pm_new_s3_i[6]
port 36 nsew signal input
flabel metal3 s 0 25032 800 25152 0 FreeSans 480 0 0 0 pm_new_s3_i[7]
port 37 nsew signal input
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 rst_n
port 38 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 valid_i
port 39 nsew signal input
flabel metal3 s 29200 22312 30000 22432 0 FreeSans 480 0 0 0 valid_o
port 40 nsew signal output
flabel metal4 s 2904 2128 3304 27792 0 FreeSans 1920 90 0 0 vccd1
port 41 nsew power bidirectional
flabel metal4 s 10904 2128 11304 27792 0 FreeSans 1920 90 0 0 vccd1
port 41 nsew power bidirectional
flabel metal4 s 18904 2128 19304 27792 0 FreeSans 1920 90 0 0 vccd1
port 41 nsew power bidirectional
flabel metal4 s 26904 2128 27304 27792 0 FreeSans 1920 90 0 0 vccd1
port 41 nsew power bidirectional
flabel metal4 s 3644 2128 4044 27792 0 FreeSans 1920 90 0 0 vssd1
port 42 nsew ground bidirectional
flabel metal4 s 11644 2128 12044 27792 0 FreeSans 1920 90 0 0 vssd1
port 42 nsew ground bidirectional
flabel metal4 s 19644 2128 20044 27792 0 FreeSans 1920 90 0 0 vssd1
port 42 nsew ground bidirectional
flabel metal4 s 27644 2128 28044 27792 0 FreeSans 1920 90 0 0 vssd1
port 42 nsew ground bidirectional
rlabel metal1 14996 27744 14996 27744 0 vccd1
rlabel metal1 14996 27200 14996 27200 0 vssd1
rlabel metal1 24104 19754 24104 19754 0 _000_
rlabel metal2 23138 17646 23138 17646 0 _001_
rlabel metal2 18170 19550 18170 19550 0 _002_
rlabel metal2 17986 14382 17986 14382 0 _003_
rlabel metal2 22126 11288 22126 11288 0 _004_
rlabel metal2 22126 8942 22126 8942 0 _005_
rlabel metal1 22172 6970 22172 6970 0 _006_
rlabel metal1 21528 5338 21528 5338 0 _007_
rlabel metal2 15686 4318 15686 4318 0 _008_
rlabel metal2 11914 3740 11914 3740 0 _009_
rlabel metal1 7360 4250 7360 4250 0 _010_
rlabel metal1 2162 4250 2162 4250 0 _011_
rlabel metal2 7130 10404 7130 10404 0 _012_
rlabel metal1 11730 10234 11730 10234 0 _013_
rlabel metal1 14950 15674 14950 15674 0 _014_
rlabel metal1 14628 17850 14628 17850 0 _015_
rlabel metal1 21666 14280 21666 14280 0 _016_
rlabel metal1 24334 13498 24334 13498 0 _017_
rlabel metal2 24702 8092 24702 8092 0 _018_
rlabel metal2 25162 4964 25162 4964 0 _019_
rlabel metal1 19826 3162 19826 3162 0 _020_
rlabel metal2 17894 3298 17894 3298 0 _021_
rlabel metal1 11224 3094 11224 3094 0 _022_
rlabel metal1 4278 3162 4278 3162 0 _023_
rlabel metal1 4738 6970 4738 6970 0 _024_
rlabel metal2 10258 8738 10258 8738 0 _025_
rlabel metal2 14398 9180 14398 9180 0 _026_
rlabel metal2 15318 12002 15318 12002 0 _027_
rlabel metal1 16146 17850 16146 17850 0 _028_
rlabel metal1 18124 17102 18124 17102 0 _029_
rlabel metal1 17473 16762 17473 16762 0 _030_
rlabel metal1 19274 14484 19274 14484 0 _031_
rlabel metal2 17618 11356 17618 11356 0 _032_
rlabel metal2 18170 9758 18170 9758 0 _033_
rlabel metal2 19550 8194 19550 8194 0 _034_
rlabel metal1 16882 7514 16882 7514 0 _035_
rlabel metal2 14398 6562 14398 6562 0 _036_
rlabel metal2 12834 6290 12834 6290 0 _037_
rlabel metal2 10350 6426 10350 6426 0 _038_
rlabel metal1 3450 7276 3450 7276 0 _039_
rlabel metal1 7084 9690 7084 9690 0 _040_
rlabel metal2 9706 11220 9706 11220 0 _041_
rlabel metal1 11960 12886 11960 12886 0 _042_
rlabel metal1 12144 18394 12144 18394 0 _043_
rlabel metal1 22126 15096 22126 15096 0 _044_
rlabel metal2 23322 11934 23322 11934 0 _045_
rlabel metal2 23690 10030 23690 10030 0 _046_
rlabel metal1 21436 3434 21436 3434 0 _047_
rlabel metal1 17848 5270 17848 5270 0 _048_
rlabel metal2 14398 4012 14398 4012 0 _049_
rlabel metal1 7222 3162 7222 3162 0 _050_
rlabel metal1 4416 4658 4416 4658 0 _051_
rlabel metal1 6992 7514 6992 7514 0 _052_
rlabel metal1 2346 8602 2346 8602 0 _053_
rlabel metal2 14122 10404 14122 10404 0 _054_
rlabel metal2 14490 13668 14490 13668 0 _055_
rlabel metal2 12098 16422 12098 16422 0 _056_
rlabel metal1 20102 17544 20102 17544 0 _057_
rlabel metal1 24610 16626 24610 16626 0 _058_
rlabel metal1 23092 19278 23092 19278 0 _059_
rlabel metal1 21613 20026 21613 20026 0 _060_
rlabel metal2 19918 16830 19918 16830 0 _061_
rlabel metal1 4370 13498 4370 13498 0 _062_
rlabel metal1 4002 11152 4002 11152 0 _063_
rlabel via2 3910 13923 3910 13923 0 _064_
rlabel metal1 2254 16048 2254 16048 0 _065_
rlabel metal1 7912 13498 7912 13498 0 _066_
rlabel metal2 2438 13260 2438 13260 0 _067_
rlabel metal1 3266 23086 3266 23086 0 _068_
rlabel metal2 4922 21794 4922 21794 0 _069_
rlabel metal1 2438 21556 2438 21556 0 _070_
rlabel metal1 5290 21930 5290 21930 0 _071_
rlabel metal2 2714 19958 2714 19958 0 _072_
rlabel metal1 5520 19142 5520 19142 0 _073_
rlabel metal1 2438 20434 2438 20434 0 _074_
rlabel metal1 5980 21998 5980 21998 0 _075_
rlabel metal1 9568 14926 9568 14926 0 _076_
rlabel metal1 5014 23154 5014 23154 0 _077_
rlabel metal1 7222 23494 7222 23494 0 _078_
rlabel metal1 6670 20026 6670 20026 0 _079_
rlabel metal1 7130 19380 7130 19380 0 _080_
rlabel metal1 5658 23562 5658 23562 0 _081_
rlabel metal1 4600 16966 4600 16966 0 _082_
rlabel metal1 7084 17102 7084 17102 0 _083_
rlabel metal1 22816 18258 22816 18258 0 _084_
rlabel metal1 9614 19380 9614 19380 0 _085_
rlabel metal2 10258 20026 10258 20026 0 _086_
rlabel metal1 9752 19482 9752 19482 0 _087_
rlabel via1 9627 19754 9627 19754 0 _088_
rlabel metal2 8234 19686 8234 19686 0 _089_
rlabel metal2 10074 20060 10074 20060 0 _090_
rlabel metal2 9430 19618 9430 19618 0 _091_
rlabel metal1 8418 19278 8418 19278 0 _092_
rlabel metal2 6210 19618 6210 19618 0 _093_
rlabel metal1 9936 18258 9936 18258 0 _094_
rlabel metal2 7130 13498 7130 13498 0 _095_
rlabel metal1 6624 13226 6624 13226 0 _096_
rlabel metal1 7084 12954 7084 12954 0 _097_
rlabel metal2 8050 14518 8050 14518 0 _098_
rlabel metal1 9430 13158 9430 13158 0 _099_
rlabel metal1 9016 13362 9016 13362 0 _100_
rlabel metal1 9430 13294 9430 13294 0 _101_
rlabel metal2 9614 14518 9614 14518 0 _102_
rlabel metal2 8970 13668 8970 13668 0 _103_
rlabel metal2 7038 13702 7038 13702 0 _104_
rlabel metal1 8464 14042 8464 14042 0 _105_
rlabel metal1 9982 18326 9982 18326 0 _106_
rlabel metal1 9706 18224 9706 18224 0 _107_
rlabel metal1 9752 15130 9752 15130 0 _108_
rlabel metal1 9476 16150 9476 16150 0 _109_
rlabel metal1 10350 15878 10350 15878 0 _110_
rlabel metal2 9614 15878 9614 15878 0 _111_
rlabel metal1 8786 16218 8786 16218 0 _112_
rlabel metal1 8004 23630 8004 23630 0 _113_
rlabel metal2 7958 22406 7958 22406 0 _114_
rlabel metal1 7912 22474 7912 22474 0 _115_
rlabel metal2 7958 23494 7958 23494 0 _116_
rlabel metal1 7774 23834 7774 23834 0 _117_
rlabel metal2 8418 23868 8418 23868 0 _118_
rlabel metal1 9016 17238 9016 17238 0 _119_
rlabel metal1 6670 15674 6670 15674 0 _120_
rlabel metal1 6586 16218 6586 16218 0 _121_
rlabel metal1 7130 15606 7130 15606 0 _122_
rlabel metal1 8216 16558 8216 16558 0 _123_
rlabel metal1 8878 22066 8878 22066 0 _124_
rlabel metal2 7130 16388 7130 16388 0 _125_
rlabel metal2 8602 19312 8602 19312 0 _126_
rlabel metal1 9568 21862 9568 21862 0 _127_
rlabel metal1 10258 15674 10258 15674 0 _128_
rlabel metal2 9890 16728 9890 16728 0 _129_
rlabel metal1 9384 17306 9384 17306 0 _130_
rlabel metal2 12466 19108 12466 19108 0 _131_
rlabel metal1 7498 21488 7498 21488 0 _132_
rlabel metal1 6486 21590 6486 21590 0 _133_
rlabel metal1 6118 21420 6118 21420 0 _134_
rlabel metal1 6532 21522 6532 21522 0 _135_
rlabel metal1 6532 21114 6532 21114 0 _136_
rlabel metal1 6578 17136 6578 17136 0 _137_
rlabel metal1 6532 16762 6532 16762 0 _138_
rlabel metal2 6394 17340 6394 17340 0 _139_
rlabel metal2 7130 17476 7130 17476 0 _140_
rlabel metal2 7774 17442 7774 17442 0 _141_
rlabel metal1 7360 17850 7360 17850 0 _142_
rlabel metal1 6670 21488 6670 21488 0 _143_
rlabel metal1 7268 20910 7268 20910 0 _144_
rlabel metal2 12926 20060 12926 20060 0 _145_
rlabel metal2 12558 19584 12558 19584 0 _146_
rlabel metal2 2622 23290 2622 23290 0 _147_
rlabel metal1 2898 22032 2898 22032 0 _148_
rlabel metal1 2944 16218 2944 16218 0 _149_
rlabel metal1 2622 15504 2622 15504 0 _150_
rlabel metal1 2530 15062 2530 15062 0 _151_
rlabel metal1 2438 15130 2438 15130 0 _152_
rlabel metal1 3174 15674 3174 15674 0 _153_
rlabel metal1 3358 16524 3358 16524 0 _154_
rlabel metal1 2622 16762 2622 16762 0 _155_
rlabel metal1 3680 22066 3680 22066 0 _156_
rlabel metal1 2484 22202 2484 22202 0 _157_
rlabel metal1 3726 20774 3726 20774 0 _158_
rlabel metal1 3818 18802 3818 18802 0 _159_
rlabel metal1 3818 18938 3818 18938 0 _160_
rlabel metal1 3818 18734 3818 18734 0 _161_
rlabel metal2 3818 18938 3818 18938 0 _162_
rlabel metal1 3128 18938 3128 18938 0 _163_
rlabel metal1 3680 19346 3680 19346 0 _164_
rlabel metal1 3956 18326 3956 18326 0 _165_
rlabel metal1 3680 17646 3680 17646 0 _166_
rlabel metal2 4094 13056 4094 13056 0 _167_
rlabel metal1 3220 12818 3220 12818 0 _168_
rlabel metal1 2530 11322 2530 11322 0 _169_
rlabel metal1 3450 11118 3450 11118 0 _170_
rlabel metal1 3726 10982 3726 10982 0 _171_
rlabel metal1 4462 10778 4462 10778 0 _172_
rlabel metal2 4370 11186 4370 11186 0 _173_
rlabel metal1 3818 13362 3818 13362 0 _174_
rlabel metal2 3450 13090 3450 13090 0 _175_
rlabel metal1 4186 13158 4186 13158 0 _176_
rlabel metal1 3818 18258 3818 18258 0 _177_
rlabel metal2 3450 17884 3450 17884 0 _178_
rlabel via2 3818 11339 3818 11339 0 _179_
rlabel metal1 3772 17850 3772 17850 0 _180_
rlabel metal1 4278 22984 4278 22984 0 _181_
rlabel metal1 3174 20944 3174 20944 0 _182_
rlabel metal1 3128 20570 3128 20570 0 _183_
rlabel metal1 3864 14042 3864 14042 0 _184_
rlabel metal2 3542 14212 3542 14212 0 _185_
rlabel metal1 4094 14348 4094 14348 0 _186_
rlabel metal2 4278 15334 4278 15334 0 _187_
rlabel metal3 2829 19924 2829 19924 0 _188_
rlabel metal1 3588 20910 3588 20910 0 _189_
rlabel metal1 3726 21114 3726 21114 0 _190_
rlabel metal1 13110 19924 13110 19924 0 _191_
rlabel metal1 13156 19754 13156 19754 0 _192_
rlabel metal1 16192 19754 16192 19754 0 _193_
rlabel metal1 19182 15062 19182 15062 0 _194_
rlabel metal2 22310 12954 22310 12954 0 _195_
rlabel metal1 22954 9690 22954 9690 0 _196_
rlabel metal1 23184 6766 23184 6766 0 _197_
rlabel metal2 21942 4964 21942 4964 0 _198_
rlabel metal2 17894 4386 17894 4386 0 _199_
rlabel metal1 12236 3706 12236 3706 0 _200_
rlabel metal1 8142 3978 8142 3978 0 _201_
rlabel metal1 3634 3978 3634 3978 0 _202_
rlabel metal1 7452 9146 7452 9146 0 _203_
rlabel metal1 12190 9690 12190 9690 0 _204_
rlabel metal1 14444 11322 14444 11322 0 _205_
rlabel metal2 16238 16082 16238 16082 0 _206_
rlabel metal1 24380 13362 24380 13362 0 _207_
rlabel metal1 24380 8602 24380 8602 0 _208_
rlabel metal1 24610 7174 24610 7174 0 _209_
rlabel metal2 22678 3536 22678 3536 0 _210_
rlabel metal2 17434 3502 17434 3502 0 _211_
rlabel metal1 11500 3162 11500 3162 0 _212_
rlabel metal1 6946 3094 6946 3094 0 _213_
rlabel metal2 5566 6256 5566 6256 0 _214_
rlabel metal1 8418 8364 8418 8364 0 _215_
rlabel metal1 13340 9146 13340 9146 0 _216_
rlabel metal1 15916 11322 15916 11322 0 _217_
rlabel metal1 16008 14586 16008 14586 0 _218_
rlabel metal1 18768 11866 18768 11866 0 _219_
rlabel metal1 19642 10098 19642 10098 0 _220_
rlabel metal1 20194 7718 20194 7718 0 _221_
rlabel metal1 17802 7514 17802 7514 0 _222_
rlabel metal1 15778 6426 15778 6426 0 _223_
rlabel metal2 12742 5882 12742 5882 0 _224_
rlabel metal1 10626 6188 10626 6188 0 _225_
rlabel metal1 6808 5882 6808 5882 0 _226_
rlabel metal1 5474 8602 5474 8602 0 _227_
rlabel metal1 9430 10540 9430 10540 0 _228_
rlabel metal1 12696 12410 12696 12410 0 _229_
rlabel metal1 12696 15130 12696 15130 0 _230_
rlabel metal1 21160 12614 21160 12614 0 _231_
rlabel metal1 23000 10778 23000 10778 0 _232_
rlabel metal2 22310 5916 22310 5916 0 _233_
rlabel metal2 18538 6188 18538 6188 0 _234_
rlabel metal1 15410 4590 15410 4590 0 _235_
rlabel metal2 14122 4352 14122 4352 0 _236_
rlabel metal1 8050 5338 8050 5338 0 _237_
rlabel metal1 7774 6426 7774 6426 0 _238_
rlabel metal1 3772 8058 3772 8058 0 _239_
rlabel metal1 9706 9928 9706 9928 0 _240_
rlabel metal1 14398 13226 14398 13226 0 _241_
rlabel metal1 12650 15674 12650 15674 0 _242_
rlabel metal1 23306 18666 23306 18666 0 _243_
rlabel metal1 20976 17306 20976 17306 0 _244_
rlabel metal2 22770 19142 22770 19142 0 _245_
rlabel metal1 22954 19380 22954 19380 0 _246_
rlabel metal3 866 4420 866 4420 0 clk
rlabel metal1 17894 15470 17894 15470 0 clknet_0_clk
rlabel metal2 1610 8160 1610 8160 0 clknet_3_0__leaf_clk
rlabel metal2 14122 7888 14122 7888 0 clknet_3_1__leaf_clk
rlabel metal2 9430 9996 9430 9996 0 clknet_3_2__leaf_clk
rlabel metal1 13846 10710 13846 10710 0 clknet_3_3__leaf_clk
rlabel metal1 17618 9554 17618 9554 0 clknet_3_4__leaf_clk
rlabel metal1 24748 5338 24748 5338 0 clknet_3_5__leaf_clk
rlabel metal1 14214 13940 14214 13940 0 clknet_3_6__leaf_clk
rlabel metal2 23046 19618 23046 19618 0 clknet_3_7__leaf_clk
rlabel metal1 1426 6290 1426 6290 0 dec_bits_i[0]
rlabel metal1 1564 6766 1564 6766 0 dec_bits_i[1]
rlabel metal1 1380 6698 1380 6698 0 dec_bits_i[2]
rlabel metal1 1794 7854 1794 7854 0 dec_bits_i[3]
rlabel metal2 28382 7599 28382 7599 0 decoded_bit_o
rlabel metal2 6118 6970 6118 6970 0 history_s0\[10\]
rlabel metal1 11592 8806 11592 8806 0 history_s0\[11\]
rlabel metal1 15134 9554 15134 9554 0 history_s0\[12\]
rlabel metal1 16192 14246 16192 14246 0 history_s0\[13\]
rlabel metal2 14490 19380 14490 19380 0 history_s0\[14\]
rlabel metal1 22908 13906 22908 13906 0 history_s0\[2\]
rlabel metal2 24794 13566 24794 13566 0 history_s0\[3\]
rlabel metal1 24840 7514 24840 7514 0 history_s0\[4\]
rlabel metal2 23322 4794 23322 4794 0 history_s0\[5\]
rlabel metal1 18676 4182 18676 4182 0 history_s0\[6\]
rlabel metal2 16330 3264 16330 3264 0 history_s0\[7\]
rlabel metal2 9338 3842 9338 3842 0 history_s0\[8\]
rlabel metal1 4876 4182 4876 4182 0 history_s0\[9\]
rlabel metal1 7866 8602 7866 8602 0 history_s1\[10\]
rlabel metal2 12006 9248 12006 9248 0 history_s1\[11\]
rlabel metal1 15134 10982 15134 10982 0 history_s1\[12\]
rlabel metal2 15962 13566 15962 13566 0 history_s1\[13\]
rlabel metal1 12512 16218 12512 16218 0 history_s1\[14\]
rlabel metal2 18722 17170 18722 17170 0 history_s1\[1\]
rlabel metal1 22908 14042 22908 14042 0 history_s1\[2\]
rlabel metal1 24196 11866 24196 11866 0 history_s1\[3\]
rlabel metal1 25116 9486 25116 9486 0 history_s1\[4\]
rlabel metal1 22310 4250 22310 4250 0 history_s1\[5\]
rlabel metal1 18814 5338 18814 5338 0 history_s1\[6\]
rlabel metal1 14720 4454 14720 4454 0 history_s1\[7\]
rlabel metal2 8326 3264 8326 3264 0 history_s1\[8\]
rlabel metal1 5520 4454 5520 4454 0 history_s1\[9\]
rlabel metal2 18630 17408 18630 17408 0 history_s2\[0\]
rlabel metal1 4048 7718 4048 7718 0 history_s2\[10\]
rlabel metal2 8142 10200 8142 10200 0 history_s2\[11\]
rlabel metal2 13294 10234 13294 10234 0 history_s2\[12\]
rlabel metal2 13570 15674 13570 15674 0 history_s2\[13\]
rlabel metal2 15134 18462 15134 18462 0 history_s2\[14\]
rlabel metal1 19136 14042 19136 14042 0 history_s2\[2\]
rlabel metal1 20700 10982 20700 10982 0 history_s2\[3\]
rlabel metal1 23506 8330 23506 8330 0 history_s2\[4\]
rlabel metal1 22586 6732 22586 6732 0 history_s2\[5\]
rlabel metal1 20562 5542 20562 5542 0 history_s2\[6\]
rlabel metal1 14214 5678 14214 5678 0 history_s2\[7\]
rlabel metal1 11868 4182 11868 4182 0 history_s2\[8\]
rlabel metal1 8096 5678 8096 5678 0 history_s2\[9\]
rlabel metal1 3772 7378 3772 7378 0 history_s3\[10\]
rlabel metal2 6762 9758 6762 9758 0 history_s3\[11\]
rlabel metal1 10994 11526 10994 11526 0 history_s3\[12\]
rlabel metal1 12880 13906 12880 13906 0 history_s3\[13\]
rlabel metal1 13018 18938 13018 18938 0 history_s3\[14\]
rlabel metal1 19458 14314 19458 14314 0 history_s3\[2\]
rlabel metal1 19274 11322 19274 11322 0 history_s3\[3\]
rlabel metal1 19596 9690 19596 9690 0 history_s3\[4\]
rlabel metal1 18860 7514 18860 7514 0 history_s3\[5\]
rlabel metal1 17020 7378 17020 7378 0 history_s3\[6\]
rlabel metal2 14766 6528 14766 6528 0 history_s3\[7\]
rlabel metal1 11086 6188 11086 6188 0 history_s3\[8\]
rlabel metal1 8188 6222 8188 6222 0 history_s3\[9\]
rlabel metal1 21712 17850 21712 17850 0 latency_counter\[0\]
rlabel via1 23414 18173 23414 18173 0 latency_counter\[1\]
rlabel metal2 23414 19210 23414 19210 0 latency_counter\[2\]
rlabel metal1 22264 19686 22264 19686 0 latency_counter\[3\]
rlabel metal1 15364 14450 15364 14450 0 net1
rlabel metal1 2438 18190 2438 18190 0 net10
rlabel metal3 2047 12036 2047 12036 0 net11
rlabel metal1 2392 19754 2392 19754 0 net12
rlabel metal1 4048 13906 4048 13906 0 net13
rlabel metal2 2944 13702 2944 13702 0 net14
rlabel metal1 5980 15470 5980 15470 0 net15
rlabel metal2 2622 14722 2622 14722 0 net16
rlabel metal3 4094 19380 4094 19380 0 net17
rlabel metal1 1702 20332 1702 20332 0 net18
rlabel via2 1610 16235 1610 16235 0 net19
rlabel metal1 1978 6868 1978 6868 0 net2
rlabel metal1 1748 16694 1748 16694 0 net20
rlabel metal2 2622 16830 2622 16830 0 net21
rlabel metal1 5842 17714 5842 17714 0 net22
rlabel metal1 6804 17170 6804 17170 0 net23
rlabel metal2 6762 18156 6762 18156 0 net24
rlabel metal1 1610 19448 1610 19448 0 net25
rlabel metal1 2346 19686 2346 19686 0 net26
rlabel metal1 9821 20434 9821 20434 0 net27
rlabel metal1 1702 21012 1702 21012 0 net28
rlabel metal3 2139 20740 2139 20740 0 net29
rlabel metal1 16468 14450 16468 14450 0 net3
rlabel metal1 1748 21862 1748 21862 0 net30
rlabel metal1 1840 22406 1840 22406 0 net31
rlabel metal2 2392 20468 2392 20468 0 net32
rlabel metal1 2070 22610 2070 22610 0 net33
rlabel metal1 2346 22542 2346 22542 0 net34
rlabel metal2 2714 24140 2714 24140 0 net35
rlabel metal1 2852 23562 2852 23562 0 net36
rlabel metal1 2070 5338 2070 5338 0 net37
rlabel metal1 1610 5576 1610 5576 0 net38
rlabel metal1 28014 7854 28014 7854 0 net39
rlabel metal2 4186 8228 4186 8228 0 net4
rlabel metal2 28106 21318 28106 21318 0 net40
rlabel metal1 19412 12750 19412 12750 0 net41
rlabel metal1 13616 12274 13616 12274 0 net42
rlabel metal2 13754 6460 13754 6460 0 net43
rlabel metal2 8142 3502 8142 3502 0 net44
rlabel metal1 6578 9520 6578 9520 0 net45
rlabel metal1 11546 8398 11546 8398 0 net46
rlabel metal1 12742 18156 12742 18156 0 net47
rlabel metal2 14858 8432 14858 8432 0 net48
rlabel metal1 17940 7990 17940 7990 0 net49
rlabel metal2 4462 14178 4462 14178 0 net5
rlabel metal1 24518 4692 24518 4692 0 net50
rlabel metal1 24794 10540 24794 10540 0 net51
rlabel metal1 17894 7854 17894 7854 0 net52
rlabel metal1 14536 15538 14536 15538 0 net53
rlabel metal1 15594 17714 15594 17714 0 net54
rlabel metal1 22172 18598 22172 18598 0 net55
rlabel metal1 21942 17238 21942 17238 0 net56
rlabel metal1 12742 16116 12742 16116 0 net57
rlabel metal1 5481 4522 5481 4522 0 net58
rlabel metal1 2438 5270 2438 5270 0 net59
rlabel metal1 2300 14926 2300 14926 0 net6
rlabel metal2 12466 9826 12466 9826 0 net60
rlabel metal2 12742 14756 12742 14756 0 net61
rlabel metal2 15410 8194 15410 8194 0 net62
rlabel metal2 18078 10880 18078 10880 0 net63
rlabel metal2 21666 9248 21666 9248 0 net64
rlabel metal1 25031 9622 25031 9622 0 net65
rlabel metal2 21298 7650 21298 7650 0 net66
rlabel metal2 18722 15181 18722 15181 0 net67
rlabel metal2 18262 16830 18262 16830 0 net68
rlabel metal2 24242 18428 24242 18428 0 net69
rlabel metal1 1794 11118 1794 11118 0 net7
rlabel via1 24058 19397 24058 19397 0 net70
rlabel metal1 16376 18258 16376 18258 0 net71
rlabel metal1 14306 7174 14306 7174 0 net72
rlabel via1 2645 21998 2645 21998 0 net73
rlabel metal1 23414 4658 23414 4658 0 net74
rlabel metal1 12512 4114 12512 4114 0 net75
rlabel metal1 7176 16762 7176 16762 0 net76
rlabel metal1 20470 12750 20470 12750 0 net77
rlabel metal2 13662 14178 13662 14178 0 net78
rlabel metal1 13432 12818 13432 12818 0 net79
rlabel via1 2637 12818 2637 12818 0 net8
rlabel viali 6655 13906 6655 13906 0 net80
rlabel metal1 24058 4046 24058 4046 0 net81
rlabel metal1 17710 3366 17710 3366 0 net82
rlabel metal1 2438 18666 2438 18666 0 net9
rlabel metal2 24610 18020 24610 18020 0 pipeline_full
rlabel metal1 1380 7922 1380 7922 0 pm_new_s0_i[0]
rlabel metal1 1380 8806 1380 8806 0 pm_new_s0_i[1]
rlabel metal1 1380 9554 1380 9554 0 pm_new_s0_i[2]
rlabel metal1 1380 10030 1380 10030 0 pm_new_s0_i[3]
rlabel metal1 1380 10642 1380 10642 0 pm_new_s0_i[4]
rlabel metal2 1426 11033 1426 11033 0 pm_new_s0_i[5]
rlabel metal1 1794 11662 1794 11662 0 pm_new_s0_i[6]
rlabel metal1 1794 12206 1794 12206 0 pm_new_s0_i[7]
rlabel metal1 1380 12818 1380 12818 0 pm_new_s1_i[0]
rlabel metal1 1334 13294 1334 13294 0 pm_new_s1_i[1]
rlabel metal1 1426 13906 1426 13906 0 pm_new_s1_i[2]
rlabel metal1 1380 14382 1380 14382 0 pm_new_s1_i[3]
rlabel metal1 1426 14994 1426 14994 0 pm_new_s1_i[4]
rlabel metal2 1426 15385 1426 15385 0 pm_new_s1_i[5]
rlabel metal1 1426 16082 1426 16082 0 pm_new_s1_i[6]
rlabel metal2 1518 16439 1518 16439 0 pm_new_s1_i[7]
rlabel metal1 1426 17170 1426 17170 0 pm_new_s2_i[0]
rlabel metal1 1380 17578 1380 17578 0 pm_new_s2_i[1]
rlabel metal1 1426 18258 1426 18258 0 pm_new_s2_i[2]
rlabel metal1 1380 18734 1380 18734 0 pm_new_s2_i[3]
rlabel metal2 1426 19227 1426 19227 0 pm_new_s2_i[4]
rlabel metal1 1380 19822 1380 19822 0 pm_new_s2_i[5]
rlabel metal1 1380 20434 1380 20434 0 pm_new_s2_i[6]
rlabel metal1 1380 20910 1380 20910 0 pm_new_s2_i[7]
rlabel metal1 1380 21522 1380 21522 0 pm_new_s3_i[0]
rlabel metal1 1380 21930 1380 21930 0 pm_new_s3_i[1]
rlabel metal1 1380 22610 1380 22610 0 pm_new_s3_i[2]
rlabel metal2 1426 23001 1426 23001 0 pm_new_s3_i[3]
rlabel metal1 1426 23698 1426 23698 0 pm_new_s3_i[4]
rlabel metal1 1380 24174 1380 24174 0 pm_new_s3_i[5]
rlabel metal1 1426 24786 1426 24786 0 pm_new_s3_i[6]
rlabel metal1 1380 25194 1380 25194 0 pm_new_s3_i[7]
rlabel metal1 1380 5202 1380 5202 0 rst_n
rlabel metal1 1380 5678 1380 5678 0 valid_i
rlabel metal2 28382 22457 28382 22457 0 valid_o
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
