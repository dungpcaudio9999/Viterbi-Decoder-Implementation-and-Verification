module sipo (byte_ready_o,
    clk,
    data_serial_i,
    rst_n,
    valid_serial_i,
    data_parallel_o);
 output byte_ready_o;
 input clk;
 input data_serial_i;
 input rst_n;
 input valid_serial_i;
 output [7:0] data_parallel_o;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire \count[0] ;
 wire \count[1] ;
 wire \count[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 sky130_fd_sc_hd__and3_1 _14_ (.A(\count[0] ),
    .B(\count[1] ),
    .C(net14),
    .X(_12_));
 sky130_fd_sc_hd__and2_1 _15_ (.A(\count[2] ),
    .B(_12_),
    .X(_00_));
 sky130_fd_sc_hd__xor2_1 _16_ (.A(\count[0] ),
    .B(net14),
    .X(_01_));
 sky130_fd_sc_hd__a21oi_1 _17_ (.A1(\count[0] ),
    .A2(net14),
    .B1(\count[1] ),
    .Y(_13_));
 sky130_fd_sc_hd__nor2_1 _18_ (.A(_12_),
    .B(_13_),
    .Y(_02_));
 sky130_fd_sc_hd__xor2_1 _19_ (.A(\count[2] ),
    .B(_12_),
    .X(_03_));
 sky130_fd_sc_hd__mux2_1 _20_ (.A0(net5),
    .A1(net6),
    .S(net13),
    .X(_04_));
 sky130_fd_sc_hd__mux2_1 _21_ (.A0(net6),
    .A1(net7),
    .S(net13),
    .X(_05_));
 sky130_fd_sc_hd__mux2_1 _22_ (.A0(net7),
    .A1(net8),
    .S(net13),
    .X(_06_));
 sky130_fd_sc_hd__mux2_1 _23_ (.A0(net8),
    .A1(net9),
    .S(net13),
    .X(_07_));
 sky130_fd_sc_hd__mux2_1 _24_ (.A0(net9),
    .A1(net10),
    .S(net13),
    .X(_08_));
 sky130_fd_sc_hd__mux2_1 _25_ (.A0(net10),
    .A1(net11),
    .S(net13),
    .X(_09_));
 sky130_fd_sc_hd__mux2_1 _26_ (.A0(net11),
    .A1(net12),
    .S(net14),
    .X(_10_));
 sky130_fd_sc_hd__mux2_1 _27_ (.A0(net12),
    .A1(net1),
    .S(net14),
    .X(_11_));
 sky130_fd_sc_hd__dfrtp_1 _28_ (.CLK(clknet_1_0__leaf_clk),
    .D(_00_),
    .RESET_B(net15),
    .Q(net4));
 sky130_fd_sc_hd__dfrtp_1 _29_ (.CLK(clknet_1_0__leaf_clk),
    .D(_01_),
    .RESET_B(net16),
    .Q(\count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _30_ (.CLK(clknet_1_0__leaf_clk),
    .D(_02_),
    .RESET_B(net15),
    .Q(\count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _31_ (.CLK(clknet_1_0__leaf_clk),
    .D(_03_),
    .RESET_B(net15),
    .Q(\count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _32_ (.CLK(clknet_1_1__leaf_clk),
    .D(_04_),
    .RESET_B(net16),
    .Q(net5));
 sky130_fd_sc_hd__dfrtp_1 _33_ (.CLK(clknet_1_1__leaf_clk),
    .D(_05_),
    .RESET_B(net16),
    .Q(net6));
 sky130_fd_sc_hd__dfrtp_1 _34_ (.CLK(clknet_1_1__leaf_clk),
    .D(_06_),
    .RESET_B(net16),
    .Q(net7));
 sky130_fd_sc_hd__dfrtp_1 _35_ (.CLK(clknet_1_1__leaf_clk),
    .D(_07_),
    .RESET_B(net16),
    .Q(net8));
 sky130_fd_sc_hd__dfrtp_1 _36_ (.CLK(clknet_1_0__leaf_clk),
    .D(_08_),
    .RESET_B(net15),
    .Q(net9));
 sky130_fd_sc_hd__dfrtp_1 _37_ (.CLK(clknet_1_1__leaf_clk),
    .D(_09_),
    .RESET_B(net15),
    .Q(net10));
 sky130_fd_sc_hd__dfrtp_1 _38_ (.CLK(clknet_1_1__leaf_clk),
    .D(_10_),
    .RESET_B(net2),
    .Q(net11));
 sky130_fd_sc_hd__dfrtp_1 _39_ (.CLK(clknet_1_0__leaf_clk),
    .D(_11_),
    .RESET_B(net15),
    .Q(net12));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_37 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(data_serial_i),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(rst_n),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(valid_serial_i),
    .X(net3));
 sky130_fd_sc_hd__buf_4 output4 (.A(net4),
    .X(byte_ready_o));
 sky130_fd_sc_hd__buf_4 output5 (.A(net5),
    .X(data_parallel_o[0]));
 sky130_fd_sc_hd__buf_4 output6 (.A(net6),
    .X(data_parallel_o[1]));
 sky130_fd_sc_hd__buf_4 output7 (.A(net7),
    .X(data_parallel_o[2]));
 sky130_fd_sc_hd__buf_4 output8 (.A(net8),
    .X(data_parallel_o[3]));
 sky130_fd_sc_hd__buf_4 output9 (.A(net9),
    .X(data_parallel_o[4]));
 sky130_fd_sc_hd__buf_4 output10 (.A(net10),
    .X(data_parallel_o[5]));
 sky130_fd_sc_hd__buf_4 output11 (.A(net11),
    .X(data_parallel_o[6]));
 sky130_fd_sc_hd__buf_4 output12 (.A(net12),
    .X(data_parallel_o[7]));
 sky130_fd_sc_hd__clkbuf_2 fanout13 (.A(net14),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 fanout14 (.A(net3),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 fanout15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 fanout16 (.A(net2),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(data_serial_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(rst_n));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(valid_serial_i));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
endmodule
