module acsu (bm_s0_s0_i,
    bm_s0_s2_i,
    bm_s1_s0_i,
    bm_s1_s2_i,
    bm_s2_s1_i,
    bm_s2_s3_i,
    bm_s3_s1_i,
    bm_s3_s3_i,
    dec_bits_o,
    pm_s0_i,
    pm_s0_o,
    pm_s1_i,
    pm_s1_o,
    pm_s2_i,
    pm_s2_o,
    pm_s3_i,
    pm_s3_o);
 input [1:0] bm_s0_s0_i;
 input [1:0] bm_s0_s2_i;
 input [1:0] bm_s1_s0_i;
 input [1:0] bm_s1_s2_i;
 input [1:0] bm_s2_s1_i;
 input [1:0] bm_s2_s3_i;
 input [1:0] bm_s3_s1_i;
 input [1:0] bm_s3_s3_i;
 output [3:0] dec_bits_o;
 input [7:0] pm_s0_i;
 output [7:0] pm_s0_o;
 input [7:0] pm_s1_i;
 output [7:0] pm_s1_o;
 input [7:0] pm_s2_i;
 output [7:0] pm_s2_o;
 input [7:0] pm_s3_i;
 output [7:0] pm_s3_o;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;

 sky130_fd_sc_hd__inv_2 _227_ (.A(net103),
    .Y(_212_));
 sky130_fd_sc_hd__inv_2 _228_ (.A(net109),
    .Y(_213_));
 sky130_fd_sc_hd__inv_2 _229_ (.A(net110),
    .Y(_214_));
 sky130_fd_sc_hd__inv_2 _230_ (.A(net107),
    .Y(_215_));
 sky130_fd_sc_hd__inv_2 _231_ (.A(net21),
    .Y(_216_));
 sky130_fd_sc_hd__nand2_1 _232_ (.A(net16),
    .B(net42),
    .Y(_217_));
 sky130_fd_sc_hd__nand2_1 _233_ (.A(net15),
    .B(net41),
    .Y(_218_));
 sky130_fd_sc_hd__xnor2_2 _234_ (.A(net16),
    .B(net42),
    .Y(_219_));
 sky130_fd_sc_hd__o21ai_4 _235_ (.A1(_218_),
    .A2(_219_),
    .B1(_217_),
    .Y(_220_));
 sky130_fd_sc_hd__nand3_1 _236_ (.A(net96),
    .B(net99),
    .C(_220_),
    .Y(_221_));
 sky130_fd_sc_hd__a21o_1 _237_ (.A1(net99),
    .A2(_220_),
    .B1(net96),
    .X(_222_));
 sky130_fd_sc_hd__and2_1 _238_ (.A(_221_),
    .B(_222_),
    .X(_223_));
 sky130_fd_sc_hd__and2_1 _239_ (.A(net12),
    .B(net34),
    .X(_224_));
 sky130_fd_sc_hd__nand2_1 _240_ (.A(net11),
    .B(net33),
    .Y(_225_));
 sky130_fd_sc_hd__xor2_1 _241_ (.A(net12),
    .B(net34),
    .X(_226_));
 sky130_fd_sc_hd__a31o_1 _242_ (.A1(net11),
    .A2(net33),
    .A3(_226_),
    .B1(_224_),
    .X(_000_));
 sky130_fd_sc_hd__and3_1 _243_ (.A(net101),
    .B(net103),
    .C(_000_),
    .X(_001_));
 sky130_fd_sc_hd__a21oi_1 _244_ (.A1(net103),
    .A2(_000_),
    .B1(net101),
    .Y(_002_));
 sky130_fd_sc_hd__nor2_1 _245_ (.A(_001_),
    .B(_002_),
    .Y(_003_));
 sky130_fd_sc_hd__o211a_1 _246_ (.A1(_001_),
    .A2(_002_),
    .B1(_221_),
    .C1(_222_),
    .X(_004_));
 sky130_fd_sc_hd__xnor2_1 _247_ (.A(net99),
    .B(_220_),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _248_ (.A(_005_),
    .Y(_006_));
 sky130_fd_sc_hd__xnor2_1 _249_ (.A(_212_),
    .B(_000_),
    .Y(_007_));
 sky130_fd_sc_hd__xnor2_1 _250_ (.A(_218_),
    .B(_219_),
    .Y(_008_));
 sky130_fd_sc_hd__xor2_1 _251_ (.A(net15),
    .B(net41),
    .X(_009_));
 sky130_fd_sc_hd__xor2_1 _252_ (.A(net11),
    .B(net33),
    .X(_010_));
 sky130_fd_sc_hd__and2b_1 _253_ (.A_N(_009_),
    .B(_010_),
    .X(_011_));
 sky130_fd_sc_hd__and3b_1 _254_ (.A_N(_009_),
    .B(_010_),
    .C(_226_),
    .X(_012_));
 sky130_fd_sc_hd__xnor2_1 _255_ (.A(_225_),
    .B(_226_),
    .Y(_013_));
 sky130_fd_sc_hd__o22a_1 _256_ (.A1(_008_),
    .A2(_012_),
    .B1(_013_),
    .B2(_011_),
    .X(_014_));
 sky130_fd_sc_hd__a21oi_1 _257_ (.A1(_005_),
    .A2(_007_),
    .B1(_014_),
    .Y(_015_));
 sky130_fd_sc_hd__nor2_1 _258_ (.A(_005_),
    .B(_007_),
    .Y(_016_));
 sky130_fd_sc_hd__and4_1 _259_ (.A(net45),
    .B(net97),
    .C(net99),
    .D(_220_),
    .X(_017_));
 sky130_fd_sc_hd__nand4_2 _260_ (.A(net45),
    .B(net97),
    .C(net99),
    .D(_220_),
    .Y(_018_));
 sky130_fd_sc_hd__a31o_1 _261_ (.A1(net97),
    .A2(net99),
    .A3(_220_),
    .B1(net45),
    .X(_019_));
 sky130_fd_sc_hd__and2_1 _262_ (.A(_018_),
    .B(_019_),
    .X(_020_));
 sky130_fd_sc_hd__and4_1 _263_ (.A(net37),
    .B(net101),
    .C(net103),
    .D(_000_),
    .X(_021_));
 sky130_fd_sc_hd__a31oi_2 _264_ (.A1(net101),
    .A2(net104),
    .A3(_000_),
    .B1(net37),
    .Y(_022_));
 sky130_fd_sc_hd__nor2_1 _265_ (.A(net94),
    .B(_022_),
    .Y(_023_));
 sky130_fd_sc_hd__a211o_1 _266_ (.A1(_018_),
    .A2(_019_),
    .B1(net94),
    .C1(_022_),
    .X(_024_));
 sky130_fd_sc_hd__a211o_1 _267_ (.A1(_221_),
    .A2(_222_),
    .B1(_001_),
    .C1(_002_),
    .X(_025_));
 sky130_fd_sc_hd__o311a_1 _268_ (.A1(_004_),
    .A2(_015_),
    .A3(_016_),
    .B1(_024_),
    .C1(_025_),
    .X(_026_));
 sky130_fd_sc_hd__xor2_1 _269_ (.A(net100),
    .B(net94),
    .X(_027_));
 sky130_fd_sc_hd__xnor2_1 _270_ (.A(net38),
    .B(_021_),
    .Y(_028_));
 sky130_fd_sc_hd__xnor2_1 _271_ (.A(net95),
    .B(_018_),
    .Y(_029_));
 sky130_fd_sc_hd__o211a_1 _272_ (.A1(net94),
    .A2(_022_),
    .B1(_018_),
    .C1(_019_),
    .X(_030_));
 sky130_fd_sc_hd__a21o_1 _273_ (.A1(_028_),
    .A2(_029_),
    .B1(_030_),
    .X(_031_));
 sky130_fd_sc_hd__and3_1 _274_ (.A(net47),
    .B(net95),
    .C(_017_),
    .X(_032_));
 sky130_fd_sc_hd__a21oi_1 _275_ (.A1(net95),
    .A2(_017_),
    .B1(net47),
    .Y(_033_));
 sky130_fd_sc_hd__nor2_1 _276_ (.A(_032_),
    .B(_033_),
    .Y(_034_));
 sky130_fd_sc_hd__and3_1 _277_ (.A(net39),
    .B(net100),
    .C(net94),
    .X(_035_));
 sky130_fd_sc_hd__a21oi_1 _278_ (.A1(net100),
    .A2(net94),
    .B1(net39),
    .Y(_036_));
 sky130_fd_sc_hd__or2_1 _279_ (.A(_035_),
    .B(_036_),
    .X(_037_));
 sky130_fd_sc_hd__inv_2 _280_ (.A(_037_),
    .Y(_038_));
 sky130_fd_sc_hd__or2_1 _281_ (.A(_028_),
    .B(_029_),
    .X(_039_));
 sky130_fd_sc_hd__o221a_1 _282_ (.A1(_026_),
    .A2(_031_),
    .B1(_034_),
    .B2(_037_),
    .C1(_039_),
    .X(_040_));
 sky130_fd_sc_hd__xor2_2 _283_ (.A(net48),
    .B(_032_),
    .X(_041_));
 sky130_fd_sc_hd__inv_2 _284_ (.A(_041_),
    .Y(_042_));
 sky130_fd_sc_hd__xnor2_2 _285_ (.A(net40),
    .B(_035_),
    .Y(_043_));
 sky130_fd_sc_hd__a22o_1 _286_ (.A1(_034_),
    .A2(_037_),
    .B1(_041_),
    .B2(_043_),
    .X(_044_));
 sky130_fd_sc_hd__o22a_1 _287_ (.A1(_041_),
    .A2(_043_),
    .B1(_044_),
    .B2(_040_),
    .X(_045_));
 sky130_fd_sc_hd__inv_2 _288_ (.A(_045_),
    .Y(net52));
 sky130_fd_sc_hd__mux2_1 _289_ (.A0(_009_),
    .A1(_010_),
    .S(net91),
    .X(net77));
 sky130_fd_sc_hd__o221a_1 _290_ (.A1(_041_),
    .A2(_043_),
    .B1(_044_),
    .B2(_040_),
    .C1(_013_),
    .X(_046_));
 sky130_fd_sc_hd__o21bai_1 _291_ (.A1(_008_),
    .A2(net91),
    .B1_N(_046_),
    .Y(net78));
 sky130_fd_sc_hd__mux2_1 _292_ (.A0(_006_),
    .A1(_007_),
    .S(net91),
    .X(net79));
 sky130_fd_sc_hd__mux2_1 _293_ (.A0(_223_),
    .A1(_003_),
    .S(net91),
    .X(net80));
 sky130_fd_sc_hd__mux2_1 _294_ (.A0(_020_),
    .A1(_023_),
    .S(_045_),
    .X(net81));
 sky130_fd_sc_hd__mux2_1 _295_ (.A0(_029_),
    .A1(_027_),
    .S(net91),
    .X(net82));
 sky130_fd_sc_hd__mux2_1 _296_ (.A0(_034_),
    .A1(_038_),
    .S(net91),
    .X(net83));
 sky130_fd_sc_hd__nor2_1 _297_ (.A(_042_),
    .B(_043_),
    .Y(net84));
 sky130_fd_sc_hd__nand2_1 _298_ (.A(net111),
    .B(net3),
    .Y(_047_));
 sky130_fd_sc_hd__or2_1 _299_ (.A(net111),
    .B(net3),
    .X(_048_));
 sky130_fd_sc_hd__and2_1 _300_ (.A(_047_),
    .B(_048_),
    .X(_049_));
 sky130_fd_sc_hd__xnor2_1 _301_ (.A(net111),
    .B(net3),
    .Y(_050_));
 sky130_fd_sc_hd__and2_1 _302_ (.A(net18),
    .B(net4),
    .X(_051_));
 sky130_fd_sc_hd__xor2_2 _303_ (.A(net18),
    .B(net4),
    .X(_052_));
 sky130_fd_sc_hd__a31o_1 _304_ (.A1(net17),
    .A2(net3),
    .A3(_052_),
    .B1(_051_),
    .X(_053_));
 sky130_fd_sc_hd__xnor2_1 _305_ (.A(_214_),
    .B(_053_),
    .Y(_054_));
 sky130_fd_sc_hd__and2_1 _306_ (.A(net8),
    .B(net26),
    .X(_055_));
 sky130_fd_sc_hd__nand2_1 _307_ (.A(net7),
    .B(net25),
    .Y(_056_));
 sky130_fd_sc_hd__xor2_1 _308_ (.A(net8),
    .B(net26),
    .X(_057_));
 sky130_fd_sc_hd__a31o_2 _309_ (.A1(net7),
    .A2(net25),
    .A3(_057_),
    .B1(_055_),
    .X(_058_));
 sky130_fd_sc_hd__xnor2_1 _310_ (.A(_215_),
    .B(_058_),
    .Y(_059_));
 sky130_fd_sc_hd__xnor2_1 _311_ (.A(_056_),
    .B(_057_),
    .Y(_060_));
 sky130_fd_sc_hd__xor2_2 _312_ (.A(net7),
    .B(net25),
    .X(_061_));
 sky130_fd_sc_hd__nor2_1 _313_ (.A(_050_),
    .B(_061_),
    .Y(_062_));
 sky130_fd_sc_hd__or3b_1 _314_ (.A(_050_),
    .B(_061_),
    .C_N(_052_),
    .X(_063_));
 sky130_fd_sc_hd__xnor2_1 _315_ (.A(_047_),
    .B(_052_),
    .Y(_064_));
 sky130_fd_sc_hd__a2bb2o_1 _316_ (.A1_N(_062_),
    .A2_N(_064_),
    .B1(_063_),
    .B2(_060_),
    .X(_065_));
 sky130_fd_sc_hd__a21boi_1 _317_ (.A1(_059_),
    .A2(_065_),
    .B1_N(_054_),
    .Y(_066_));
 sky130_fd_sc_hd__and3_1 _318_ (.A(net109),
    .B(net110),
    .C(_053_),
    .X(_067_));
 sky130_fd_sc_hd__a21oi_1 _319_ (.A1(net110),
    .A2(_053_),
    .B1(net109),
    .Y(_068_));
 sky130_fd_sc_hd__nor2_1 _320_ (.A(_067_),
    .B(_068_),
    .Y(_069_));
 sky130_fd_sc_hd__nand3_1 _321_ (.A(net107),
    .B(net106),
    .C(_058_),
    .Y(_070_));
 sky130_fd_sc_hd__a21o_1 _322_ (.A1(net107),
    .A2(_058_),
    .B1(net106),
    .X(_071_));
 sky130_fd_sc_hd__and2_1 _323_ (.A(_070_),
    .B(_071_),
    .X(_072_));
 sky130_fd_sc_hd__a211oi_1 _324_ (.A1(_070_),
    .A2(_071_),
    .B1(_067_),
    .C1(_068_),
    .Y(_073_));
 sky130_fd_sc_hd__nor2_1 _325_ (.A(_059_),
    .B(_065_),
    .Y(_074_));
 sky130_fd_sc_hd__o211ai_1 _326_ (.A1(_067_),
    .A2(_068_),
    .B1(_070_),
    .C1(_071_),
    .Y(_075_));
 sky130_fd_sc_hd__and4_1 _327_ (.A(net20),
    .B(net19),
    .C(net21),
    .D(_053_),
    .X(_076_));
 sky130_fd_sc_hd__or4b_2 _328_ (.A(_213_),
    .B(_214_),
    .C(_216_),
    .D_N(_053_),
    .X(_077_));
 sky130_fd_sc_hd__a31o_1 _329_ (.A1(net20),
    .A2(net19),
    .A3(_053_),
    .B1(net21),
    .X(_078_));
 sky130_fd_sc_hd__and2_1 _330_ (.A(_077_),
    .B(_078_),
    .X(_079_));
 sky130_fd_sc_hd__and4_1 _331_ (.A(net108),
    .B(net28),
    .C(net29),
    .D(_058_),
    .X(_080_));
 sky130_fd_sc_hd__a31oi_2 _332_ (.A1(net108),
    .A2(net28),
    .A3(_058_),
    .B1(net29),
    .Y(_081_));
 sky130_fd_sc_hd__nor2_1 _333_ (.A(net93),
    .B(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__a211o_1 _334_ (.A1(_077_),
    .A2(_078_),
    .B1(net93),
    .C1(_081_),
    .X(_083_));
 sky130_fd_sc_hd__o311a_1 _335_ (.A1(_066_),
    .A2(_073_),
    .A3(_074_),
    .B1(_075_),
    .C1(_083_),
    .X(_084_));
 sky130_fd_sc_hd__xor2_1 _336_ (.A(net105),
    .B(net93),
    .X(_085_));
 sky130_fd_sc_hd__xnor2_1 _337_ (.A(net105),
    .B(net93),
    .Y(_086_));
 sky130_fd_sc_hd__xnor2_1 _338_ (.A(net22),
    .B(_077_),
    .Y(_087_));
 sky130_fd_sc_hd__o211a_1 _339_ (.A1(net93),
    .A2(_081_),
    .B1(_077_),
    .C1(_078_),
    .X(_088_));
 sky130_fd_sc_hd__a21o_1 _340_ (.A1(_086_),
    .A2(_087_),
    .B1(_088_),
    .X(_089_));
 sky130_fd_sc_hd__or2_1 _341_ (.A(_086_),
    .B(_087_),
    .X(_090_));
 sky130_fd_sc_hd__and3_1 _342_ (.A(net23),
    .B(net22),
    .C(_076_),
    .X(_091_));
 sky130_fd_sc_hd__a21oi_1 _343_ (.A1(net22),
    .A2(_076_),
    .B1(net23),
    .Y(_092_));
 sky130_fd_sc_hd__nor2_1 _344_ (.A(_091_),
    .B(_092_),
    .Y(_093_));
 sky130_fd_sc_hd__and3_1 _345_ (.A(net31),
    .B(net105),
    .C(net93),
    .X(_094_));
 sky130_fd_sc_hd__a21oi_1 _346_ (.A1(net30),
    .A2(_080_),
    .B1(net31),
    .Y(_095_));
 sky130_fd_sc_hd__or2_1 _347_ (.A(_094_),
    .B(_095_),
    .X(_096_));
 sky130_fd_sc_hd__inv_2 _348_ (.A(_096_),
    .Y(_097_));
 sky130_fd_sc_hd__o221a_1 _349_ (.A1(_084_),
    .A2(_089_),
    .B1(_093_),
    .B2(_096_),
    .C1(_090_),
    .X(_098_));
 sky130_fd_sc_hd__xnor2_1 _350_ (.A(net32),
    .B(_094_),
    .Y(_099_));
 sky130_fd_sc_hd__xor2_1 _351_ (.A(net24),
    .B(_091_),
    .X(_100_));
 sky130_fd_sc_hd__a22o_1 _352_ (.A1(_093_),
    .A2(_096_),
    .B1(_099_),
    .B2(_100_),
    .X(_101_));
 sky130_fd_sc_hd__o22a_1 _353_ (.A1(_099_),
    .A2(_100_),
    .B1(_101_),
    .B2(_098_),
    .X(net51));
 sky130_fd_sc_hd__mux2_1 _354_ (.A0(_049_),
    .A1(_061_),
    .S(net89),
    .X(net69));
 sky130_fd_sc_hd__mux2_1 _355_ (.A0(_064_),
    .A1(_060_),
    .S(net89),
    .X(net70));
 sky130_fd_sc_hd__mux2_1 _356_ (.A0(_054_),
    .A1(_059_),
    .S(net89),
    .X(net71));
 sky130_fd_sc_hd__mux2_1 _357_ (.A0(_069_),
    .A1(_072_),
    .S(net89),
    .X(net72));
 sky130_fd_sc_hd__mux2_1 _358_ (.A0(_079_),
    .A1(_082_),
    .S(net89),
    .X(net73));
 sky130_fd_sc_hd__mux2_1 _359_ (.A0(_087_),
    .A1(_085_),
    .S(net90),
    .X(net74));
 sky130_fd_sc_hd__mux2_1 _360_ (.A0(_093_),
    .A1(_097_),
    .S(net89),
    .X(net75));
 sky130_fd_sc_hd__and2b_1 _361_ (.A_N(_099_),
    .B(_100_),
    .X(net76));
 sky130_fd_sc_hd__nand2_1 _362_ (.A(net42),
    .B(net14),
    .Y(_102_));
 sky130_fd_sc_hd__xnor2_2 _363_ (.A(net42),
    .B(net14),
    .Y(_103_));
 sky130_fd_sc_hd__nand2_1 _364_ (.A(net41),
    .B(net13),
    .Y(_104_));
 sky130_fd_sc_hd__o21ai_4 _365_ (.A1(_103_),
    .A2(_104_),
    .B1(_102_),
    .Y(_105_));
 sky130_fd_sc_hd__xor2_1 _366_ (.A(net98),
    .B(_105_),
    .X(_106_));
 sky130_fd_sc_hd__xnor2_1 _367_ (.A(net98),
    .B(_105_),
    .Y(_107_));
 sky130_fd_sc_hd__and2_1 _368_ (.A(net34),
    .B(net10),
    .X(_108_));
 sky130_fd_sc_hd__xor2_1 _369_ (.A(net34),
    .B(net10),
    .X(_109_));
 sky130_fd_sc_hd__nand2_1 _370_ (.A(net33),
    .B(net9),
    .Y(_110_));
 sky130_fd_sc_hd__a31o_2 _371_ (.A1(net33),
    .A2(net9),
    .A3(_109_),
    .B1(_108_),
    .X(_111_));
 sky130_fd_sc_hd__xnor2_1 _372_ (.A(_212_),
    .B(_111_),
    .Y(_112_));
 sky130_fd_sc_hd__xnor2_1 _373_ (.A(_109_),
    .B(_110_),
    .Y(_113_));
 sky130_fd_sc_hd__xnor2_1 _374_ (.A(_103_),
    .B(_104_),
    .Y(_114_));
 sky130_fd_sc_hd__inv_2 _375_ (.A(_114_),
    .Y(_115_));
 sky130_fd_sc_hd__or2_1 _376_ (.A(_113_),
    .B(_114_),
    .X(_116_));
 sky130_fd_sc_hd__xor2_1 _377_ (.A(net41),
    .B(net13),
    .X(_117_));
 sky130_fd_sc_hd__xor2_1 _378_ (.A(net33),
    .B(net9),
    .X(_118_));
 sky130_fd_sc_hd__and2b_1 _379_ (.A_N(_117_),
    .B(_118_),
    .X(_119_));
 sky130_fd_sc_hd__a21o_1 _380_ (.A1(_113_),
    .A2(_114_),
    .B1(_119_),
    .X(_120_));
 sky130_fd_sc_hd__a22o_1 _381_ (.A1(_107_),
    .A2(_112_),
    .B1(_116_),
    .B2(_120_),
    .X(_121_));
 sky130_fd_sc_hd__nand3_1 _382_ (.A(net101),
    .B(net103),
    .C(_111_),
    .Y(_122_));
 sky130_fd_sc_hd__a21o_1 _383_ (.A1(net103),
    .A2(_111_),
    .B1(net101),
    .X(_123_));
 sky130_fd_sc_hd__and2_1 _384_ (.A(_122_),
    .B(_123_),
    .X(_124_));
 sky130_fd_sc_hd__and3_1 _385_ (.A(net96),
    .B(net98),
    .C(_105_),
    .X(_125_));
 sky130_fd_sc_hd__a21oi_1 _386_ (.A1(net98),
    .A2(_105_),
    .B1(net96),
    .Y(_126_));
 sky130_fd_sc_hd__nor2_1 _387_ (.A(_125_),
    .B(_126_),
    .Y(_127_));
 sky130_fd_sc_hd__a211o_1 _388_ (.A1(_122_),
    .A2(_123_),
    .B1(_125_),
    .C1(_126_),
    .X(_128_));
 sky130_fd_sc_hd__or2_1 _389_ (.A(_107_),
    .B(_112_),
    .X(_129_));
 sky130_fd_sc_hd__and4_1 _390_ (.A(net45),
    .B(net96),
    .C(net98),
    .D(_105_),
    .X(_130_));
 sky130_fd_sc_hd__a31oi_2 _391_ (.A1(net96),
    .A2(net98),
    .A3(_105_),
    .B1(net45),
    .Y(_131_));
 sky130_fd_sc_hd__nor2_1 _392_ (.A(net92),
    .B(_131_),
    .Y(_132_));
 sky130_fd_sc_hd__and4_1 _393_ (.A(net37),
    .B(net102),
    .C(net104),
    .D(_111_),
    .X(_133_));
 sky130_fd_sc_hd__nand4_2 _394_ (.A(net37),
    .B(net102),
    .C(net104),
    .D(_111_),
    .Y(_134_));
 sky130_fd_sc_hd__a31o_1 _395_ (.A1(net102),
    .A2(net104),
    .A3(_111_),
    .B1(net37),
    .X(_135_));
 sky130_fd_sc_hd__and2_1 _396_ (.A(_134_),
    .B(_135_),
    .X(_136_));
 sky130_fd_sc_hd__o211a_1 _397_ (.A1(net92),
    .A2(_131_),
    .B1(_134_),
    .C1(_135_),
    .X(_137_));
 sky130_fd_sc_hd__o211a_1 _398_ (.A1(_125_),
    .A2(_126_),
    .B1(_122_),
    .C1(_123_),
    .X(_138_));
 sky130_fd_sc_hd__a311o_1 _399_ (.A1(_121_),
    .A2(_128_),
    .A3(_129_),
    .B1(_137_),
    .C1(_138_),
    .X(_139_));
 sky130_fd_sc_hd__xnor2_1 _400_ (.A(net100),
    .B(_134_),
    .Y(_140_));
 sky130_fd_sc_hd__xor2_1 _401_ (.A(net95),
    .B(net92),
    .X(_141_));
 sky130_fd_sc_hd__xnor2_1 _402_ (.A(net95),
    .B(net92),
    .Y(_142_));
 sky130_fd_sc_hd__o32a_1 _403_ (.A1(net92),
    .A2(_131_),
    .A3(_136_),
    .B1(_140_),
    .B2(_142_),
    .X(_143_));
 sky130_fd_sc_hd__and3_1 _404_ (.A(net47),
    .B(net46),
    .C(net92),
    .X(_144_));
 sky130_fd_sc_hd__a21oi_1 _405_ (.A1(net95),
    .A2(_130_),
    .B1(net47),
    .Y(_145_));
 sky130_fd_sc_hd__or2_1 _406_ (.A(_144_),
    .B(_145_),
    .X(_146_));
 sky130_fd_sc_hd__inv_2 _407_ (.A(_146_),
    .Y(_147_));
 sky130_fd_sc_hd__and3_1 _408_ (.A(net39),
    .B(net100),
    .C(_133_),
    .X(_148_));
 sky130_fd_sc_hd__a21oi_1 _409_ (.A1(net100),
    .A2(_133_),
    .B1(net39),
    .Y(_149_));
 sky130_fd_sc_hd__nor2_1 _410_ (.A(_148_),
    .B(_149_),
    .Y(_150_));
 sky130_fd_sc_hd__and2_1 _411_ (.A(_140_),
    .B(_142_),
    .X(_151_));
 sky130_fd_sc_hd__a221o_1 _412_ (.A1(_139_),
    .A2(_143_),
    .B1(_146_),
    .B2(_150_),
    .C1(_151_),
    .X(_152_));
 sky130_fd_sc_hd__xnor2_1 _413_ (.A(net48),
    .B(_144_),
    .Y(_153_));
 sky130_fd_sc_hd__xor2_1 _414_ (.A(net40),
    .B(_148_),
    .X(_154_));
 sky130_fd_sc_hd__o22a_1 _415_ (.A1(_146_),
    .A2(_150_),
    .B1(_153_),
    .B2(_154_),
    .X(_155_));
 sky130_fd_sc_hd__a22o_1 _416_ (.A1(_153_),
    .A2(_154_),
    .B1(_155_),
    .B2(_152_),
    .X(net50));
 sky130_fd_sc_hd__mux2_1 _417_ (.A0(_118_),
    .A1(_117_),
    .S(net87),
    .X(net61));
 sky130_fd_sc_hd__mux2_1 _418_ (.A0(_113_),
    .A1(_115_),
    .S(net87),
    .X(net62));
 sky130_fd_sc_hd__mux2_1 _419_ (.A0(_112_),
    .A1(_106_),
    .S(net87),
    .X(net63));
 sky130_fd_sc_hd__mux2_1 _420_ (.A0(_124_),
    .A1(_127_),
    .S(net87),
    .X(net64));
 sky130_fd_sc_hd__mux2_1 _421_ (.A0(_136_),
    .A1(_132_),
    .S(net87),
    .X(net65));
 sky130_fd_sc_hd__mux2_1 _422_ (.A0(_140_),
    .A1(_141_),
    .S(net87),
    .X(net66));
 sky130_fd_sc_hd__mux2_1 _423_ (.A0(_150_),
    .A1(_147_),
    .S(net88),
    .X(net67));
 sky130_fd_sc_hd__and2b_1 _424_ (.A_N(_153_),
    .B(_154_),
    .X(net68));
 sky130_fd_sc_hd__nand2_1 _425_ (.A(net111),
    .B(net1),
    .Y(_156_));
 sky130_fd_sc_hd__or2_1 _426_ (.A(net111),
    .B(net1),
    .X(_157_));
 sky130_fd_sc_hd__and2_1 _427_ (.A(_156_),
    .B(_157_),
    .X(_158_));
 sky130_fd_sc_hd__and2_1 _428_ (.A(net18),
    .B(net2),
    .X(_159_));
 sky130_fd_sc_hd__xor2_1 _429_ (.A(net18),
    .B(net2),
    .X(_160_));
 sky130_fd_sc_hd__a31o_1 _430_ (.A1(net111),
    .A2(net1),
    .A3(_160_),
    .B1(_159_),
    .X(_161_));
 sky130_fd_sc_hd__xnor2_1 _431_ (.A(_214_),
    .B(_161_),
    .Y(_162_));
 sky130_fd_sc_hd__nand2_1 _432_ (.A(net26),
    .B(net6),
    .Y(_163_));
 sky130_fd_sc_hd__nand2_2 _433_ (.A(net25),
    .B(net5),
    .Y(_164_));
 sky130_fd_sc_hd__xnor2_2 _434_ (.A(net26),
    .B(net6),
    .Y(_165_));
 sky130_fd_sc_hd__o21ai_4 _435_ (.A1(_164_),
    .A2(_165_),
    .B1(_163_),
    .Y(_166_));
 sky130_fd_sc_hd__xnor2_1 _436_ (.A(_215_),
    .B(_166_),
    .Y(_167_));
 sky130_fd_sc_hd__xnor2_1 _437_ (.A(net107),
    .B(_166_),
    .Y(_168_));
 sky130_fd_sc_hd__xor2_1 _438_ (.A(_164_),
    .B(_165_),
    .X(_169_));
 sky130_fd_sc_hd__xnor2_1 _439_ (.A(_164_),
    .B(_165_),
    .Y(_170_));
 sky130_fd_sc_hd__xnor2_1 _440_ (.A(_156_),
    .B(_160_),
    .Y(_171_));
 sky130_fd_sc_hd__or2_1 _441_ (.A(net25),
    .B(net5),
    .X(_172_));
 sky130_fd_sc_hd__and2_1 _442_ (.A(_164_),
    .B(_172_),
    .X(_173_));
 sky130_fd_sc_hd__nand2_1 _443_ (.A(_164_),
    .B(_172_),
    .Y(_174_));
 sky130_fd_sc_hd__a22o_1 _444_ (.A1(_170_),
    .A2(_171_),
    .B1(_174_),
    .B2(_158_),
    .X(_175_));
 sky130_fd_sc_hd__o221a_1 _445_ (.A1(_162_),
    .A2(_168_),
    .B1(_170_),
    .B2(_171_),
    .C1(_175_),
    .X(_176_));
 sky130_fd_sc_hd__or3b_1 _446_ (.A(_213_),
    .B(_214_),
    .C_N(_161_),
    .X(_177_));
 sky130_fd_sc_hd__a21o_1 _447_ (.A1(net110),
    .A2(_161_),
    .B1(net109),
    .X(_178_));
 sky130_fd_sc_hd__and2_1 _448_ (.A(_177_),
    .B(_178_),
    .X(_179_));
 sky130_fd_sc_hd__and3_1 _449_ (.A(net107),
    .B(net106),
    .C(_166_),
    .X(_180_));
 sky130_fd_sc_hd__a21oi_1 _450_ (.A1(net107),
    .A2(_166_),
    .B1(net106),
    .Y(_181_));
 sky130_fd_sc_hd__nor2_1 _451_ (.A(_180_),
    .B(_181_),
    .Y(_182_));
 sky130_fd_sc_hd__o211a_1 _452_ (.A1(_180_),
    .A2(_181_),
    .B1(_177_),
    .C1(_178_),
    .X(_183_));
 sky130_fd_sc_hd__and2_1 _453_ (.A(_162_),
    .B(_168_),
    .X(_184_));
 sky130_fd_sc_hd__a211o_1 _454_ (.A1(_177_),
    .A2(_178_),
    .B1(_180_),
    .C1(_181_),
    .X(_185_));
 sky130_fd_sc_hd__and4_1 _455_ (.A(net109),
    .B(net110),
    .C(net21),
    .D(_161_),
    .X(_186_));
 sky130_fd_sc_hd__or4b_2 _456_ (.A(_213_),
    .B(_214_),
    .C(_216_),
    .D_N(_161_),
    .X(_187_));
 sky130_fd_sc_hd__a31o_1 _457_ (.A1(net109),
    .A2(net110),
    .A3(_161_),
    .B1(net21),
    .X(_188_));
 sky130_fd_sc_hd__and2_1 _458_ (.A(_187_),
    .B(_188_),
    .X(_189_));
 sky130_fd_sc_hd__and4_2 _459_ (.A(net108),
    .B(net106),
    .C(net29),
    .D(_166_),
    .X(_190_));
 sky130_fd_sc_hd__a31oi_2 _460_ (.A1(net108),
    .A2(net106),
    .A3(_166_),
    .B1(net29),
    .Y(_191_));
 sky130_fd_sc_hd__nor2_1 _461_ (.A(_190_),
    .B(_191_),
    .Y(_192_));
 sky130_fd_sc_hd__a211o_1 _462_ (.A1(_187_),
    .A2(_188_),
    .B1(_190_),
    .C1(_191_),
    .X(_193_));
 sky130_fd_sc_hd__o311a_1 _463_ (.A1(_176_),
    .A2(_183_),
    .A3(_184_),
    .B1(_185_),
    .C1(_193_),
    .X(_194_));
 sky130_fd_sc_hd__xnor2_1 _464_ (.A(net105),
    .B(_190_),
    .Y(_195_));
 sky130_fd_sc_hd__inv_2 _465_ (.A(_195_),
    .Y(_196_));
 sky130_fd_sc_hd__xnor2_1 _466_ (.A(net22),
    .B(_187_),
    .Y(_197_));
 sky130_fd_sc_hd__o211a_1 _467_ (.A1(_190_),
    .A2(_191_),
    .B1(_187_),
    .C1(_188_),
    .X(_198_));
 sky130_fd_sc_hd__a21o_1 _468_ (.A1(_195_),
    .A2(_197_),
    .B1(_198_),
    .X(_199_));
 sky130_fd_sc_hd__or2_1 _469_ (.A(_195_),
    .B(_197_),
    .X(_200_));
 sky130_fd_sc_hd__and3_1 _470_ (.A(net23),
    .B(net22),
    .C(_186_),
    .X(_201_));
 sky130_fd_sc_hd__a21oi_1 _471_ (.A1(net22),
    .A2(_186_),
    .B1(net23),
    .Y(_202_));
 sky130_fd_sc_hd__nor2_1 _472_ (.A(_201_),
    .B(_202_),
    .Y(_203_));
 sky130_fd_sc_hd__and3_1 _473_ (.A(net31),
    .B(net105),
    .C(_190_),
    .X(_204_));
 sky130_fd_sc_hd__a21oi_1 _474_ (.A1(net105),
    .A2(_190_),
    .B1(net31),
    .Y(_205_));
 sky130_fd_sc_hd__or2_1 _475_ (.A(_204_),
    .B(_205_),
    .X(_206_));
 sky130_fd_sc_hd__inv_2 _476_ (.A(_206_),
    .Y(_207_));
 sky130_fd_sc_hd__o221a_1 _477_ (.A1(_194_),
    .A2(_199_),
    .B1(_203_),
    .B2(_206_),
    .C1(_200_),
    .X(_208_));
 sky130_fd_sc_hd__xnor2_1 _478_ (.A(net32),
    .B(_204_),
    .Y(_209_));
 sky130_fd_sc_hd__xor2_1 _479_ (.A(net24),
    .B(_201_),
    .X(_210_));
 sky130_fd_sc_hd__a22o_1 _480_ (.A1(_203_),
    .A2(_206_),
    .B1(_209_),
    .B2(_210_),
    .X(_211_));
 sky130_fd_sc_hd__o22a_1 _481_ (.A1(_209_),
    .A2(_210_),
    .B1(_211_),
    .B2(_208_),
    .X(net49));
 sky130_fd_sc_hd__mux2_1 _482_ (.A0(_158_),
    .A1(_173_),
    .S(net85),
    .X(net53));
 sky130_fd_sc_hd__mux2_1 _483_ (.A0(_171_),
    .A1(_169_),
    .S(net85),
    .X(net54));
 sky130_fd_sc_hd__mux2_1 _484_ (.A0(_162_),
    .A1(_167_),
    .S(net85),
    .X(net55));
 sky130_fd_sc_hd__mux2_1 _485_ (.A0(_179_),
    .A1(_182_),
    .S(net85),
    .X(net56));
 sky130_fd_sc_hd__mux2_1 _486_ (.A0(_189_),
    .A1(_192_),
    .S(net85),
    .X(net57));
 sky130_fd_sc_hd__mux2_1 _487_ (.A0(_197_),
    .A1(_196_),
    .S(net85),
    .X(net58));
 sky130_fd_sc_hd__mux2_1 _488_ (.A0(_203_),
    .A1(_207_),
    .S(net86),
    .X(net59));
 sky130_fd_sc_hd__and2b_1 _489_ (.A_N(_209_),
    .B(_210_),
    .X(net60));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_145 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(bm_s0_s0_i[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(bm_s0_s0_i[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(bm_s0_s2_i[0]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(bm_s0_s2_i[1]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(bm_s1_s0_i[0]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(bm_s1_s0_i[1]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(bm_s1_s2_i[0]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(bm_s1_s2_i[1]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(bm_s2_s1_i[0]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(bm_s2_s1_i[1]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(bm_s2_s3_i[0]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(bm_s2_s3_i[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(bm_s3_s1_i[0]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(bm_s3_s1_i[1]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(bm_s3_s3_i[0]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(bm_s3_s3_i[1]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(pm_s0_i[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(pm_s0_i[1]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(pm_s0_i[2]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(pm_s0_i[3]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(pm_s0_i[4]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(pm_s0_i[5]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(pm_s0_i[6]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(pm_s0_i[7]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(pm_s1_i[0]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(pm_s1_i[1]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(pm_s1_i[2]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(pm_s1_i[3]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(pm_s1_i[4]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(pm_s1_i[5]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(pm_s1_i[6]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(pm_s1_i[7]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(pm_s2_i[0]),
    .X(net33));
 sky130_fd_sc_hd__dlymetal6s2s_1 input34 (.A(pm_s2_i[1]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(pm_s2_i[2]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(pm_s2_i[3]),
    .X(net36));
 sky130_fd_sc_hd__dlymetal6s2s_1 input37 (.A(pm_s2_i[4]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(pm_s2_i[5]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(pm_s2_i[6]),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 input40 (.A(pm_s2_i[7]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(pm_s3_i[0]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input42 (.A(pm_s3_i[1]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(pm_s3_i[2]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(pm_s3_i[3]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(pm_s3_i[4]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(pm_s3_i[5]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(pm_s3_i[6]),
    .X(net47));
 sky130_fd_sc_hd__dlymetal6s2s_1 input48 (.A(pm_s3_i[7]),
    .X(net48));
 sky130_fd_sc_hd__buf_4 output49 (.A(net86),
    .X(dec_bits_o[0]));
 sky130_fd_sc_hd__buf_4 output50 (.A(net88),
    .X(dec_bits_o[1]));
 sky130_fd_sc_hd__buf_4 output51 (.A(net90),
    .X(dec_bits_o[2]));
 sky130_fd_sc_hd__buf_4 output52 (.A(net52),
    .X(dec_bits_o[3]));
 sky130_fd_sc_hd__buf_4 output53 (.A(net53),
    .X(pm_s0_o[0]));
 sky130_fd_sc_hd__buf_4 output54 (.A(net54),
    .X(pm_s0_o[1]));
 sky130_fd_sc_hd__buf_4 output55 (.A(net55),
    .X(pm_s0_o[2]));
 sky130_fd_sc_hd__buf_4 output56 (.A(net56),
    .X(pm_s0_o[3]));
 sky130_fd_sc_hd__buf_4 output57 (.A(net57),
    .X(pm_s0_o[4]));
 sky130_fd_sc_hd__buf_4 output58 (.A(net58),
    .X(pm_s0_o[5]));
 sky130_fd_sc_hd__buf_4 output59 (.A(net59),
    .X(pm_s0_o[6]));
 sky130_fd_sc_hd__buf_4 output60 (.A(net60),
    .X(pm_s0_o[7]));
 sky130_fd_sc_hd__buf_4 output61 (.A(net61),
    .X(pm_s1_o[0]));
 sky130_fd_sc_hd__buf_4 output62 (.A(net62),
    .X(pm_s1_o[1]));
 sky130_fd_sc_hd__buf_4 output63 (.A(net63),
    .X(pm_s1_o[2]));
 sky130_fd_sc_hd__buf_4 output64 (.A(net64),
    .X(pm_s1_o[3]));
 sky130_fd_sc_hd__buf_4 output65 (.A(net65),
    .X(pm_s1_o[4]));
 sky130_fd_sc_hd__buf_4 output66 (.A(net66),
    .X(pm_s1_o[5]));
 sky130_fd_sc_hd__buf_4 output67 (.A(net67),
    .X(pm_s1_o[6]));
 sky130_fd_sc_hd__buf_4 output68 (.A(net68),
    .X(pm_s1_o[7]));
 sky130_fd_sc_hd__buf_4 output69 (.A(net69),
    .X(pm_s2_o[0]));
 sky130_fd_sc_hd__buf_4 output70 (.A(net70),
    .X(pm_s2_o[1]));
 sky130_fd_sc_hd__buf_4 output71 (.A(net71),
    .X(pm_s2_o[2]));
 sky130_fd_sc_hd__buf_4 output72 (.A(net72),
    .X(pm_s2_o[3]));
 sky130_fd_sc_hd__buf_4 output73 (.A(net73),
    .X(pm_s2_o[4]));
 sky130_fd_sc_hd__buf_4 output74 (.A(net74),
    .X(pm_s2_o[5]));
 sky130_fd_sc_hd__buf_4 output75 (.A(net75),
    .X(pm_s2_o[6]));
 sky130_fd_sc_hd__buf_4 output76 (.A(net76),
    .X(pm_s2_o[7]));
 sky130_fd_sc_hd__buf_4 output77 (.A(net77),
    .X(pm_s3_o[0]));
 sky130_fd_sc_hd__buf_4 output78 (.A(net78),
    .X(pm_s3_o[1]));
 sky130_fd_sc_hd__buf_4 output79 (.A(net79),
    .X(pm_s3_o[2]));
 sky130_fd_sc_hd__buf_4 output80 (.A(net80),
    .X(pm_s3_o[3]));
 sky130_fd_sc_hd__buf_4 output81 (.A(net81),
    .X(pm_s3_o[4]));
 sky130_fd_sc_hd__buf_4 output82 (.A(net82),
    .X(pm_s3_o[5]));
 sky130_fd_sc_hd__buf_4 output83 (.A(net83),
    .X(pm_s3_o[6]));
 sky130_fd_sc_hd__buf_4 output84 (.A(net84),
    .X(pm_s3_o[7]));
 sky130_fd_sc_hd__clkbuf_2 fanout85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout86 (.A(net49),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 fanout87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout88 (.A(net50),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 fanout89 (.A(net90),
    .X(net89));
 sky130_fd_sc_hd__buf_1 fanout90 (.A(net51),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 fanout91 (.A(_045_),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 fanout92 (.A(_130_),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 fanout93 (.A(_080_),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 fanout94 (.A(_021_),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 fanout95 (.A(net46),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 fanout96 (.A(net44),
    .X(net96));
 sky130_fd_sc_hd__buf_1 fanout97 (.A(net44),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 fanout98 (.A(net43),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 fanout99 (.A(net43),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 fanout100 (.A(net38),
    .X(net100));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout101 (.A(net36),
    .X(net101));
 sky130_fd_sc_hd__buf_1 fanout102 (.A(net36),
    .X(net102));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout103 (.A(net35),
    .X(net103));
 sky130_fd_sc_hd__buf_1 fanout104 (.A(net35),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 fanout105 (.A(net30),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 fanout106 (.A(net28),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 fanout107 (.A(net27),
    .X(net107));
 sky130_fd_sc_hd__buf_1 fanout108 (.A(net27),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 fanout109 (.A(net20),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 fanout110 (.A(net19),
    .X(net110));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout111 (.A(net17),
    .X(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(bm_s0_s0_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(bm_s0_s0_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(bm_s0_s2_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(bm_s0_s2_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(bm_s1_s0_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(bm_s1_s0_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(bm_s1_s2_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(bm_s1_s2_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(bm_s2_s1_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(bm_s2_s1_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(bm_s2_s3_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(bm_s2_s3_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(bm_s3_s1_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(bm_s3_s1_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(bm_s3_s3_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(bm_s3_s3_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(pm_s0_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(pm_s0_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(pm_s0_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(pm_s0_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(pm_s0_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(pm_s0_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(pm_s0_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(pm_s0_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(pm_s1_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(pm_s1_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(pm_s1_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(pm_s1_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(pm_s1_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(pm_s1_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(pm_s1_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(pm_s1_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(pm_s2_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(pm_s2_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(pm_s2_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(pm_s2_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(pm_s2_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(pm_s2_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(pm_s2_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(pm_s2_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(pm_s3_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(pm_s3_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(pm_s3_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(pm_s3_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(pm_s3_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(pm_s3_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(pm_s3_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(pm_s3_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_X (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__304__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_X (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__488__S (.DIODE(net86));
 sky130_fd_sc_hd__decap_3 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_5 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_141 ();
endmodule
