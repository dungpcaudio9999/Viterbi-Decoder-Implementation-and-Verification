VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO system_top
  CLASS BLOCK ;
  FOREIGN system_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN busy_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END busy_o
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 374.990 1496.000 375.270 1500.000 ;
    END
  END clk
  PIN data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 149.640 1500.000 150.240 ;
    END
  END data_i[0]
  PIN data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 720.840 1500.000 721.440 ;
    END
  END data_i[10]
  PIN data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 777.960 1500.000 778.560 ;
    END
  END data_i[11]
  PIN data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 835.080 1500.000 835.680 ;
    END
  END data_i[12]
  PIN data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 892.200 1500.000 892.800 ;
    END
  END data_i[13]
  PIN data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 949.320 1500.000 949.920 ;
    END
  END data_i[14]
  PIN data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1006.440 1500.000 1007.040 ;
    END
  END data_i[15]
  PIN data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 206.760 1500.000 207.360 ;
    END
  END data_i[1]
  PIN data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 263.880 1500.000 264.480 ;
    END
  END data_i[2]
  PIN data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 321.000 1500.000 321.600 ;
    END
  END data_i[3]
  PIN data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 378.120 1500.000 378.720 ;
    END
  END data_i[4]
  PIN data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 435.240 1500.000 435.840 ;
    END
  END data_i[5]
  PIN data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 492.360 1500.000 492.960 ;
    END
  END data_i[6]
  PIN data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 549.480 1500.000 550.080 ;
    END
  END data_i[7]
  PIN data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 606.600 1500.000 607.200 ;
    END
  END data_i[8]
  PIN data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 663.720 1500.000 664.320 ;
    END
  END data_i[9]
  PIN data_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1063.560 1500.000 1064.160 ;
    END
  END data_o[0]
  PIN data_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1120.680 1500.000 1121.280 ;
    END
  END data_o[1]
  PIN data_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1177.800 1500.000 1178.400 ;
    END
  END data_o[2]
  PIN data_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1234.920 1500.000 1235.520 ;
    END
  END data_o[3]
  PIN data_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1292.040 1500.000 1292.640 ;
    END
  END data_o[4]
  PIN data_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1349.160 1500.000 1349.760 ;
    END
  END data_o[5]
  PIN data_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1406.280 1500.000 1406.880 ;
    END
  END data_o[6]
  PIN data_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1463.400 1500.000 1464.000 ;
    END
  END data_o[7]
  PIN dvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 35.400 1500.000 36.000 ;
    END
  END dvalid_i
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 1124.790 1496.000 1125.070 1500.000 ;
    END
  END rst_n
  PIN valid_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1496.000 92.520 1500.000 93.120 ;
    END
  END valid_o
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -47.480 -42.120 -44.480 1540.840 ;
    END
    PORT
      LAYER met5 ;
        RECT -47.480 -42.120 1547.080 -39.120 ;
    END
    PORT
      LAYER met5 ;
        RECT -47.480 1537.840 1547.080 1540.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1544.080 -42.120 1547.080 1540.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 -46.820 22.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 -46.820 72.640 74.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 925.800 72.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 -46.820 122.640 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 910.125 122.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 -46.820 172.640 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 910.125 172.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 -46.820 222.640 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 910.125 222.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 -46.820 272.640 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 910.125 272.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 -46.820 322.640 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 910.125 322.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 -46.820 372.640 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 910.125 372.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 -46.820 422.640 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 910.125 422.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 -46.820 472.640 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 910.125 472.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 -46.820 522.640 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 910.125 522.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 -46.820 572.640 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 910.125 572.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 -46.820 622.640 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 910.125 622.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.040 -46.820 672.640 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.040 910.125 672.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 721.040 -46.820 722.640 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 721.040 910.125 722.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 -46.820 772.640 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 910.125 772.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.040 -46.820 822.640 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.040 910.125 822.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 871.040 -46.820 872.640 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 871.040 910.125 872.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 -46.820 922.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 971.040 -46.820 972.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.040 -46.820 1022.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 -46.820 1072.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.040 -46.820 1122.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1171.040 -46.820 1172.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1221.040 -46.820 1222.640 50.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1221.040 240.360 1222.640 400.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1221.040 454.360 1222.640 750.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1221.040 820.680 1222.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1271.040 -46.820 1272.640 73.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1271.040 237.605 1272.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1321.040 -46.820 1322.640 73.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1321.040 237.605 1322.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.040 -46.820 1372.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1421.040 -46.820 1422.640 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1471.040 -46.820 1472.640 1545.540 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 26.730 1551.780 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 76.730 1551.780 78.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 126.730 42.080 128.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 176.730 88.660 178.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 226.730 88.660 228.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 276.730 42.080 278.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 326.730 88.660 328.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 376.730 88.660 378.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 426.730 42.080 428.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 476.730 88.660 478.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 526.730 88.660 528.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 576.730 42.080 578.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 626.730 88.660 628.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 676.730 88.660 678.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 726.730 42.080 728.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 776.730 88.660 778.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 826.730 88.660 828.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 876.730 42.080 878.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 926.730 1551.780 928.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 976.730 1551.780 978.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1026.730 42.080 1028.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1076.730 1551.780 1078.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1126.730 1551.780 1128.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1176.730 1551.780 1178.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1226.730 1551.780 1228.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1276.730 1551.780 1278.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1326.730 1551.780 1328.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1376.730 1551.780 1378.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1426.730 1551.780 1428.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1476.730 1551.780 1478.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 176.730 1551.780 178.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 226.730 1551.780 228.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 326.730 1551.780 328.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 376.730 1551.780 378.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 476.730 1551.780 478.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 526.730 1551.780 528.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 626.730 1551.780 628.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 676.730 1551.780 678.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 776.730 1551.780 778.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 826.730 1551.780 828.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 1057.500 126.730 1551.780 128.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 1057.500 276.730 1551.780 278.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 1057.500 426.730 1551.780 428.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 1057.500 576.730 1551.780 578.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 1057.500 726.730 1551.780 728.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 1057.500 876.730 1551.780 878.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 1057.500 1026.730 1551.780 1028.330 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -52.180 -46.820 -49.180 1545.540 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 -46.820 1551.780 -43.820 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1542.540 1551.780 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1548.780 -46.820 1551.780 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.340 -46.820 25.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.340 -46.820 75.940 74.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.340 925.800 75.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 124.340 -46.820 125.940 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 124.340 910.125 125.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.340 -46.820 175.940 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.340 910.125 175.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 224.340 -46.820 225.940 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 224.340 910.125 225.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 274.340 -46.820 275.940 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 274.340 910.125 275.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 324.340 -46.820 325.940 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 324.340 910.125 325.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 374.340 -46.820 375.940 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 374.340 910.125 375.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.340 -46.820 425.940 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.340 910.125 425.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 474.340 -46.820 475.940 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 474.340 910.125 475.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 524.340 -46.820 525.940 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 524.340 910.125 525.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 574.340 -46.820 575.940 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 574.340 910.125 575.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 624.340 -46.820 625.940 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 624.340 910.125 625.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 674.340 -46.820 675.940 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 674.340 910.125 675.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.340 -46.820 725.940 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.340 910.125 725.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 774.340 -46.820 775.940 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 774.340 910.125 775.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 824.340 -46.820 825.940 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 824.340 910.125 825.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.340 -46.820 875.940 45.995 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.340 910.125 875.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 924.340 -46.820 925.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 974.340 -46.820 975.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1024.340 -46.820 1025.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1074.340 -46.820 1075.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1124.340 -46.820 1125.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1174.340 -46.820 1175.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1224.340 -46.820 1225.940 50.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1224.340 240.360 1225.940 400.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1224.340 454.360 1225.940 750.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1224.340 820.680 1225.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1274.340 -46.820 1275.940 73.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1274.340 237.605 1275.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.340 -46.820 1325.940 73.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.340 237.605 1325.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1374.340 -46.820 1375.940 50.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1374.340 240.360 1375.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1424.340 -46.820 1425.940 1545.540 ;
    END
    PORT
      LAYER met4 ;
        RECT 1474.340 -46.820 1475.940 1545.540 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 30.030 1551.780 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 80.030 1551.780 81.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 130.030 1551.780 131.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 180.030 88.660 181.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 230.030 88.660 231.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 280.030 88.660 281.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 330.030 88.660 331.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 380.030 88.660 381.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 430.030 88.660 431.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 480.030 88.660 481.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 530.030 88.660 531.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 580.030 88.660 581.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 630.030 88.660 631.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 680.030 88.660 681.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 730.030 88.660 731.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 780.030 88.660 781.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 830.030 88.660 831.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 880.030 88.660 881.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 930.030 1551.780 931.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 980.030 1551.780 981.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1030.030 1551.780 1031.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1080.030 1551.780 1081.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1130.030 1551.780 1131.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1180.030 1551.780 1181.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1230.030 1551.780 1231.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1280.030 1551.780 1281.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1330.030 1551.780 1331.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1380.030 1551.780 1381.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1430.030 1551.780 1431.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -52.180 1480.030 1551.780 1481.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 180.030 1551.780 181.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 230.030 1551.780 231.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 280.030 1551.780 281.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 330.030 1551.780 331.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 380.030 1551.780 381.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 430.030 1551.780 431.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 480.030 1551.780 481.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 530.030 1551.780 531.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 580.030 1551.780 581.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 630.030 1551.780 631.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 680.030 1551.780 681.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 730.030 1551.780 731.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 780.030 1551.780 781.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 830.030 1551.780 831.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 909.260 880.030 1551.780 881.630 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 1494.270 1488.030 ;
      LAYER li1 ;
        RECT 5.520 10.795 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 5.520 10.640 1494.080 1496.640 ;
      LAYER met2 ;
        RECT 21.070 1495.720 374.710 1496.670 ;
        RECT 375.550 1495.720 1124.510 1496.670 ;
        RECT 1125.350 1495.720 1492.150 1496.670 ;
        RECT 21.070 4.280 1492.150 1495.720 ;
        RECT 21.070 4.000 749.610 4.280 ;
        RECT 750.450 4.000 1492.150 4.280 ;
      LAYER met3 ;
        RECT 21.050 1464.400 1496.000 1488.005 ;
        RECT 21.050 1463.000 1495.600 1464.400 ;
        RECT 21.050 1407.280 1496.000 1463.000 ;
        RECT 21.050 1405.880 1495.600 1407.280 ;
        RECT 21.050 1350.160 1496.000 1405.880 ;
        RECT 21.050 1348.760 1495.600 1350.160 ;
        RECT 21.050 1293.040 1496.000 1348.760 ;
        RECT 21.050 1291.640 1495.600 1293.040 ;
        RECT 21.050 1235.920 1496.000 1291.640 ;
        RECT 21.050 1234.520 1495.600 1235.920 ;
        RECT 21.050 1178.800 1496.000 1234.520 ;
        RECT 21.050 1177.400 1495.600 1178.800 ;
        RECT 21.050 1121.680 1496.000 1177.400 ;
        RECT 21.050 1120.280 1495.600 1121.680 ;
        RECT 21.050 1064.560 1496.000 1120.280 ;
        RECT 21.050 1063.160 1495.600 1064.560 ;
        RECT 21.050 1007.440 1496.000 1063.160 ;
        RECT 21.050 1006.040 1495.600 1007.440 ;
        RECT 21.050 950.320 1496.000 1006.040 ;
        RECT 21.050 948.920 1495.600 950.320 ;
        RECT 21.050 893.200 1496.000 948.920 ;
        RECT 21.050 891.800 1495.600 893.200 ;
        RECT 21.050 836.080 1496.000 891.800 ;
        RECT 21.050 834.680 1495.600 836.080 ;
        RECT 21.050 778.960 1496.000 834.680 ;
        RECT 21.050 777.560 1495.600 778.960 ;
        RECT 21.050 721.840 1496.000 777.560 ;
        RECT 21.050 720.440 1495.600 721.840 ;
        RECT 21.050 664.720 1496.000 720.440 ;
        RECT 21.050 663.320 1495.600 664.720 ;
        RECT 21.050 607.600 1496.000 663.320 ;
        RECT 21.050 606.200 1495.600 607.600 ;
        RECT 21.050 550.480 1496.000 606.200 ;
        RECT 21.050 549.080 1495.600 550.480 ;
        RECT 21.050 493.360 1496.000 549.080 ;
        RECT 21.050 491.960 1495.600 493.360 ;
        RECT 21.050 436.240 1496.000 491.960 ;
        RECT 21.050 434.840 1495.600 436.240 ;
        RECT 21.050 379.120 1496.000 434.840 ;
        RECT 21.050 377.720 1495.600 379.120 ;
        RECT 21.050 322.000 1496.000 377.720 ;
        RECT 21.050 320.600 1495.600 322.000 ;
        RECT 21.050 264.880 1496.000 320.600 ;
        RECT 21.050 263.480 1495.600 264.880 ;
        RECT 21.050 207.760 1496.000 263.480 ;
        RECT 21.050 206.360 1495.600 207.760 ;
        RECT 21.050 150.640 1496.000 206.360 ;
        RECT 21.050 149.240 1495.600 150.640 ;
        RECT 21.050 93.520 1496.000 149.240 ;
        RECT 21.050 92.120 1495.600 93.520 ;
        RECT 21.050 36.400 1496.000 92.120 ;
        RECT 21.050 35.000 1495.600 36.400 ;
        RECT 21.050 10.715 1496.000 35.000 ;
      LAYER met4 ;
        RECT 69.900 925.400 70.640 1037.600 ;
        RECT 73.040 925.400 73.940 1037.600 ;
        RECT 76.340 925.400 120.640 1037.600 ;
        RECT 69.900 909.725 120.640 925.400 ;
        RECT 123.040 909.725 123.940 1037.600 ;
        RECT 126.340 909.725 170.640 1037.600 ;
        RECT 173.040 909.725 173.940 1037.600 ;
        RECT 176.340 909.725 220.640 1037.600 ;
        RECT 223.040 909.725 223.940 1037.600 ;
        RECT 226.340 909.725 270.640 1037.600 ;
        RECT 273.040 909.725 273.940 1037.600 ;
        RECT 276.340 909.725 320.640 1037.600 ;
        RECT 323.040 909.725 323.940 1037.600 ;
        RECT 326.340 909.725 370.640 1037.600 ;
        RECT 373.040 909.725 373.940 1037.600 ;
        RECT 376.340 909.725 420.640 1037.600 ;
        RECT 423.040 909.725 423.940 1037.600 ;
        RECT 426.340 909.725 470.640 1037.600 ;
        RECT 473.040 909.725 473.940 1037.600 ;
        RECT 476.340 909.725 520.640 1037.600 ;
        RECT 523.040 909.725 523.940 1037.600 ;
        RECT 526.340 909.725 570.640 1037.600 ;
        RECT 573.040 909.725 573.940 1037.600 ;
        RECT 576.340 909.725 620.640 1037.600 ;
        RECT 623.040 909.725 623.940 1037.600 ;
        RECT 626.340 909.725 670.640 1037.600 ;
        RECT 673.040 909.725 673.940 1037.600 ;
        RECT 676.340 909.725 720.640 1037.600 ;
        RECT 723.040 909.725 723.940 1037.600 ;
        RECT 726.340 909.725 770.640 1037.600 ;
        RECT 773.040 909.725 773.940 1037.600 ;
        RECT 776.340 909.725 820.640 1037.600 ;
        RECT 823.040 909.725 823.940 1037.600 ;
        RECT 826.340 909.725 870.640 1037.600 ;
        RECT 873.040 909.725 873.940 1037.600 ;
        RECT 876.340 909.725 920.640 1037.600 ;
        RECT 69.900 74.920 920.640 909.725 ;
        RECT 69.900 54.575 70.640 74.920 ;
        RECT 73.040 54.575 73.940 74.920 ;
        RECT 76.340 54.575 920.640 74.920 ;
        RECT 923.040 54.575 923.940 1037.600 ;
        RECT 926.340 54.575 970.640 1037.600 ;
        RECT 973.040 54.575 973.940 1037.600 ;
        RECT 976.340 54.575 1020.640 1037.600 ;
        RECT 1023.040 54.575 1023.940 1037.600 ;
        RECT 1026.340 54.575 1070.640 1037.600 ;
        RECT 1073.040 54.575 1073.940 1037.600 ;
        RECT 1076.340 54.575 1120.640 1037.600 ;
        RECT 1123.040 54.575 1123.940 1037.600 ;
        RECT 1126.340 54.575 1170.640 1037.600 ;
        RECT 1173.040 54.575 1173.940 1037.600 ;
        RECT 1176.340 820.280 1220.640 1037.600 ;
        RECT 1223.040 820.280 1223.940 1037.600 ;
        RECT 1226.340 820.280 1270.640 1037.600 ;
        RECT 1176.340 750.440 1270.640 820.280 ;
        RECT 1176.340 453.960 1220.640 750.440 ;
        RECT 1223.040 453.960 1223.940 750.440 ;
        RECT 1226.340 453.960 1270.640 750.440 ;
        RECT 1176.340 400.440 1270.640 453.960 ;
        RECT 1176.340 239.960 1220.640 400.440 ;
        RECT 1223.040 239.960 1223.940 400.440 ;
        RECT 1226.340 239.960 1270.640 400.440 ;
        RECT 1176.340 237.205 1270.640 239.960 ;
        RECT 1273.040 237.205 1273.940 1037.600 ;
        RECT 1276.340 237.205 1320.640 1037.600 ;
        RECT 1323.040 237.205 1323.940 1037.600 ;
        RECT 1326.340 237.205 1370.640 1037.600 ;
        RECT 1176.340 74.275 1370.640 237.205 ;
        RECT 1176.340 54.575 1270.640 74.275 ;
        RECT 1273.040 54.575 1273.940 74.275 ;
        RECT 1276.340 54.575 1320.640 74.275 ;
        RECT 1323.040 54.575 1323.940 74.275 ;
        RECT 1326.340 54.575 1370.640 74.275 ;
        RECT 1373.040 239.960 1373.940 1037.600 ;
        RECT 1376.340 239.960 1382.465 1037.600 ;
        RECT 1373.040 54.575 1382.465 239.960 ;
      LAYER met5 ;
        RECT 55.280 983.230 1212.900 1024.980 ;
        RECT 55.280 933.230 1212.900 975.130 ;
        RECT 55.280 883.230 1212.900 925.130 ;
        RECT 90.260 878.430 907.660 883.230 ;
        RECT 55.280 875.130 1055.900 878.430 ;
        RECT 55.280 833.230 1212.900 875.130 ;
        RECT 90.260 825.130 907.660 833.230 ;
        RECT 55.280 783.230 1212.900 825.130 ;
        RECT 90.260 775.130 907.660 783.230 ;
        RECT 55.280 733.230 1212.900 775.130 ;
        RECT 90.260 728.430 907.660 733.230 ;
        RECT 55.280 725.130 1055.900 728.430 ;
        RECT 55.280 683.230 1212.900 725.130 ;
        RECT 90.260 675.130 907.660 683.230 ;
        RECT 55.280 633.230 1212.900 675.130 ;
        RECT 90.260 625.130 907.660 633.230 ;
        RECT 55.280 583.230 1212.900 625.130 ;
        RECT 90.260 578.430 907.660 583.230 ;
        RECT 55.280 575.130 1055.900 578.430 ;
        RECT 55.280 533.230 1212.900 575.130 ;
        RECT 90.260 525.130 907.660 533.230 ;
        RECT 55.280 483.230 1212.900 525.130 ;
        RECT 90.260 475.130 907.660 483.230 ;
        RECT 55.280 433.230 1212.900 475.130 ;
        RECT 90.260 428.430 907.660 433.230 ;
        RECT 55.280 425.130 1055.900 428.430 ;
        RECT 55.280 383.230 1212.900 425.130 ;
        RECT 90.260 375.130 907.660 383.230 ;
        RECT 55.280 333.230 1212.900 375.130 ;
        RECT 90.260 325.130 907.660 333.230 ;
        RECT 55.280 283.230 1212.900 325.130 ;
        RECT 90.260 278.430 907.660 283.230 ;
        RECT 55.280 275.130 1055.900 278.430 ;
        RECT 55.280 233.230 1212.900 275.130 ;
        RECT 90.260 225.130 907.660 233.230 ;
        RECT 55.280 183.230 1212.900 225.130 ;
        RECT 90.260 175.130 907.660 183.230 ;
        RECT 55.280 133.230 1212.900 175.130 ;
        RECT 55.280 125.130 1055.900 128.430 ;
        RECT 55.280 113.100 1212.900 125.130 ;
  END
END system_top
END LIBRARY

