VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sipo
  CLASS BLOCK ;
  FOREIGN sipo ;
  ORIGIN 0.000 0.000 ;
  SIZE 45.245 BY 55.965 ;
  PIN byte_ready_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 41.245 49.000 45.245 49.600 ;
    END
  END byte_ready_o
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END clk
  PIN data_parallel_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 41.245 5.480 45.245 6.080 ;
    END
  END data_parallel_o[0]
  PIN data_parallel_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 41.245 10.920 45.245 11.520 ;
    END
  END data_parallel_o[1]
  PIN data_parallel_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 41.245 16.360 45.245 16.960 ;
    END
  END data_parallel_o[2]
  PIN data_parallel_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 41.245 21.800 45.245 22.400 ;
    END
  END data_parallel_o[3]
  PIN data_parallel_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 41.245 27.240 45.245 27.840 ;
    END
  END data_parallel_o[4]
  PIN data_parallel_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 41.245 32.680 45.245 33.280 ;
    END
  END data_parallel_o[5]
  PIN data_parallel_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 41.245 38.120 45.245 38.720 ;
    END
  END data_parallel_o[6]
  PIN data_parallel_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 41.245 43.560 45.245 44.160 ;
    END
  END data_parallel_o[7]
  PIN data_serial_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END data_serial_i
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END rst_n
  PIN valid_serial_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END valid_serial_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.840 10.640 22.840 43.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.540 10.640 26.540 43.760 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 39.750 43.605 ;
      LAYER li1 ;
        RECT 5.520 10.795 39.560 43.605 ;
      LAYER met1 ;
        RECT 5.520 10.240 39.560 43.760 ;
      LAYER met2 ;
        RECT 6.530 5.595 38.090 49.485 ;
      LAYER met3 ;
        RECT 4.000 48.640 40.845 49.465 ;
        RECT 4.400 48.600 40.845 48.640 ;
        RECT 4.400 47.240 41.245 48.600 ;
        RECT 4.000 44.560 41.245 47.240 ;
        RECT 4.000 43.160 40.845 44.560 ;
        RECT 4.000 39.120 41.245 43.160 ;
        RECT 4.000 37.720 40.845 39.120 ;
        RECT 4.000 35.040 41.245 37.720 ;
        RECT 4.400 33.680 41.245 35.040 ;
        RECT 4.400 33.640 40.845 33.680 ;
        RECT 4.000 32.280 40.845 33.640 ;
        RECT 4.000 28.240 41.245 32.280 ;
        RECT 4.000 26.840 40.845 28.240 ;
        RECT 4.000 22.800 41.245 26.840 ;
        RECT 4.000 21.440 40.845 22.800 ;
        RECT 4.400 21.400 40.845 21.440 ;
        RECT 4.400 20.040 41.245 21.400 ;
        RECT 4.000 17.360 41.245 20.040 ;
        RECT 4.000 15.960 40.845 17.360 ;
        RECT 4.000 11.920 41.245 15.960 ;
        RECT 4.000 10.520 40.845 11.920 ;
        RECT 4.000 7.840 41.245 10.520 ;
        RECT 4.400 6.480 41.245 7.840 ;
        RECT 4.400 6.440 40.845 6.480 ;
        RECT 4.000 5.615 40.845 6.440 ;
  END
END sipo
END LIBRARY

