magic
tech sky130A
magscale 1 2
timestamp 1769196443
<< viali >>
rect 6837 8517 6871 8551
rect 7389 8517 7423 8551
rect 1409 8449 1443 8483
rect 1685 8449 1719 8483
rect 6561 8449 6595 8483
rect 7113 8449 7147 8483
rect 1593 8313 1627 8347
rect 2605 7905 2639 7939
rect 6745 7905 6779 7939
rect 2881 7837 2915 7871
rect 7113 7837 7147 7871
rect 2421 7769 2455 7803
rect 3065 7769 3099 7803
rect 6469 7769 6503 7803
rect 7389 7769 7423 7803
rect 1961 7701 1995 7735
rect 2329 7701 2363 7735
rect 6101 7701 6135 7735
rect 6561 7701 6595 7735
rect 6837 7497 6871 7531
rect 1777 7429 1811 7463
rect 6745 7361 6779 7395
rect 7389 7361 7423 7395
rect 1501 7293 1535 7327
rect 3249 7293 3283 7327
rect 4261 7293 4295 7327
rect 4537 7293 4571 7327
rect 6009 7293 6043 7327
rect 7021 7293 7055 7327
rect 7205 7225 7239 7259
rect 6377 7157 6411 7191
rect 1593 6953 1627 6987
rect 4169 6953 4203 6987
rect 5536 6953 5570 6987
rect 7021 6953 7055 6987
rect 1869 6817 1903 6851
rect 1409 6749 1443 6783
rect 1685 6749 1719 6783
rect 3801 6749 3835 6783
rect 3985 6749 4019 6783
rect 5273 6749 5307 6783
rect 7113 6749 7147 6783
rect 2145 6681 2179 6715
rect 7389 6681 7423 6715
rect 3617 6613 3651 6647
rect 6193 6409 6227 6443
rect 6745 6409 6779 6443
rect 6837 6409 6871 6443
rect 4261 6341 4295 6375
rect 1593 6273 1627 6307
rect 1777 6273 1811 6307
rect 2237 6273 2271 6307
rect 2697 6273 2731 6307
rect 4445 6273 4479 6307
rect 1869 6205 1903 6239
rect 2329 6205 2363 6239
rect 4721 6205 4755 6239
rect 6929 6205 6963 6239
rect 6377 6137 6411 6171
rect 1777 6069 1811 6103
rect 2126 5865 2160 5899
rect 3617 5865 3651 5899
rect 3985 5865 4019 5899
rect 4261 5865 4295 5899
rect 7113 5865 7147 5899
rect 3801 5797 3835 5831
rect 1869 5729 1903 5763
rect 5365 5729 5399 5763
rect 4261 5661 4295 5695
rect 4537 5661 4571 5695
rect 3969 5593 4003 5627
rect 4169 5593 4203 5627
rect 4445 5593 4479 5627
rect 4813 5593 4847 5627
rect 5641 5593 5675 5627
rect 4721 5525 4755 5559
rect 3709 5321 3743 5355
rect 5181 5321 5215 5355
rect 6653 5321 6687 5355
rect 5917 5253 5951 5287
rect 1685 5185 1719 5219
rect 3617 5185 3651 5219
rect 3893 5185 3927 5219
rect 6193 5185 6227 5219
rect 6745 5185 6779 5219
rect 1961 5117 1995 5151
rect 6561 5117 6595 5151
rect 3433 4981 3467 5015
rect 7113 4981 7147 5015
rect 1777 4777 1811 4811
rect 7113 4777 7147 4811
rect 1593 4709 1627 4743
rect 2237 4641 2271 4675
rect 1409 4573 1443 4607
rect 2145 4573 2179 4607
rect 5825 4573 5859 4607
rect 3801 4437 3835 4471
rect 6837 4233 6871 4267
rect 1409 4165 1443 4199
rect 6193 4097 6227 4131
rect 6745 4097 6779 4131
rect 5917 4029 5951 4063
rect 6929 4029 6963 4063
rect 4445 3893 4479 3927
rect 6377 3893 6411 3927
rect 5365 3689 5399 3723
rect 5089 3553 5123 3587
rect 6837 3553 6871 3587
rect 7113 3553 7147 3587
rect 5273 3485 5307 3519
rect 6377 3145 6411 3179
rect 6837 3145 6871 3179
rect 5917 3077 5951 3111
rect 6745 3077 6779 3111
rect 4353 3009 4387 3043
rect 6193 3009 6227 3043
rect 4169 2941 4203 2975
rect 6929 2941 6963 2975
rect 4445 2805 4479 2839
rect 4445 2533 4479 2567
rect 6377 2533 6411 2567
rect 4077 2465 4111 2499
rect 5917 2465 5951 2499
rect 6193 2465 6227 2499
rect 6929 2465 6963 2499
rect 3617 2397 3651 2431
rect 4353 2397 4387 2431
rect 6745 2397 6779 2431
rect 3341 2329 3375 2363
rect 6837 2261 6871 2295
<< metal1 >>
rect 1104 8730 7912 8752
rect 1104 8678 4922 8730
rect 4974 8678 4986 8730
rect 5038 8678 5050 8730
rect 5102 8678 5114 8730
rect 5166 8678 5178 8730
rect 5230 8678 5242 8730
rect 5294 8678 7912 8730
rect 1104 8656 7912 8678
rect 6822 8508 6828 8560
rect 6880 8508 6886 8560
rect 7374 8508 7380 8560
rect 7432 8508 7438 8560
rect 1302 8440 1308 8492
rect 1360 8480 1366 8492
rect 1397 8483 1455 8489
rect 1397 8480 1409 8483
rect 1360 8452 1409 8480
rect 1360 8440 1366 8452
rect 1397 8449 1409 8452
rect 1443 8480 1455 8483
rect 1673 8483 1731 8489
rect 1673 8480 1685 8483
rect 1443 8452 1685 8480
rect 1443 8449 1455 8452
rect 1397 8443 1455 8449
rect 1673 8449 1685 8452
rect 1719 8449 1731 8483
rect 1673 8443 1731 8449
rect 6546 8440 6552 8492
rect 6604 8440 6610 8492
rect 6638 8440 6644 8492
rect 6696 8480 6702 8492
rect 7101 8483 7159 8489
rect 7101 8480 7113 8483
rect 6696 8452 7113 8480
rect 6696 8440 6702 8452
rect 7101 8449 7113 8452
rect 7147 8449 7159 8483
rect 7101 8443 7159 8449
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 2866 8344 2872 8356
rect 1627 8316 2872 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 2866 8304 2872 8316
rect 2924 8304 2930 8356
rect 1104 8186 7912 8208
rect 1104 8134 4182 8186
rect 4234 8134 4246 8186
rect 4298 8134 4310 8186
rect 4362 8134 4374 8186
rect 4426 8134 4438 8186
rect 4490 8134 4502 8186
rect 4554 8134 7912 8186
rect 1104 8112 7912 8134
rect 2593 7939 2651 7945
rect 2593 7905 2605 7939
rect 2639 7905 2651 7939
rect 2593 7899 2651 7905
rect 1578 7760 1584 7812
rect 1636 7800 1642 7812
rect 2409 7803 2467 7809
rect 2409 7800 2421 7803
rect 1636 7772 2421 7800
rect 1636 7760 1642 7772
rect 2409 7769 2421 7772
rect 2455 7769 2467 7803
rect 2608 7800 2636 7899
rect 6730 7896 6736 7948
rect 6788 7896 6794 7948
rect 2866 7828 2872 7880
rect 2924 7828 2930 7880
rect 7101 7871 7159 7877
rect 7101 7868 7113 7871
rect 6932 7840 7113 7868
rect 2958 7800 2964 7812
rect 2608 7772 2964 7800
rect 2409 7763 2467 7769
rect 2958 7760 2964 7772
rect 3016 7800 3022 7812
rect 3053 7803 3111 7809
rect 3053 7800 3065 7803
rect 3016 7772 3065 7800
rect 3016 7760 3022 7772
rect 3053 7769 3065 7772
rect 3099 7800 3111 7803
rect 5810 7800 5816 7812
rect 3099 7772 5816 7800
rect 3099 7769 3111 7772
rect 3053 7763 3111 7769
rect 5810 7760 5816 7772
rect 5868 7760 5874 7812
rect 6457 7803 6515 7809
rect 6457 7769 6469 7803
rect 6503 7800 6515 7803
rect 6822 7800 6828 7812
rect 6503 7772 6828 7800
rect 6503 7769 6515 7772
rect 6457 7763 6515 7769
rect 6822 7760 6828 7772
rect 6880 7760 6886 7812
rect 6932 7744 6960 7840
rect 7101 7837 7113 7840
rect 7147 7837 7159 7871
rect 7101 7831 7159 7837
rect 7374 7760 7380 7812
rect 7432 7760 7438 7812
rect 1762 7692 1768 7744
rect 1820 7732 1826 7744
rect 1949 7735 2007 7741
rect 1949 7732 1961 7735
rect 1820 7704 1961 7732
rect 1820 7692 1826 7704
rect 1949 7701 1961 7704
rect 1995 7701 2007 7735
rect 1949 7695 2007 7701
rect 2317 7735 2375 7741
rect 2317 7701 2329 7735
rect 2363 7732 2375 7735
rect 2498 7732 2504 7744
rect 2363 7704 2504 7732
rect 2363 7701 2375 7704
rect 2317 7695 2375 7701
rect 2498 7692 2504 7704
rect 2556 7692 2562 7744
rect 5718 7692 5724 7744
rect 5776 7732 5782 7744
rect 6089 7735 6147 7741
rect 6089 7732 6101 7735
rect 5776 7704 6101 7732
rect 5776 7692 5782 7704
rect 6089 7701 6101 7704
rect 6135 7701 6147 7735
rect 6089 7695 6147 7701
rect 6549 7735 6607 7741
rect 6549 7701 6561 7735
rect 6595 7732 6607 7735
rect 6914 7732 6920 7744
rect 6595 7704 6920 7732
rect 6595 7701 6607 7704
rect 6549 7695 6607 7701
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 1104 7642 7912 7664
rect 1104 7590 4922 7642
rect 4974 7590 4986 7642
rect 5038 7590 5050 7642
rect 5102 7590 5114 7642
rect 5166 7590 5178 7642
rect 5230 7590 5242 7642
rect 5294 7590 7912 7642
rect 1104 7568 7912 7590
rect 2498 7488 2504 7540
rect 2556 7528 2562 7540
rect 6638 7528 6644 7540
rect 2556 7500 6644 7528
rect 2556 7488 2562 7500
rect 1762 7420 1768 7472
rect 1820 7420 1826 7472
rect 3234 7460 3240 7472
rect 2990 7432 3240 7460
rect 3234 7420 3240 7432
rect 3292 7420 3298 7472
rect 1486 7284 1492 7336
rect 1544 7284 1550 7336
rect 3237 7327 3295 7333
rect 3237 7293 3249 7327
rect 3283 7324 3295 7327
rect 3344 7324 3372 7500
rect 6638 7488 6644 7500
rect 6696 7528 6702 7540
rect 6825 7531 6883 7537
rect 6825 7528 6837 7531
rect 6696 7500 6837 7528
rect 6696 7488 6702 7500
rect 6825 7497 6837 7500
rect 6871 7497 6883 7531
rect 6825 7491 6883 7497
rect 5994 7460 6000 7472
rect 5750 7432 6000 7460
rect 5994 7420 6000 7432
rect 6052 7420 6058 7472
rect 5810 7352 5816 7404
rect 5868 7392 5874 7404
rect 6733 7395 6791 7401
rect 5868 7364 6684 7392
rect 5868 7352 5874 7364
rect 3283 7296 3372 7324
rect 4249 7327 4307 7333
rect 3283 7293 3295 7296
rect 3237 7287 3295 7293
rect 4249 7293 4261 7327
rect 4295 7293 4307 7327
rect 4249 7287 4307 7293
rect 4525 7327 4583 7333
rect 4525 7293 4537 7327
rect 4571 7324 4583 7327
rect 4614 7324 4620 7336
rect 4571 7296 4620 7324
rect 4571 7293 4583 7296
rect 4525 7287 4583 7293
rect 4264 7188 4292 7287
rect 4614 7284 4620 7296
rect 4672 7284 4678 7336
rect 5997 7327 6055 7333
rect 5997 7293 6009 7327
rect 6043 7324 6055 7327
rect 6546 7324 6552 7336
rect 6043 7296 6552 7324
rect 6043 7293 6055 7296
rect 5997 7287 6055 7293
rect 6546 7284 6552 7296
rect 6604 7284 6610 7336
rect 6656 7324 6684 7364
rect 6733 7361 6745 7395
rect 6779 7392 6791 7395
rect 6914 7392 6920 7404
rect 6779 7364 6920 7392
rect 6779 7361 6791 7364
rect 6733 7355 6791 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 7024 7364 7389 7392
rect 7024 7333 7052 7364
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 7009 7327 7067 7333
rect 7009 7324 7021 7327
rect 6656 7296 7021 7324
rect 7009 7293 7021 7296
rect 7055 7293 7067 7327
rect 7009 7287 7067 7293
rect 6730 7216 6736 7268
rect 6788 7256 6794 7268
rect 7193 7259 7251 7265
rect 7193 7256 7205 7259
rect 6788 7228 7205 7256
rect 6788 7216 6794 7228
rect 7193 7225 7205 7228
rect 7239 7225 7251 7259
rect 7193 7219 7251 7225
rect 4614 7188 4620 7200
rect 4264 7160 4620 7188
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 6086 7148 6092 7200
rect 6144 7188 6150 7200
rect 6365 7191 6423 7197
rect 6365 7188 6377 7191
rect 6144 7160 6377 7188
rect 6144 7148 6150 7160
rect 6365 7157 6377 7160
rect 6411 7157 6423 7191
rect 6365 7151 6423 7157
rect 1104 7098 7912 7120
rect 1104 7046 4182 7098
rect 4234 7046 4246 7098
rect 4298 7046 4310 7098
rect 4362 7046 4374 7098
rect 4426 7046 4438 7098
rect 4490 7046 4502 7098
rect 4554 7046 7912 7098
rect 1104 7024 7912 7046
rect 1578 6944 1584 6996
rect 1636 6944 1642 6996
rect 4157 6987 4215 6993
rect 4157 6953 4169 6987
rect 4203 6984 4215 6987
rect 4706 6984 4712 6996
rect 4203 6956 4712 6984
rect 4203 6953 4215 6956
rect 4157 6947 4215 6953
rect 4706 6944 4712 6956
rect 4764 6944 4770 6996
rect 5524 6987 5582 6993
rect 5524 6953 5536 6987
rect 5570 6984 5582 6987
rect 6086 6984 6092 6996
rect 5570 6956 6092 6984
rect 5570 6953 5582 6956
rect 5524 6947 5582 6953
rect 6086 6944 6092 6956
rect 6144 6944 6150 6996
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 7009 6987 7067 6993
rect 7009 6984 7021 6987
rect 6972 6956 7021 6984
rect 6972 6944 6978 6956
rect 7009 6953 7021 6956
rect 7055 6953 7067 6987
rect 7009 6947 7067 6953
rect 1486 6808 1492 6860
rect 1544 6848 1550 6860
rect 1857 6851 1915 6857
rect 1857 6848 1869 6851
rect 1544 6820 1869 6848
rect 1544 6808 1550 6820
rect 1857 6817 1869 6820
rect 1903 6848 1915 6851
rect 2682 6848 2688 6860
rect 1903 6820 2688 6848
rect 1903 6817 1915 6820
rect 1857 6811 1915 6817
rect 2682 6808 2688 6820
rect 2740 6808 2746 6860
rect 3602 6808 3608 6860
rect 3660 6848 3666 6860
rect 3660 6820 6684 6848
rect 3660 6808 3666 6820
rect 1302 6740 1308 6792
rect 1360 6780 1366 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 1360 6752 1409 6780
rect 1360 6740 1366 6752
rect 1397 6749 1409 6752
rect 1443 6780 1455 6783
rect 1673 6783 1731 6789
rect 1673 6780 1685 6783
rect 1443 6752 1685 6780
rect 1443 6749 1455 6752
rect 1397 6743 1455 6749
rect 1673 6749 1685 6752
rect 1719 6749 1731 6783
rect 1673 6743 1731 6749
rect 3234 6740 3240 6792
rect 3292 6740 3298 6792
rect 3789 6783 3847 6789
rect 3789 6749 3801 6783
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 1854 6672 1860 6724
rect 1912 6712 1918 6724
rect 2133 6715 2191 6721
rect 2133 6712 2145 6715
rect 1912 6684 2145 6712
rect 1912 6672 1918 6684
rect 2133 6681 2145 6684
rect 2179 6681 2191 6715
rect 2133 6675 2191 6681
rect 2222 6604 2228 6656
rect 2280 6644 2286 6656
rect 3605 6647 3663 6653
rect 3605 6644 3617 6647
rect 2280 6616 3617 6644
rect 2280 6604 2286 6616
rect 3605 6613 3617 6616
rect 3651 6644 3663 6647
rect 3804 6644 3832 6743
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3936 6752 3985 6780
rect 3936 6740 3942 6752
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6749 5319 6783
rect 6656 6766 6684 6820
rect 5261 6743 5319 6749
rect 5276 6712 5304 6743
rect 6822 6740 6828 6792
rect 6880 6780 6886 6792
rect 7101 6783 7159 6789
rect 7101 6780 7113 6783
rect 6880 6752 7113 6780
rect 6880 6740 6886 6752
rect 7101 6749 7113 6752
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 5276 6684 5396 6712
rect 5368 6656 5396 6684
rect 7374 6672 7380 6724
rect 7432 6672 7438 6724
rect 3651 6616 3832 6644
rect 3651 6613 3663 6616
rect 3605 6607 3663 6613
rect 5350 6604 5356 6656
rect 5408 6604 5414 6656
rect 1104 6554 7912 6576
rect 1104 6502 4922 6554
rect 4974 6502 4986 6554
rect 5038 6502 5050 6554
rect 5102 6502 5114 6554
rect 5166 6502 5178 6554
rect 5230 6502 5242 6554
rect 5294 6502 7912 6554
rect 1104 6480 7912 6502
rect 6181 6443 6239 6449
rect 6181 6409 6193 6443
rect 6227 6440 6239 6443
rect 6638 6440 6644 6452
rect 6227 6412 6644 6440
rect 6227 6409 6239 6412
rect 6181 6403 6239 6409
rect 6638 6400 6644 6412
rect 6696 6440 6702 6452
rect 6733 6443 6791 6449
rect 6733 6440 6745 6443
rect 6696 6412 6745 6440
rect 6696 6400 6702 6412
rect 6733 6409 6745 6412
rect 6779 6409 6791 6443
rect 6733 6403 6791 6409
rect 6822 6400 6828 6452
rect 6880 6400 6886 6452
rect 4249 6375 4307 6381
rect 1596 6344 2360 6372
rect 1596 6313 1624 6344
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6273 1639 6307
rect 1581 6267 1639 6273
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 1780 6168 1808 6267
rect 2222 6264 2228 6316
rect 2280 6264 2286 6316
rect 1854 6196 1860 6248
rect 1912 6196 1918 6248
rect 2332 6245 2360 6344
rect 4249 6341 4261 6375
rect 4295 6372 4307 6375
rect 4798 6372 4804 6384
rect 4295 6344 4804 6372
rect 4295 6341 4307 6344
rect 4249 6335 4307 6341
rect 4798 6332 4804 6344
rect 4856 6332 4862 6384
rect 6086 6372 6092 6384
rect 5934 6344 6092 6372
rect 6086 6332 6092 6344
rect 6144 6332 6150 6384
rect 2682 6264 2688 6316
rect 2740 6304 2746 6316
rect 4430 6304 4436 6316
rect 2740 6276 4436 6304
rect 2740 6264 2746 6276
rect 4430 6264 4436 6276
rect 4488 6264 4494 6316
rect 2317 6239 2375 6245
rect 2317 6205 2329 6239
rect 2363 6236 2375 6239
rect 3878 6236 3884 6248
rect 2363 6208 3884 6236
rect 2363 6205 2375 6208
rect 2317 6199 2375 6205
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6236 4767 6239
rect 4755 6208 6408 6236
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 4062 6168 4068 6180
rect 1780 6140 4068 6168
rect 4062 6128 4068 6140
rect 4120 6128 4126 6180
rect 6380 6177 6408 6208
rect 6546 6196 6552 6248
rect 6604 6236 6610 6248
rect 6730 6236 6736 6248
rect 6604 6208 6736 6236
rect 6604 6196 6610 6208
rect 6730 6196 6736 6208
rect 6788 6236 6794 6248
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 6788 6208 6929 6236
rect 6788 6196 6794 6208
rect 6917 6205 6929 6208
rect 6963 6205 6975 6239
rect 6917 6199 6975 6205
rect 6365 6171 6423 6177
rect 6365 6137 6377 6171
rect 6411 6137 6423 6171
rect 6365 6131 6423 6137
rect 1762 6060 1768 6112
rect 1820 6060 1826 6112
rect 3234 6060 3240 6112
rect 3292 6100 3298 6112
rect 6086 6100 6092 6112
rect 3292 6072 6092 6100
rect 3292 6060 3298 6072
rect 6086 6060 6092 6072
rect 6144 6060 6150 6112
rect 1104 6010 7912 6032
rect 1104 5958 4182 6010
rect 4234 5958 4246 6010
rect 4298 5958 4310 6010
rect 4362 5958 4374 6010
rect 4426 5958 4438 6010
rect 4490 5958 4502 6010
rect 4554 5958 7912 6010
rect 1104 5936 7912 5958
rect 1762 5856 1768 5908
rect 1820 5896 1826 5908
rect 2114 5899 2172 5905
rect 2114 5896 2126 5899
rect 1820 5868 2126 5896
rect 1820 5856 1826 5868
rect 2114 5865 2126 5868
rect 2160 5865 2172 5899
rect 2114 5859 2172 5865
rect 3605 5899 3663 5905
rect 3605 5865 3617 5899
rect 3651 5896 3663 5899
rect 3973 5899 4031 5905
rect 3973 5896 3985 5899
rect 3651 5868 3985 5896
rect 3651 5865 3663 5868
rect 3605 5859 3663 5865
rect 3973 5865 3985 5868
rect 4019 5865 4031 5899
rect 3973 5859 4031 5865
rect 3789 5831 3847 5837
rect 3789 5797 3801 5831
rect 3835 5828 3847 5831
rect 3878 5828 3884 5840
rect 3835 5800 3884 5828
rect 3835 5797 3847 5800
rect 3789 5791 3847 5797
rect 3878 5788 3884 5800
rect 3936 5788 3942 5840
rect 1670 5720 1676 5772
rect 1728 5760 1734 5772
rect 1857 5763 1915 5769
rect 1857 5760 1869 5763
rect 1728 5732 1869 5760
rect 1728 5720 1734 5732
rect 1857 5729 1869 5732
rect 1903 5760 1915 5763
rect 2682 5760 2688 5772
rect 1903 5732 2688 5760
rect 1903 5729 1915 5732
rect 1857 5723 1915 5729
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 3234 5652 3240 5704
rect 3292 5652 3298 5704
rect 3988 5692 4016 5859
rect 4062 5856 4068 5908
rect 4120 5896 4126 5908
rect 4249 5899 4307 5905
rect 4249 5896 4261 5899
rect 4120 5868 4261 5896
rect 4120 5856 4126 5868
rect 4249 5865 4261 5868
rect 4295 5865 4307 5899
rect 4249 5859 4307 5865
rect 6822 5856 6828 5908
rect 6880 5896 6886 5908
rect 7101 5899 7159 5905
rect 7101 5896 7113 5899
rect 6880 5868 7113 5896
rect 6880 5856 6886 5868
rect 7101 5865 7113 5868
rect 7147 5865 7159 5899
rect 7101 5859 7159 5865
rect 4062 5720 4068 5772
rect 4120 5760 4126 5772
rect 4120 5732 4568 5760
rect 4120 5720 4126 5732
rect 4540 5701 4568 5732
rect 5350 5720 5356 5772
rect 5408 5760 5414 5772
rect 7098 5760 7104 5772
rect 5408 5732 7104 5760
rect 5408 5720 5414 5732
rect 7098 5720 7104 5732
rect 7156 5720 7162 5772
rect 4249 5695 4307 5701
rect 4249 5692 4261 5695
rect 3988 5664 4261 5692
rect 4249 5661 4261 5664
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 3970 5633 3976 5636
rect 3957 5627 3976 5633
rect 3957 5593 3969 5627
rect 3957 5587 3976 5593
rect 3970 5584 3976 5587
rect 4028 5584 4034 5636
rect 4154 5584 4160 5636
rect 4212 5624 4218 5636
rect 4433 5627 4491 5633
rect 4433 5624 4445 5627
rect 4212 5596 4445 5624
rect 4212 5584 4218 5596
rect 4433 5593 4445 5596
rect 4479 5593 4491 5627
rect 4433 5587 4491 5593
rect 4614 5584 4620 5636
rect 4672 5624 4678 5636
rect 4801 5627 4859 5633
rect 4801 5624 4813 5627
rect 4672 5596 4813 5624
rect 4672 5584 4678 5596
rect 4801 5593 4813 5596
rect 4847 5593 4859 5627
rect 4801 5587 4859 5593
rect 5629 5627 5687 5633
rect 5629 5593 5641 5627
rect 5675 5624 5687 5627
rect 5718 5624 5724 5636
rect 5675 5596 5724 5624
rect 5675 5593 5687 5596
rect 5629 5587 5687 5593
rect 5718 5584 5724 5596
rect 5776 5584 5782 5636
rect 6086 5624 6092 5636
rect 5828 5596 6092 5624
rect 4709 5559 4767 5565
rect 4709 5525 4721 5559
rect 4755 5556 4767 5559
rect 5828 5556 5856 5596
rect 6086 5584 6092 5596
rect 6144 5584 6150 5636
rect 4755 5528 5856 5556
rect 4755 5525 4767 5528
rect 4709 5519 4767 5525
rect 1104 5466 7912 5488
rect 1104 5414 4922 5466
rect 4974 5414 4986 5466
rect 5038 5414 5050 5466
rect 5102 5414 5114 5466
rect 5166 5414 5178 5466
rect 5230 5414 5242 5466
rect 5294 5414 7912 5466
rect 1104 5392 7912 5414
rect 3697 5355 3755 5361
rect 3697 5321 3709 5355
rect 3743 5352 3755 5355
rect 4614 5352 4620 5364
rect 3743 5324 4620 5352
rect 3743 5321 3755 5324
rect 3697 5315 3755 5321
rect 3712 5284 3740 5315
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 4798 5312 4804 5364
rect 4856 5352 4862 5364
rect 5169 5355 5227 5361
rect 5169 5352 5181 5355
rect 4856 5324 5181 5352
rect 4856 5312 4862 5324
rect 5169 5321 5181 5324
rect 5215 5321 5227 5355
rect 5169 5315 5227 5321
rect 6638 5312 6644 5364
rect 6696 5312 6702 5364
rect 3174 5256 3740 5284
rect 5902 5244 5908 5296
rect 5960 5244 5966 5296
rect 1670 5176 1676 5228
rect 1728 5176 1734 5228
rect 3602 5176 3608 5228
rect 3660 5176 3666 5228
rect 3786 5176 3792 5228
rect 3844 5216 3850 5228
rect 3881 5219 3939 5225
rect 3881 5216 3893 5219
rect 3844 5188 3893 5216
rect 3844 5176 3850 5188
rect 3881 5185 3893 5188
rect 3927 5185 3939 5219
rect 3881 5179 3939 5185
rect 6181 5219 6239 5225
rect 6181 5185 6193 5219
rect 6227 5216 6239 5219
rect 6656 5216 6684 5312
rect 6227 5188 6684 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 6730 5176 6736 5228
rect 6788 5176 6794 5228
rect 1946 5108 1952 5160
rect 2004 5108 2010 5160
rect 6546 5108 6552 5160
rect 6604 5108 6610 5160
rect 3418 4972 3424 5024
rect 3476 5012 3482 5024
rect 4154 5012 4160 5024
rect 3476 4984 4160 5012
rect 3476 4972 3482 4984
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 6822 4972 6828 5024
rect 6880 5012 6886 5024
rect 7101 5015 7159 5021
rect 7101 5012 7113 5015
rect 6880 4984 7113 5012
rect 6880 4972 6886 4984
rect 7101 4981 7113 4984
rect 7147 4981 7159 5015
rect 7101 4975 7159 4981
rect 1104 4922 7912 4944
rect 1104 4870 4182 4922
rect 4234 4870 4246 4922
rect 4298 4870 4310 4922
rect 4362 4870 4374 4922
rect 4426 4870 4438 4922
rect 4490 4870 4502 4922
rect 4554 4870 7912 4922
rect 1104 4848 7912 4870
rect 1765 4811 1823 4817
rect 1765 4777 1777 4811
rect 1811 4808 1823 4811
rect 1946 4808 1952 4820
rect 1811 4780 1952 4808
rect 1811 4777 1823 4780
rect 1765 4771 1823 4777
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 7098 4768 7104 4820
rect 7156 4768 7162 4820
rect 1581 4743 1639 4749
rect 1581 4709 1593 4743
rect 1627 4740 1639 4743
rect 3602 4740 3608 4752
rect 1627 4712 3608 4740
rect 1627 4709 1639 4712
rect 1581 4703 1639 4709
rect 3602 4700 3608 4712
rect 3660 4700 3666 4752
rect 2225 4675 2283 4681
rect 2225 4641 2237 4675
rect 2271 4672 2283 4675
rect 2958 4672 2964 4684
rect 2271 4644 2964 4672
rect 2271 4641 2283 4644
rect 2225 4635 2283 4641
rect 2958 4632 2964 4644
rect 3016 4672 3022 4684
rect 3970 4672 3976 4684
rect 3016 4644 3976 4672
rect 3016 4632 3022 4644
rect 3970 4632 3976 4644
rect 4028 4632 4034 4684
rect 1394 4564 1400 4616
rect 1452 4564 1458 4616
rect 2133 4607 2191 4613
rect 2133 4573 2145 4607
rect 2179 4604 2191 4607
rect 3418 4604 3424 4616
rect 2179 4576 3424 4604
rect 2179 4573 2191 4576
rect 2133 4567 2191 4573
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 4798 4564 4804 4616
rect 4856 4604 4862 4616
rect 5813 4607 5871 4613
rect 5813 4604 5825 4607
rect 4856 4576 5825 4604
rect 4856 4564 4862 4576
rect 5813 4573 5825 4576
rect 5859 4573 5871 4607
rect 5813 4567 5871 4573
rect 3786 4428 3792 4480
rect 3844 4428 3850 4480
rect 1104 4378 7912 4400
rect 1104 4326 4922 4378
rect 4974 4326 4986 4378
rect 5038 4326 5050 4378
rect 5102 4326 5114 4378
rect 5166 4326 5178 4378
rect 5230 4326 5242 4378
rect 5294 4326 7912 4378
rect 1104 4304 7912 4326
rect 6730 4224 6736 4276
rect 6788 4264 6794 4276
rect 6825 4267 6883 4273
rect 6825 4264 6837 4267
rect 6788 4236 6837 4264
rect 6788 4224 6794 4236
rect 6825 4233 6837 4236
rect 6871 4233 6883 4267
rect 6825 4227 6883 4233
rect 1394 4156 1400 4208
rect 1452 4156 1458 4208
rect 4614 4156 4620 4208
rect 4672 4196 4678 4208
rect 4672 4168 4738 4196
rect 4672 4156 4678 4168
rect 6178 4088 6184 4140
rect 6236 4128 6242 4140
rect 6236 4100 6408 4128
rect 6236 4088 6242 4100
rect 5810 4020 5816 4072
rect 5868 4060 5874 4072
rect 5905 4063 5963 4069
rect 5905 4060 5917 4063
rect 5868 4032 5917 4060
rect 5868 4020 5874 4032
rect 5905 4029 5917 4032
rect 5951 4029 5963 4063
rect 5905 4023 5963 4029
rect 6380 3992 6408 4100
rect 6638 4088 6644 4140
rect 6696 4128 6702 4140
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 6696 4100 6745 4128
rect 6696 4088 6702 4100
rect 6733 4097 6745 4100
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 6546 4020 6552 4072
rect 6604 4060 6610 4072
rect 6917 4063 6975 4069
rect 6917 4060 6929 4063
rect 6604 4032 6929 4060
rect 6604 4020 6610 4032
rect 6917 4029 6929 4032
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 7098 3992 7104 4004
rect 6380 3964 7104 3992
rect 7098 3952 7104 3964
rect 7156 3952 7162 4004
rect 4433 3927 4491 3933
rect 4433 3893 4445 3927
rect 4479 3924 4491 3927
rect 4614 3924 4620 3936
rect 4479 3896 4620 3924
rect 4479 3893 4491 3896
rect 4433 3887 4491 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 5902 3884 5908 3936
rect 5960 3924 5966 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 5960 3896 6377 3924
rect 5960 3884 5966 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 1104 3834 7912 3856
rect 1104 3782 4182 3834
rect 4234 3782 4246 3834
rect 4298 3782 4310 3834
rect 4362 3782 4374 3834
rect 4426 3782 4438 3834
rect 4490 3782 4502 3834
rect 4554 3782 7912 3834
rect 1104 3760 7912 3782
rect 5353 3723 5411 3729
rect 5353 3689 5365 3723
rect 5399 3720 5411 3723
rect 6730 3720 6736 3732
rect 5399 3692 6736 3720
rect 5399 3689 5411 3692
rect 5353 3683 5411 3689
rect 5077 3587 5135 3593
rect 5077 3553 5089 3587
rect 5123 3584 5135 3587
rect 5442 3584 5448 3596
rect 5123 3556 5448 3584
rect 5123 3553 5135 3556
rect 5077 3547 5135 3553
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3516 5319 3519
rect 5539 3516 5567 3692
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 6822 3544 6828 3596
rect 6880 3544 6886 3596
rect 7098 3544 7104 3596
rect 7156 3544 7162 3596
rect 5307 3488 5567 3516
rect 5307 3485 5319 3488
rect 5261 3479 5319 3485
rect 4798 3408 4804 3460
rect 4856 3448 4862 3460
rect 4856 3420 5658 3448
rect 4856 3408 4862 3420
rect 4614 3340 4620 3392
rect 4672 3380 4678 3392
rect 6730 3380 6736 3392
rect 4672 3352 6736 3380
rect 4672 3340 4678 3352
rect 6730 3340 6736 3352
rect 6788 3340 6794 3392
rect 1104 3290 7912 3312
rect 1104 3238 4922 3290
rect 4974 3238 4986 3290
rect 5038 3238 5050 3290
rect 5102 3238 5114 3290
rect 5166 3238 5178 3290
rect 5230 3238 5242 3290
rect 5294 3238 7912 3290
rect 1104 3216 7912 3238
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 6365 3179 6423 3185
rect 6365 3176 6377 3179
rect 5868 3148 6377 3176
rect 5868 3136 5874 3148
rect 6365 3145 6377 3148
rect 6411 3145 6423 3179
rect 6365 3139 6423 3145
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 6825 3179 6883 3185
rect 6825 3176 6837 3179
rect 6696 3148 6837 3176
rect 6696 3136 6702 3148
rect 6825 3145 6837 3148
rect 6871 3145 6883 3179
rect 6825 3139 6883 3145
rect 5902 3068 5908 3120
rect 5960 3068 5966 3120
rect 6730 3068 6736 3120
rect 6788 3068 6794 3120
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3040 4399 3043
rect 4614 3040 4620 3052
rect 4387 3012 4620 3040
rect 4387 3009 4399 3012
rect 4341 3003 4399 3009
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 4798 3000 4804 3052
rect 4856 3000 4862 3052
rect 6178 3000 6184 3052
rect 6236 3000 6242 3052
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2972 4215 2975
rect 4203 2944 6132 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 6104 2904 6132 2944
rect 6546 2932 6552 2984
rect 6604 2972 6610 2984
rect 6917 2975 6975 2981
rect 6917 2972 6929 2975
rect 6604 2944 6929 2972
rect 6604 2932 6610 2944
rect 6917 2941 6929 2944
rect 6963 2941 6975 2975
rect 6917 2935 6975 2941
rect 7558 2904 7564 2916
rect 6104 2876 7564 2904
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 4433 2839 4491 2845
rect 4433 2805 4445 2839
rect 4479 2836 4491 2839
rect 4614 2836 4620 2848
rect 4479 2808 4620 2836
rect 4479 2805 4491 2808
rect 4433 2799 4491 2805
rect 4614 2796 4620 2808
rect 4672 2836 4678 2848
rect 6638 2836 6644 2848
rect 4672 2808 6644 2836
rect 4672 2796 4678 2808
rect 6638 2796 6644 2808
rect 6696 2796 6702 2848
rect 1104 2746 7912 2768
rect 1104 2694 4182 2746
rect 4234 2694 4246 2746
rect 4298 2694 4310 2746
rect 4362 2694 4374 2746
rect 4426 2694 4438 2746
rect 4490 2694 4502 2746
rect 4554 2694 7912 2746
rect 1104 2672 7912 2694
rect 7190 2632 7196 2644
rect 4908 2604 7196 2632
rect 4430 2524 4436 2576
rect 4488 2524 4494 2576
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 4908 2496 4936 2604
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 6365 2567 6423 2573
rect 6365 2564 6377 2567
rect 6104 2536 6377 2564
rect 4111 2468 4936 2496
rect 5905 2499 5963 2505
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 5905 2465 5917 2499
rect 5951 2496 5963 2499
rect 6104 2496 6132 2536
rect 6365 2533 6377 2536
rect 6411 2533 6423 2567
rect 6365 2527 6423 2533
rect 5951 2468 6132 2496
rect 5951 2465 5963 2468
rect 5905 2459 5963 2465
rect 6178 2456 6184 2508
rect 6236 2456 6242 2508
rect 6546 2456 6552 2508
rect 6604 2496 6610 2508
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6604 2468 6929 2496
rect 6604 2456 6610 2468
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2397 3663 2431
rect 3605 2391 3663 2397
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 4614 2428 4620 2440
rect 4387 2400 4620 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 3329 2363 3387 2369
rect 3329 2329 3341 2363
rect 3375 2329 3387 2363
rect 3620 2360 3648 2391
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 4798 2388 4804 2440
rect 4856 2388 4862 2440
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 6512 2400 6745 2428
rect 6512 2388 6518 2400
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 4430 2360 4436 2372
rect 3620 2332 4436 2360
rect 3329 2323 3387 2329
rect 3344 2292 3372 2323
rect 4430 2320 4436 2332
rect 4488 2320 4494 2372
rect 7374 2360 7380 2372
rect 6012 2332 7380 2360
rect 6012 2292 6040 2332
rect 7374 2320 7380 2332
rect 7432 2320 7438 2372
rect 3344 2264 6040 2292
rect 6730 2252 6736 2304
rect 6788 2292 6794 2304
rect 6825 2295 6883 2301
rect 6825 2292 6837 2295
rect 6788 2264 6837 2292
rect 6788 2252 6794 2264
rect 6825 2261 6837 2264
rect 6871 2261 6883 2295
rect 6825 2255 6883 2261
rect 1104 2202 7912 2224
rect 1104 2150 4922 2202
rect 4974 2150 4986 2202
rect 5038 2150 5050 2202
rect 5102 2150 5114 2202
rect 5166 2150 5178 2202
rect 5230 2150 5242 2202
rect 5294 2150 7912 2202
rect 1104 2128 7912 2150
rect 4430 2048 4436 2100
rect 4488 2088 4494 2100
rect 6454 2088 6460 2100
rect 4488 2060 6460 2088
rect 4488 2048 4494 2060
rect 6454 2048 6460 2060
rect 6512 2048 6518 2100
<< via1 >>
rect 4922 8678 4974 8730
rect 4986 8678 5038 8730
rect 5050 8678 5102 8730
rect 5114 8678 5166 8730
rect 5178 8678 5230 8730
rect 5242 8678 5294 8730
rect 6828 8551 6880 8560
rect 6828 8517 6837 8551
rect 6837 8517 6871 8551
rect 6871 8517 6880 8551
rect 6828 8508 6880 8517
rect 7380 8551 7432 8560
rect 7380 8517 7389 8551
rect 7389 8517 7423 8551
rect 7423 8517 7432 8551
rect 7380 8508 7432 8517
rect 1308 8440 1360 8492
rect 6552 8483 6604 8492
rect 6552 8449 6561 8483
rect 6561 8449 6595 8483
rect 6595 8449 6604 8483
rect 6552 8440 6604 8449
rect 6644 8440 6696 8492
rect 2872 8304 2924 8356
rect 4182 8134 4234 8186
rect 4246 8134 4298 8186
rect 4310 8134 4362 8186
rect 4374 8134 4426 8186
rect 4438 8134 4490 8186
rect 4502 8134 4554 8186
rect 1584 7760 1636 7812
rect 6736 7939 6788 7948
rect 6736 7905 6745 7939
rect 6745 7905 6779 7939
rect 6779 7905 6788 7939
rect 6736 7896 6788 7905
rect 2872 7871 2924 7880
rect 2872 7837 2881 7871
rect 2881 7837 2915 7871
rect 2915 7837 2924 7871
rect 2872 7828 2924 7837
rect 2964 7760 3016 7812
rect 5816 7760 5868 7812
rect 6828 7760 6880 7812
rect 7380 7803 7432 7812
rect 7380 7769 7389 7803
rect 7389 7769 7423 7803
rect 7423 7769 7432 7803
rect 7380 7760 7432 7769
rect 1768 7692 1820 7744
rect 2504 7692 2556 7744
rect 5724 7692 5776 7744
rect 6920 7692 6972 7744
rect 4922 7590 4974 7642
rect 4986 7590 5038 7642
rect 5050 7590 5102 7642
rect 5114 7590 5166 7642
rect 5178 7590 5230 7642
rect 5242 7590 5294 7642
rect 2504 7488 2556 7540
rect 1768 7463 1820 7472
rect 1768 7429 1777 7463
rect 1777 7429 1811 7463
rect 1811 7429 1820 7463
rect 1768 7420 1820 7429
rect 3240 7420 3292 7472
rect 1492 7327 1544 7336
rect 1492 7293 1501 7327
rect 1501 7293 1535 7327
rect 1535 7293 1544 7327
rect 1492 7284 1544 7293
rect 6644 7488 6696 7540
rect 6000 7420 6052 7472
rect 5816 7352 5868 7404
rect 4620 7284 4672 7336
rect 6552 7284 6604 7336
rect 6920 7352 6972 7404
rect 6736 7216 6788 7268
rect 4620 7148 4672 7200
rect 6092 7148 6144 7200
rect 4182 7046 4234 7098
rect 4246 7046 4298 7098
rect 4310 7046 4362 7098
rect 4374 7046 4426 7098
rect 4438 7046 4490 7098
rect 4502 7046 4554 7098
rect 1584 6987 1636 6996
rect 1584 6953 1593 6987
rect 1593 6953 1627 6987
rect 1627 6953 1636 6987
rect 1584 6944 1636 6953
rect 4712 6944 4764 6996
rect 6092 6944 6144 6996
rect 6920 6944 6972 6996
rect 1492 6808 1544 6860
rect 2688 6808 2740 6860
rect 3608 6808 3660 6860
rect 1308 6740 1360 6792
rect 3240 6740 3292 6792
rect 1860 6672 1912 6724
rect 2228 6604 2280 6656
rect 3884 6740 3936 6792
rect 6828 6740 6880 6792
rect 7380 6715 7432 6724
rect 7380 6681 7389 6715
rect 7389 6681 7423 6715
rect 7423 6681 7432 6715
rect 7380 6672 7432 6681
rect 5356 6604 5408 6656
rect 4922 6502 4974 6554
rect 4986 6502 5038 6554
rect 5050 6502 5102 6554
rect 5114 6502 5166 6554
rect 5178 6502 5230 6554
rect 5242 6502 5294 6554
rect 6644 6400 6696 6452
rect 6828 6443 6880 6452
rect 6828 6409 6837 6443
rect 6837 6409 6871 6443
rect 6871 6409 6880 6443
rect 6828 6400 6880 6409
rect 2228 6307 2280 6316
rect 2228 6273 2237 6307
rect 2237 6273 2271 6307
rect 2271 6273 2280 6307
rect 2228 6264 2280 6273
rect 1860 6239 1912 6248
rect 1860 6205 1869 6239
rect 1869 6205 1903 6239
rect 1903 6205 1912 6239
rect 1860 6196 1912 6205
rect 4804 6332 4856 6384
rect 6092 6332 6144 6384
rect 2688 6307 2740 6316
rect 2688 6273 2697 6307
rect 2697 6273 2731 6307
rect 2731 6273 2740 6307
rect 4436 6307 4488 6316
rect 2688 6264 2740 6273
rect 4436 6273 4445 6307
rect 4445 6273 4479 6307
rect 4479 6273 4488 6307
rect 4436 6264 4488 6273
rect 3884 6196 3936 6248
rect 4068 6128 4120 6180
rect 6552 6196 6604 6248
rect 6736 6196 6788 6248
rect 1768 6103 1820 6112
rect 1768 6069 1777 6103
rect 1777 6069 1811 6103
rect 1811 6069 1820 6103
rect 1768 6060 1820 6069
rect 3240 6060 3292 6112
rect 6092 6060 6144 6112
rect 4182 5958 4234 6010
rect 4246 5958 4298 6010
rect 4310 5958 4362 6010
rect 4374 5958 4426 6010
rect 4438 5958 4490 6010
rect 4502 5958 4554 6010
rect 1768 5856 1820 5908
rect 3884 5788 3936 5840
rect 1676 5720 1728 5772
rect 2688 5720 2740 5772
rect 3240 5652 3292 5704
rect 4068 5856 4120 5908
rect 6828 5856 6880 5908
rect 4068 5720 4120 5772
rect 5356 5763 5408 5772
rect 5356 5729 5365 5763
rect 5365 5729 5399 5763
rect 5399 5729 5408 5763
rect 5356 5720 5408 5729
rect 7104 5720 7156 5772
rect 3976 5627 4028 5636
rect 3976 5593 4003 5627
rect 4003 5593 4028 5627
rect 3976 5584 4028 5593
rect 4160 5627 4212 5636
rect 4160 5593 4169 5627
rect 4169 5593 4203 5627
rect 4203 5593 4212 5627
rect 4160 5584 4212 5593
rect 4620 5584 4672 5636
rect 5724 5584 5776 5636
rect 6092 5584 6144 5636
rect 4922 5414 4974 5466
rect 4986 5414 5038 5466
rect 5050 5414 5102 5466
rect 5114 5414 5166 5466
rect 5178 5414 5230 5466
rect 5242 5414 5294 5466
rect 4620 5312 4672 5364
rect 4804 5312 4856 5364
rect 6644 5355 6696 5364
rect 6644 5321 6653 5355
rect 6653 5321 6687 5355
rect 6687 5321 6696 5355
rect 6644 5312 6696 5321
rect 5908 5287 5960 5296
rect 5908 5253 5917 5287
rect 5917 5253 5951 5287
rect 5951 5253 5960 5287
rect 5908 5244 5960 5253
rect 1676 5219 1728 5228
rect 1676 5185 1685 5219
rect 1685 5185 1719 5219
rect 1719 5185 1728 5219
rect 1676 5176 1728 5185
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 3792 5176 3844 5228
rect 6736 5219 6788 5228
rect 6736 5185 6745 5219
rect 6745 5185 6779 5219
rect 6779 5185 6788 5219
rect 6736 5176 6788 5185
rect 1952 5151 2004 5160
rect 1952 5117 1961 5151
rect 1961 5117 1995 5151
rect 1995 5117 2004 5151
rect 1952 5108 2004 5117
rect 6552 5151 6604 5160
rect 6552 5117 6561 5151
rect 6561 5117 6595 5151
rect 6595 5117 6604 5151
rect 6552 5108 6604 5117
rect 3424 5015 3476 5024
rect 3424 4981 3433 5015
rect 3433 4981 3467 5015
rect 3467 4981 3476 5015
rect 3424 4972 3476 4981
rect 4160 4972 4212 5024
rect 6828 4972 6880 5024
rect 4182 4870 4234 4922
rect 4246 4870 4298 4922
rect 4310 4870 4362 4922
rect 4374 4870 4426 4922
rect 4438 4870 4490 4922
rect 4502 4870 4554 4922
rect 1952 4768 2004 4820
rect 7104 4811 7156 4820
rect 7104 4777 7113 4811
rect 7113 4777 7147 4811
rect 7147 4777 7156 4811
rect 7104 4768 7156 4777
rect 3608 4700 3660 4752
rect 2964 4632 3016 4684
rect 3976 4632 4028 4684
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 3424 4564 3476 4616
rect 4804 4564 4856 4616
rect 3792 4471 3844 4480
rect 3792 4437 3801 4471
rect 3801 4437 3835 4471
rect 3835 4437 3844 4471
rect 3792 4428 3844 4437
rect 4922 4326 4974 4378
rect 4986 4326 5038 4378
rect 5050 4326 5102 4378
rect 5114 4326 5166 4378
rect 5178 4326 5230 4378
rect 5242 4326 5294 4378
rect 6736 4224 6788 4276
rect 1400 4199 1452 4208
rect 1400 4165 1409 4199
rect 1409 4165 1443 4199
rect 1443 4165 1452 4199
rect 1400 4156 1452 4165
rect 4620 4156 4672 4208
rect 6184 4131 6236 4140
rect 6184 4097 6193 4131
rect 6193 4097 6227 4131
rect 6227 4097 6236 4131
rect 6184 4088 6236 4097
rect 5816 4020 5868 4072
rect 6644 4088 6696 4140
rect 6552 4020 6604 4072
rect 7104 3952 7156 4004
rect 4620 3884 4672 3936
rect 5908 3884 5960 3936
rect 4182 3782 4234 3834
rect 4246 3782 4298 3834
rect 4310 3782 4362 3834
rect 4374 3782 4426 3834
rect 4438 3782 4490 3834
rect 4502 3782 4554 3834
rect 5448 3544 5500 3596
rect 6736 3680 6788 3732
rect 6828 3587 6880 3596
rect 6828 3553 6837 3587
rect 6837 3553 6871 3587
rect 6871 3553 6880 3587
rect 6828 3544 6880 3553
rect 7104 3587 7156 3596
rect 7104 3553 7113 3587
rect 7113 3553 7147 3587
rect 7147 3553 7156 3587
rect 7104 3544 7156 3553
rect 4804 3408 4856 3460
rect 4620 3340 4672 3392
rect 6736 3340 6788 3392
rect 4922 3238 4974 3290
rect 4986 3238 5038 3290
rect 5050 3238 5102 3290
rect 5114 3238 5166 3290
rect 5178 3238 5230 3290
rect 5242 3238 5294 3290
rect 5816 3136 5868 3188
rect 6644 3136 6696 3188
rect 5908 3111 5960 3120
rect 5908 3077 5917 3111
rect 5917 3077 5951 3111
rect 5951 3077 5960 3111
rect 5908 3068 5960 3077
rect 6736 3111 6788 3120
rect 6736 3077 6745 3111
rect 6745 3077 6779 3111
rect 6779 3077 6788 3111
rect 6736 3068 6788 3077
rect 4620 3000 4672 3052
rect 4804 3000 4856 3052
rect 6184 3043 6236 3052
rect 6184 3009 6193 3043
rect 6193 3009 6227 3043
rect 6227 3009 6236 3043
rect 6184 3000 6236 3009
rect 6552 2932 6604 2984
rect 7564 2864 7616 2916
rect 4620 2796 4672 2848
rect 6644 2796 6696 2848
rect 4182 2694 4234 2746
rect 4246 2694 4298 2746
rect 4310 2694 4362 2746
rect 4374 2694 4426 2746
rect 4438 2694 4490 2746
rect 4502 2694 4554 2746
rect 4436 2567 4488 2576
rect 4436 2533 4445 2567
rect 4445 2533 4479 2567
rect 4479 2533 4488 2567
rect 4436 2524 4488 2533
rect 7196 2592 7248 2644
rect 6184 2499 6236 2508
rect 6184 2465 6193 2499
rect 6193 2465 6227 2499
rect 6227 2465 6236 2499
rect 6184 2456 6236 2465
rect 6552 2456 6604 2508
rect 4620 2388 4672 2440
rect 4804 2388 4856 2440
rect 6460 2388 6512 2440
rect 4436 2320 4488 2372
rect 7380 2320 7432 2372
rect 6736 2252 6788 2304
rect 4922 2150 4974 2202
rect 4986 2150 5038 2202
rect 5050 2150 5102 2202
rect 5114 2150 5166 2202
rect 5178 2150 5230 2202
rect 5242 2150 5294 2202
rect 4436 2048 4488 2100
rect 6460 2048 6512 2100
<< metal2 >>
rect 6826 9888 6882 9897
rect 6826 9823 6882 9832
rect 1306 9616 1362 9625
rect 1306 9551 1362 9560
rect 1320 8498 1348 9551
rect 4920 8732 5296 8741
rect 4976 8730 5000 8732
rect 5056 8730 5080 8732
rect 5136 8730 5160 8732
rect 5216 8730 5240 8732
rect 4976 8678 4986 8730
rect 5230 8678 5240 8730
rect 4976 8676 5000 8678
rect 5056 8676 5080 8678
rect 5136 8676 5160 8678
rect 5216 8676 5240 8678
rect 4920 8667 5296 8676
rect 6840 8566 6868 9823
rect 7378 8800 7434 8809
rect 7378 8735 7434 8744
rect 7392 8566 7420 8735
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 7380 8560 7432 8566
rect 7380 8502 7432 8508
rect 1308 8492 1360 8498
rect 1308 8434 1360 8440
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2884 7886 2912 8298
rect 4180 8188 4556 8197
rect 4236 8186 4260 8188
rect 4316 8186 4340 8188
rect 4396 8186 4420 8188
rect 4476 8186 4500 8188
rect 4236 8134 4246 8186
rect 4490 8134 4500 8186
rect 4236 8132 4260 8134
rect 4316 8132 4340 8134
rect 4396 8132 4420 8134
rect 4476 8132 4500 8134
rect 4180 8123 4556 8132
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 1584 7812 1636 7818
rect 1584 7754 1636 7760
rect 2964 7812 3016 7818
rect 2964 7754 3016 7760
rect 5816 7812 5868 7818
rect 5816 7754 5868 7760
rect 1492 7336 1544 7342
rect 1492 7278 1544 7284
rect 1306 6896 1362 6905
rect 1504 6866 1532 7278
rect 1596 7002 1624 7754
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 1780 7478 1808 7686
rect 2516 7546 2544 7686
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 1768 7472 1820 7478
rect 1768 7414 1820 7420
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1306 6831 1362 6840
rect 1492 6860 1544 6866
rect 1320 6798 1348 6831
rect 1492 6802 1544 6808
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 1308 6792 1360 6798
rect 1308 6734 1360 6740
rect 1860 6724 1912 6730
rect 1860 6666 1912 6672
rect 1872 6254 1900 6666
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2240 6322 2268 6598
rect 2700 6322 2728 6802
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 1780 5914 1808 6054
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 2700 5778 2728 6258
rect 1676 5772 1728 5778
rect 1676 5714 1728 5720
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 1688 5234 1716 5714
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 1964 4826 1992 5102
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 2976 4690 3004 7754
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 4920 7644 5296 7653
rect 4976 7642 5000 7644
rect 5056 7642 5080 7644
rect 5136 7642 5160 7644
rect 5216 7642 5240 7644
rect 4976 7590 4986 7642
rect 5230 7590 5240 7642
rect 4976 7588 5000 7590
rect 5056 7588 5080 7590
rect 5136 7588 5160 7590
rect 5216 7588 5240 7590
rect 4920 7579 5296 7588
rect 3240 7472 3292 7478
rect 3240 7414 3292 7420
rect 3252 6798 3280 7414
rect 4620 7336 4672 7342
rect 4672 7284 4752 7290
rect 4620 7278 4752 7284
rect 4632 7262 4752 7278
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4180 7100 4556 7109
rect 4236 7098 4260 7100
rect 4316 7098 4340 7100
rect 4396 7098 4420 7100
rect 4476 7098 4500 7100
rect 4236 7046 4246 7098
rect 4490 7046 4500 7098
rect 4236 7044 4260 7046
rect 4316 7044 4340 7046
rect 4396 7044 4420 7046
rect 4476 7044 4500 7046
rect 4180 7035 4556 7044
rect 4632 6914 4660 7142
rect 4724 7002 4752 7262
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 4448 6886 4660 6914
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3252 6118 3280 6734
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3252 5710 3280 6054
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3620 5234 3648 6802
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3896 6254 3924 6734
rect 4448 6322 4476 6886
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 4920 6556 5296 6565
rect 4976 6554 5000 6556
rect 5056 6554 5080 6556
rect 5136 6554 5160 6556
rect 5216 6554 5240 6556
rect 4976 6502 4986 6554
rect 5230 6502 5240 6554
rect 4976 6500 5000 6502
rect 5056 6500 5080 6502
rect 5136 6500 5160 6502
rect 5216 6500 5240 6502
rect 4920 6491 5296 6500
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3896 5846 3924 6190
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 4080 5914 4108 6122
rect 4180 6012 4556 6021
rect 4236 6010 4260 6012
rect 4316 6010 4340 6012
rect 4396 6010 4420 6012
rect 4476 6010 4500 6012
rect 4236 5958 4246 6010
rect 4490 5958 4500 6010
rect 4236 5956 4260 5958
rect 4316 5956 4340 5958
rect 4396 5956 4420 5958
rect 4476 5956 4500 5958
rect 4180 5947 4556 5956
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3884 5840 3936 5846
rect 3884 5782 3936 5788
rect 4068 5772 4120 5778
rect 3988 5732 4068 5760
rect 3988 5642 4016 5732
rect 4068 5714 4120 5720
rect 3976 5636 4028 5642
rect 3976 5578 4028 5584
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4620 5636 4672 5642
rect 4620 5578 4672 5584
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 3436 4622 3464 4966
rect 3620 4758 3648 5170
rect 3608 4752 3660 4758
rect 3608 4694 3660 4700
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 1412 4214 1440 4558
rect 3804 4486 3832 5170
rect 3988 4690 4016 5578
rect 4172 5030 4200 5578
rect 4632 5370 4660 5578
rect 4816 5370 4844 6326
rect 5368 5778 5396 6598
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5736 5642 5764 7686
rect 5828 7410 5856 7754
rect 6000 7472 6052 7478
rect 6000 7414 6052 7420
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 6012 6474 6040 7414
rect 6564 7342 6592 8434
rect 6656 7546 6684 8434
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6748 7274 6776 7890
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6104 7002 6132 7142
rect 6092 6996 6144 7002
rect 6092 6938 6144 6944
rect 6012 6446 6132 6474
rect 6104 6390 6132 6446
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6092 6384 6144 6390
rect 6092 6326 6144 6332
rect 6104 6118 6132 6326
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6104 5642 6132 6054
rect 5724 5636 5776 5642
rect 5724 5578 5776 5584
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 5906 5536 5962 5545
rect 4920 5468 5296 5477
rect 5906 5471 5962 5480
rect 4976 5466 5000 5468
rect 5056 5466 5080 5468
rect 5136 5466 5160 5468
rect 5216 5466 5240 5468
rect 4976 5414 4986 5466
rect 5230 5414 5240 5466
rect 4976 5412 5000 5414
rect 5056 5412 5080 5414
rect 5136 5412 5160 5414
rect 5216 5412 5240 5414
rect 4920 5403 5296 5412
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4180 4924 4556 4933
rect 4236 4922 4260 4924
rect 4316 4922 4340 4924
rect 4396 4922 4420 4924
rect 4476 4922 4500 4924
rect 4236 4870 4246 4922
rect 4490 4870 4500 4922
rect 4236 4868 4260 4870
rect 4316 4868 4340 4870
rect 4396 4868 4420 4870
rect 4476 4868 4500 4870
rect 4180 4859 4556 4868
rect 3976 4684 4028 4690
rect 3976 4626 4028 4632
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 1400 4208 1452 4214
rect 1398 4176 1400 4185
rect 1452 4176 1454 4185
rect 1398 4111 1454 4120
rect 3804 1465 3832 4422
rect 4632 4214 4660 5306
rect 4816 4622 4844 5306
rect 5920 5302 5948 5471
rect 5908 5296 5960 5302
rect 5908 5238 5960 5244
rect 6564 5166 6592 6190
rect 6656 5370 6684 6394
rect 6748 6254 6776 7210
rect 6840 6798 6868 7754
rect 6920 7744 6972 7750
rect 7392 7721 7420 7754
rect 6920 7686 6972 7692
rect 7378 7712 7434 7721
rect 6932 7410 6960 7686
rect 7378 7647 7434 7656
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6932 7002 6960 7346
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6840 6458 6868 6734
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 7392 6633 7420 6666
rect 7378 6624 7434 6633
rect 7378 6559 7434 6568
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6840 5914 6868 6394
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 5446 4448 5502 4457
rect 4920 4380 5296 4389
rect 5446 4383 5502 4392
rect 4976 4378 5000 4380
rect 5056 4378 5080 4380
rect 5136 4378 5160 4380
rect 5216 4378 5240 4380
rect 4976 4326 4986 4378
rect 5230 4326 5240 4378
rect 4976 4324 5000 4326
rect 5056 4324 5080 4326
rect 5136 4324 5160 4326
rect 5216 4324 5240 4326
rect 4920 4315 5296 4324
rect 4620 4208 4672 4214
rect 4672 4156 4844 4162
rect 4620 4150 4844 4156
rect 4632 4134 4844 4150
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4180 3836 4556 3845
rect 4236 3834 4260 3836
rect 4316 3834 4340 3836
rect 4396 3834 4420 3836
rect 4476 3834 4500 3836
rect 4236 3782 4246 3834
rect 4490 3782 4500 3834
rect 4236 3780 4260 3782
rect 4316 3780 4340 3782
rect 4396 3780 4420 3782
rect 4476 3780 4500 3782
rect 4180 3771 4556 3780
rect 4632 3398 4660 3878
rect 4816 3466 4844 4134
rect 5460 3602 5488 4383
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4632 3058 4660 3334
rect 4816 3058 4844 3402
rect 4920 3292 5296 3301
rect 4976 3290 5000 3292
rect 5056 3290 5080 3292
rect 5136 3290 5160 3292
rect 5216 3290 5240 3292
rect 4976 3238 4986 3290
rect 5230 3238 5240 3290
rect 4976 3236 5000 3238
rect 5056 3236 5080 3238
rect 5136 3236 5160 3238
rect 5216 3236 5240 3238
rect 4920 3227 5296 3236
rect 5828 3194 5856 4014
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5920 3126 5948 3878
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 6196 3058 6224 4082
rect 6564 4078 6592 5102
rect 6748 4282 6776 5170
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4180 2748 4556 2757
rect 4236 2746 4260 2748
rect 4316 2746 4340 2748
rect 4396 2746 4420 2748
rect 4476 2746 4500 2748
rect 4236 2694 4246 2746
rect 4490 2694 4500 2746
rect 4236 2692 4260 2694
rect 4316 2692 4340 2694
rect 4396 2692 4420 2694
rect 4476 2692 4500 2694
rect 4180 2683 4556 2692
rect 4436 2576 4488 2582
rect 4436 2518 4488 2524
rect 4448 2378 4476 2518
rect 4632 2446 4660 2790
rect 4816 2446 4844 2994
rect 6196 2514 6224 2994
rect 6564 2990 6592 4014
rect 6656 3194 6684 4082
rect 6748 3738 6776 4218
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6840 3602 6868 4966
rect 7116 4826 7144 5714
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7116 4010 7144 4762
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 7116 3602 7144 3946
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 7194 3360 7250 3369
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6564 2514 6592 2926
rect 6656 2854 6684 3130
rect 6748 3126 6776 3334
rect 7194 3295 7250 3304
rect 6736 3120 6788 3126
rect 6736 3062 6788 3068
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 4436 2372 4488 2378
rect 4436 2314 4488 2320
rect 4448 2106 4476 2314
rect 4920 2204 5296 2213
rect 4976 2202 5000 2204
rect 5056 2202 5080 2204
rect 5136 2202 5160 2204
rect 5216 2202 5240 2204
rect 4976 2150 4986 2202
rect 5230 2150 5240 2202
rect 4976 2148 5000 2150
rect 5056 2148 5080 2150
rect 5136 2148 5160 2150
rect 5216 2148 5240 2150
rect 4920 2139 5296 2148
rect 6472 2106 6500 2382
rect 6748 2310 6776 3062
rect 7208 2650 7236 3295
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7380 2372 7432 2378
rect 7380 2314 7432 2320
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 4436 2100 4488 2106
rect 4436 2042 4488 2048
rect 6460 2100 6512 2106
rect 6460 2042 6512 2048
rect 3790 1456 3846 1465
rect 3790 1391 3846 1400
rect 7392 1193 7420 2314
rect 7576 2281 7604 2858
rect 7562 2272 7618 2281
rect 7562 2207 7618 2216
rect 7378 1184 7434 1193
rect 7378 1119 7434 1128
<< via2 >>
rect 6826 9832 6882 9888
rect 1306 9560 1362 9616
rect 4920 8730 4976 8732
rect 5000 8730 5056 8732
rect 5080 8730 5136 8732
rect 5160 8730 5216 8732
rect 5240 8730 5296 8732
rect 4920 8678 4922 8730
rect 4922 8678 4974 8730
rect 4974 8678 4976 8730
rect 5000 8678 5038 8730
rect 5038 8678 5050 8730
rect 5050 8678 5056 8730
rect 5080 8678 5102 8730
rect 5102 8678 5114 8730
rect 5114 8678 5136 8730
rect 5160 8678 5166 8730
rect 5166 8678 5178 8730
rect 5178 8678 5216 8730
rect 5240 8678 5242 8730
rect 5242 8678 5294 8730
rect 5294 8678 5296 8730
rect 4920 8676 4976 8678
rect 5000 8676 5056 8678
rect 5080 8676 5136 8678
rect 5160 8676 5216 8678
rect 5240 8676 5296 8678
rect 7378 8744 7434 8800
rect 4180 8186 4236 8188
rect 4260 8186 4316 8188
rect 4340 8186 4396 8188
rect 4420 8186 4476 8188
rect 4500 8186 4556 8188
rect 4180 8134 4182 8186
rect 4182 8134 4234 8186
rect 4234 8134 4236 8186
rect 4260 8134 4298 8186
rect 4298 8134 4310 8186
rect 4310 8134 4316 8186
rect 4340 8134 4362 8186
rect 4362 8134 4374 8186
rect 4374 8134 4396 8186
rect 4420 8134 4426 8186
rect 4426 8134 4438 8186
rect 4438 8134 4476 8186
rect 4500 8134 4502 8186
rect 4502 8134 4554 8186
rect 4554 8134 4556 8186
rect 4180 8132 4236 8134
rect 4260 8132 4316 8134
rect 4340 8132 4396 8134
rect 4420 8132 4476 8134
rect 4500 8132 4556 8134
rect 1306 6840 1362 6896
rect 4920 7642 4976 7644
rect 5000 7642 5056 7644
rect 5080 7642 5136 7644
rect 5160 7642 5216 7644
rect 5240 7642 5296 7644
rect 4920 7590 4922 7642
rect 4922 7590 4974 7642
rect 4974 7590 4976 7642
rect 5000 7590 5038 7642
rect 5038 7590 5050 7642
rect 5050 7590 5056 7642
rect 5080 7590 5102 7642
rect 5102 7590 5114 7642
rect 5114 7590 5136 7642
rect 5160 7590 5166 7642
rect 5166 7590 5178 7642
rect 5178 7590 5216 7642
rect 5240 7590 5242 7642
rect 5242 7590 5294 7642
rect 5294 7590 5296 7642
rect 4920 7588 4976 7590
rect 5000 7588 5056 7590
rect 5080 7588 5136 7590
rect 5160 7588 5216 7590
rect 5240 7588 5296 7590
rect 4180 7098 4236 7100
rect 4260 7098 4316 7100
rect 4340 7098 4396 7100
rect 4420 7098 4476 7100
rect 4500 7098 4556 7100
rect 4180 7046 4182 7098
rect 4182 7046 4234 7098
rect 4234 7046 4236 7098
rect 4260 7046 4298 7098
rect 4298 7046 4310 7098
rect 4310 7046 4316 7098
rect 4340 7046 4362 7098
rect 4362 7046 4374 7098
rect 4374 7046 4396 7098
rect 4420 7046 4426 7098
rect 4426 7046 4438 7098
rect 4438 7046 4476 7098
rect 4500 7046 4502 7098
rect 4502 7046 4554 7098
rect 4554 7046 4556 7098
rect 4180 7044 4236 7046
rect 4260 7044 4316 7046
rect 4340 7044 4396 7046
rect 4420 7044 4476 7046
rect 4500 7044 4556 7046
rect 4920 6554 4976 6556
rect 5000 6554 5056 6556
rect 5080 6554 5136 6556
rect 5160 6554 5216 6556
rect 5240 6554 5296 6556
rect 4920 6502 4922 6554
rect 4922 6502 4974 6554
rect 4974 6502 4976 6554
rect 5000 6502 5038 6554
rect 5038 6502 5050 6554
rect 5050 6502 5056 6554
rect 5080 6502 5102 6554
rect 5102 6502 5114 6554
rect 5114 6502 5136 6554
rect 5160 6502 5166 6554
rect 5166 6502 5178 6554
rect 5178 6502 5216 6554
rect 5240 6502 5242 6554
rect 5242 6502 5294 6554
rect 5294 6502 5296 6554
rect 4920 6500 4976 6502
rect 5000 6500 5056 6502
rect 5080 6500 5136 6502
rect 5160 6500 5216 6502
rect 5240 6500 5296 6502
rect 4180 6010 4236 6012
rect 4260 6010 4316 6012
rect 4340 6010 4396 6012
rect 4420 6010 4476 6012
rect 4500 6010 4556 6012
rect 4180 5958 4182 6010
rect 4182 5958 4234 6010
rect 4234 5958 4236 6010
rect 4260 5958 4298 6010
rect 4298 5958 4310 6010
rect 4310 5958 4316 6010
rect 4340 5958 4362 6010
rect 4362 5958 4374 6010
rect 4374 5958 4396 6010
rect 4420 5958 4426 6010
rect 4426 5958 4438 6010
rect 4438 5958 4476 6010
rect 4500 5958 4502 6010
rect 4502 5958 4554 6010
rect 4554 5958 4556 6010
rect 4180 5956 4236 5958
rect 4260 5956 4316 5958
rect 4340 5956 4396 5958
rect 4420 5956 4476 5958
rect 4500 5956 4556 5958
rect 5906 5480 5962 5536
rect 4920 5466 4976 5468
rect 5000 5466 5056 5468
rect 5080 5466 5136 5468
rect 5160 5466 5216 5468
rect 5240 5466 5296 5468
rect 4920 5414 4922 5466
rect 4922 5414 4974 5466
rect 4974 5414 4976 5466
rect 5000 5414 5038 5466
rect 5038 5414 5050 5466
rect 5050 5414 5056 5466
rect 5080 5414 5102 5466
rect 5102 5414 5114 5466
rect 5114 5414 5136 5466
rect 5160 5414 5166 5466
rect 5166 5414 5178 5466
rect 5178 5414 5216 5466
rect 5240 5414 5242 5466
rect 5242 5414 5294 5466
rect 5294 5414 5296 5466
rect 4920 5412 4976 5414
rect 5000 5412 5056 5414
rect 5080 5412 5136 5414
rect 5160 5412 5216 5414
rect 5240 5412 5296 5414
rect 4180 4922 4236 4924
rect 4260 4922 4316 4924
rect 4340 4922 4396 4924
rect 4420 4922 4476 4924
rect 4500 4922 4556 4924
rect 4180 4870 4182 4922
rect 4182 4870 4234 4922
rect 4234 4870 4236 4922
rect 4260 4870 4298 4922
rect 4298 4870 4310 4922
rect 4310 4870 4316 4922
rect 4340 4870 4362 4922
rect 4362 4870 4374 4922
rect 4374 4870 4396 4922
rect 4420 4870 4426 4922
rect 4426 4870 4438 4922
rect 4438 4870 4476 4922
rect 4500 4870 4502 4922
rect 4502 4870 4554 4922
rect 4554 4870 4556 4922
rect 4180 4868 4236 4870
rect 4260 4868 4316 4870
rect 4340 4868 4396 4870
rect 4420 4868 4476 4870
rect 4500 4868 4556 4870
rect 1398 4156 1400 4176
rect 1400 4156 1452 4176
rect 1452 4156 1454 4176
rect 1398 4120 1454 4156
rect 7378 7656 7434 7712
rect 7378 6568 7434 6624
rect 5446 4392 5502 4448
rect 4920 4378 4976 4380
rect 5000 4378 5056 4380
rect 5080 4378 5136 4380
rect 5160 4378 5216 4380
rect 5240 4378 5296 4380
rect 4920 4326 4922 4378
rect 4922 4326 4974 4378
rect 4974 4326 4976 4378
rect 5000 4326 5038 4378
rect 5038 4326 5050 4378
rect 5050 4326 5056 4378
rect 5080 4326 5102 4378
rect 5102 4326 5114 4378
rect 5114 4326 5136 4378
rect 5160 4326 5166 4378
rect 5166 4326 5178 4378
rect 5178 4326 5216 4378
rect 5240 4326 5242 4378
rect 5242 4326 5294 4378
rect 5294 4326 5296 4378
rect 4920 4324 4976 4326
rect 5000 4324 5056 4326
rect 5080 4324 5136 4326
rect 5160 4324 5216 4326
rect 5240 4324 5296 4326
rect 4180 3834 4236 3836
rect 4260 3834 4316 3836
rect 4340 3834 4396 3836
rect 4420 3834 4476 3836
rect 4500 3834 4556 3836
rect 4180 3782 4182 3834
rect 4182 3782 4234 3834
rect 4234 3782 4236 3834
rect 4260 3782 4298 3834
rect 4298 3782 4310 3834
rect 4310 3782 4316 3834
rect 4340 3782 4362 3834
rect 4362 3782 4374 3834
rect 4374 3782 4396 3834
rect 4420 3782 4426 3834
rect 4426 3782 4438 3834
rect 4438 3782 4476 3834
rect 4500 3782 4502 3834
rect 4502 3782 4554 3834
rect 4554 3782 4556 3834
rect 4180 3780 4236 3782
rect 4260 3780 4316 3782
rect 4340 3780 4396 3782
rect 4420 3780 4476 3782
rect 4500 3780 4556 3782
rect 4920 3290 4976 3292
rect 5000 3290 5056 3292
rect 5080 3290 5136 3292
rect 5160 3290 5216 3292
rect 5240 3290 5296 3292
rect 4920 3238 4922 3290
rect 4922 3238 4974 3290
rect 4974 3238 4976 3290
rect 5000 3238 5038 3290
rect 5038 3238 5050 3290
rect 5050 3238 5056 3290
rect 5080 3238 5102 3290
rect 5102 3238 5114 3290
rect 5114 3238 5136 3290
rect 5160 3238 5166 3290
rect 5166 3238 5178 3290
rect 5178 3238 5216 3290
rect 5240 3238 5242 3290
rect 5242 3238 5294 3290
rect 5294 3238 5296 3290
rect 4920 3236 4976 3238
rect 5000 3236 5056 3238
rect 5080 3236 5136 3238
rect 5160 3236 5216 3238
rect 5240 3236 5296 3238
rect 4180 2746 4236 2748
rect 4260 2746 4316 2748
rect 4340 2746 4396 2748
rect 4420 2746 4476 2748
rect 4500 2746 4556 2748
rect 4180 2694 4182 2746
rect 4182 2694 4234 2746
rect 4234 2694 4236 2746
rect 4260 2694 4298 2746
rect 4298 2694 4310 2746
rect 4310 2694 4316 2746
rect 4340 2694 4362 2746
rect 4362 2694 4374 2746
rect 4374 2694 4396 2746
rect 4420 2694 4426 2746
rect 4426 2694 4438 2746
rect 4438 2694 4476 2746
rect 4500 2694 4502 2746
rect 4502 2694 4554 2746
rect 4554 2694 4556 2746
rect 4180 2692 4236 2694
rect 4260 2692 4316 2694
rect 4340 2692 4396 2694
rect 4420 2692 4476 2694
rect 4500 2692 4556 2694
rect 7194 3304 7250 3360
rect 4920 2202 4976 2204
rect 5000 2202 5056 2204
rect 5080 2202 5136 2204
rect 5160 2202 5216 2204
rect 5240 2202 5296 2204
rect 4920 2150 4922 2202
rect 4922 2150 4974 2202
rect 4974 2150 4976 2202
rect 5000 2150 5038 2202
rect 5038 2150 5050 2202
rect 5050 2150 5056 2202
rect 5080 2150 5102 2202
rect 5102 2150 5114 2202
rect 5114 2150 5136 2202
rect 5160 2150 5166 2202
rect 5166 2150 5178 2202
rect 5178 2150 5216 2202
rect 5240 2150 5242 2202
rect 5242 2150 5294 2202
rect 5294 2150 5296 2202
rect 4920 2148 4976 2150
rect 5000 2148 5056 2150
rect 5080 2148 5136 2150
rect 5160 2148 5216 2150
rect 5240 2148 5296 2150
rect 3790 1400 3846 1456
rect 7562 2216 7618 2272
rect 7378 1128 7434 1184
<< metal3 >>
rect 6821 9890 6887 9893
rect 8249 9890 9049 9920
rect 6821 9888 9049 9890
rect 6821 9832 6826 9888
rect 6882 9832 9049 9888
rect 6821 9830 9049 9832
rect 6821 9827 6887 9830
rect 8249 9800 9049 9830
rect 0 9618 800 9648
rect 1301 9618 1367 9621
rect 0 9616 1367 9618
rect 0 9560 1306 9616
rect 1362 9560 1367 9616
rect 0 9558 1367 9560
rect 0 9528 800 9558
rect 1301 9555 1367 9558
rect 7373 8802 7439 8805
rect 8249 8802 9049 8832
rect 7373 8800 9049 8802
rect 7373 8744 7378 8800
rect 7434 8744 9049 8800
rect 7373 8742 9049 8744
rect 7373 8739 7439 8742
rect 4910 8736 5306 8737
rect 4910 8672 4916 8736
rect 4980 8672 4996 8736
rect 5060 8672 5076 8736
rect 5140 8672 5156 8736
rect 5220 8672 5236 8736
rect 5300 8672 5306 8736
rect 8249 8712 9049 8742
rect 4910 8671 5306 8672
rect 4170 8192 4566 8193
rect 4170 8128 4176 8192
rect 4240 8128 4256 8192
rect 4320 8128 4336 8192
rect 4400 8128 4416 8192
rect 4480 8128 4496 8192
rect 4560 8128 4566 8192
rect 4170 8127 4566 8128
rect 7373 7714 7439 7717
rect 8249 7714 9049 7744
rect 7373 7712 9049 7714
rect 7373 7656 7378 7712
rect 7434 7656 9049 7712
rect 7373 7654 9049 7656
rect 7373 7651 7439 7654
rect 4910 7648 5306 7649
rect 4910 7584 4916 7648
rect 4980 7584 4996 7648
rect 5060 7584 5076 7648
rect 5140 7584 5156 7648
rect 5220 7584 5236 7648
rect 5300 7584 5306 7648
rect 8249 7624 9049 7654
rect 4910 7583 5306 7584
rect 4170 7104 4566 7105
rect 4170 7040 4176 7104
rect 4240 7040 4256 7104
rect 4320 7040 4336 7104
rect 4400 7040 4416 7104
rect 4480 7040 4496 7104
rect 4560 7040 4566 7104
rect 4170 7039 4566 7040
rect 0 6898 800 6928
rect 1301 6898 1367 6901
rect 0 6896 1367 6898
rect 0 6840 1306 6896
rect 1362 6840 1367 6896
rect 0 6838 1367 6840
rect 0 6808 800 6838
rect 1301 6835 1367 6838
rect 7373 6626 7439 6629
rect 8249 6626 9049 6656
rect 7373 6624 9049 6626
rect 7373 6568 7378 6624
rect 7434 6568 9049 6624
rect 7373 6566 9049 6568
rect 7373 6563 7439 6566
rect 4910 6560 5306 6561
rect 4910 6496 4916 6560
rect 4980 6496 4996 6560
rect 5060 6496 5076 6560
rect 5140 6496 5156 6560
rect 5220 6496 5236 6560
rect 5300 6496 5306 6560
rect 8249 6536 9049 6566
rect 4910 6495 5306 6496
rect 4170 6016 4566 6017
rect 4170 5952 4176 6016
rect 4240 5952 4256 6016
rect 4320 5952 4336 6016
rect 4400 5952 4416 6016
rect 4480 5952 4496 6016
rect 4560 5952 4566 6016
rect 4170 5951 4566 5952
rect 5901 5538 5967 5541
rect 8249 5538 9049 5568
rect 5901 5536 9049 5538
rect 5901 5480 5906 5536
rect 5962 5480 9049 5536
rect 5901 5478 9049 5480
rect 5901 5475 5967 5478
rect 4910 5472 5306 5473
rect 4910 5408 4916 5472
rect 4980 5408 4996 5472
rect 5060 5408 5076 5472
rect 5140 5408 5156 5472
rect 5220 5408 5236 5472
rect 5300 5408 5306 5472
rect 8249 5448 9049 5478
rect 4910 5407 5306 5408
rect 4170 4928 4566 4929
rect 4170 4864 4176 4928
rect 4240 4864 4256 4928
rect 4320 4864 4336 4928
rect 4400 4864 4416 4928
rect 4480 4864 4496 4928
rect 4560 4864 4566 4928
rect 4170 4863 4566 4864
rect 5441 4450 5507 4453
rect 8249 4450 9049 4480
rect 5441 4448 9049 4450
rect 5441 4392 5446 4448
rect 5502 4392 9049 4448
rect 5441 4390 9049 4392
rect 5441 4387 5507 4390
rect 4910 4384 5306 4385
rect 4910 4320 4916 4384
rect 4980 4320 4996 4384
rect 5060 4320 5076 4384
rect 5140 4320 5156 4384
rect 5220 4320 5236 4384
rect 5300 4320 5306 4384
rect 8249 4360 9049 4390
rect 4910 4319 5306 4320
rect 0 4178 800 4208
rect 1393 4178 1459 4181
rect 0 4176 1459 4178
rect 0 4120 1398 4176
rect 1454 4120 1459 4176
rect 0 4118 1459 4120
rect 0 4088 800 4118
rect 1393 4115 1459 4118
rect 4170 3840 4566 3841
rect 4170 3776 4176 3840
rect 4240 3776 4256 3840
rect 4320 3776 4336 3840
rect 4400 3776 4416 3840
rect 4480 3776 4496 3840
rect 4560 3776 4566 3840
rect 4170 3775 4566 3776
rect 7189 3362 7255 3365
rect 8249 3362 9049 3392
rect 7189 3360 9049 3362
rect 7189 3304 7194 3360
rect 7250 3304 9049 3360
rect 7189 3302 9049 3304
rect 7189 3299 7255 3302
rect 4910 3296 5306 3297
rect 4910 3232 4916 3296
rect 4980 3232 4996 3296
rect 5060 3232 5076 3296
rect 5140 3232 5156 3296
rect 5220 3232 5236 3296
rect 5300 3232 5306 3296
rect 8249 3272 9049 3302
rect 4910 3231 5306 3232
rect 4170 2752 4566 2753
rect 4170 2688 4176 2752
rect 4240 2688 4256 2752
rect 4320 2688 4336 2752
rect 4400 2688 4416 2752
rect 4480 2688 4496 2752
rect 4560 2688 4566 2752
rect 4170 2687 4566 2688
rect 7557 2274 7623 2277
rect 8249 2274 9049 2304
rect 7557 2272 9049 2274
rect 7557 2216 7562 2272
rect 7618 2216 9049 2272
rect 7557 2214 9049 2216
rect 7557 2211 7623 2214
rect 4910 2208 5306 2209
rect 4910 2144 4916 2208
rect 4980 2144 4996 2208
rect 5060 2144 5076 2208
rect 5140 2144 5156 2208
rect 5220 2144 5236 2208
rect 5300 2144 5306 2208
rect 8249 2184 9049 2214
rect 4910 2143 5306 2144
rect 0 1458 800 1488
rect 3785 1458 3851 1461
rect 0 1456 3851 1458
rect 0 1400 3790 1456
rect 3846 1400 3851 1456
rect 0 1398 3851 1400
rect 0 1368 800 1398
rect 3785 1395 3851 1398
rect 7373 1186 7439 1189
rect 8249 1186 9049 1216
rect 7373 1184 9049 1186
rect 7373 1128 7378 1184
rect 7434 1128 9049 1184
rect 7373 1126 9049 1128
rect 7373 1123 7439 1126
rect 8249 1096 9049 1126
<< via3 >>
rect 4916 8732 4980 8736
rect 4916 8676 4920 8732
rect 4920 8676 4976 8732
rect 4976 8676 4980 8732
rect 4916 8672 4980 8676
rect 4996 8732 5060 8736
rect 4996 8676 5000 8732
rect 5000 8676 5056 8732
rect 5056 8676 5060 8732
rect 4996 8672 5060 8676
rect 5076 8732 5140 8736
rect 5076 8676 5080 8732
rect 5080 8676 5136 8732
rect 5136 8676 5140 8732
rect 5076 8672 5140 8676
rect 5156 8732 5220 8736
rect 5156 8676 5160 8732
rect 5160 8676 5216 8732
rect 5216 8676 5220 8732
rect 5156 8672 5220 8676
rect 5236 8732 5300 8736
rect 5236 8676 5240 8732
rect 5240 8676 5296 8732
rect 5296 8676 5300 8732
rect 5236 8672 5300 8676
rect 4176 8188 4240 8192
rect 4176 8132 4180 8188
rect 4180 8132 4236 8188
rect 4236 8132 4240 8188
rect 4176 8128 4240 8132
rect 4256 8188 4320 8192
rect 4256 8132 4260 8188
rect 4260 8132 4316 8188
rect 4316 8132 4320 8188
rect 4256 8128 4320 8132
rect 4336 8188 4400 8192
rect 4336 8132 4340 8188
rect 4340 8132 4396 8188
rect 4396 8132 4400 8188
rect 4336 8128 4400 8132
rect 4416 8188 4480 8192
rect 4416 8132 4420 8188
rect 4420 8132 4476 8188
rect 4476 8132 4480 8188
rect 4416 8128 4480 8132
rect 4496 8188 4560 8192
rect 4496 8132 4500 8188
rect 4500 8132 4556 8188
rect 4556 8132 4560 8188
rect 4496 8128 4560 8132
rect 4916 7644 4980 7648
rect 4916 7588 4920 7644
rect 4920 7588 4976 7644
rect 4976 7588 4980 7644
rect 4916 7584 4980 7588
rect 4996 7644 5060 7648
rect 4996 7588 5000 7644
rect 5000 7588 5056 7644
rect 5056 7588 5060 7644
rect 4996 7584 5060 7588
rect 5076 7644 5140 7648
rect 5076 7588 5080 7644
rect 5080 7588 5136 7644
rect 5136 7588 5140 7644
rect 5076 7584 5140 7588
rect 5156 7644 5220 7648
rect 5156 7588 5160 7644
rect 5160 7588 5216 7644
rect 5216 7588 5220 7644
rect 5156 7584 5220 7588
rect 5236 7644 5300 7648
rect 5236 7588 5240 7644
rect 5240 7588 5296 7644
rect 5296 7588 5300 7644
rect 5236 7584 5300 7588
rect 4176 7100 4240 7104
rect 4176 7044 4180 7100
rect 4180 7044 4236 7100
rect 4236 7044 4240 7100
rect 4176 7040 4240 7044
rect 4256 7100 4320 7104
rect 4256 7044 4260 7100
rect 4260 7044 4316 7100
rect 4316 7044 4320 7100
rect 4256 7040 4320 7044
rect 4336 7100 4400 7104
rect 4336 7044 4340 7100
rect 4340 7044 4396 7100
rect 4396 7044 4400 7100
rect 4336 7040 4400 7044
rect 4416 7100 4480 7104
rect 4416 7044 4420 7100
rect 4420 7044 4476 7100
rect 4476 7044 4480 7100
rect 4416 7040 4480 7044
rect 4496 7100 4560 7104
rect 4496 7044 4500 7100
rect 4500 7044 4556 7100
rect 4556 7044 4560 7100
rect 4496 7040 4560 7044
rect 4916 6556 4980 6560
rect 4916 6500 4920 6556
rect 4920 6500 4976 6556
rect 4976 6500 4980 6556
rect 4916 6496 4980 6500
rect 4996 6556 5060 6560
rect 4996 6500 5000 6556
rect 5000 6500 5056 6556
rect 5056 6500 5060 6556
rect 4996 6496 5060 6500
rect 5076 6556 5140 6560
rect 5076 6500 5080 6556
rect 5080 6500 5136 6556
rect 5136 6500 5140 6556
rect 5076 6496 5140 6500
rect 5156 6556 5220 6560
rect 5156 6500 5160 6556
rect 5160 6500 5216 6556
rect 5216 6500 5220 6556
rect 5156 6496 5220 6500
rect 5236 6556 5300 6560
rect 5236 6500 5240 6556
rect 5240 6500 5296 6556
rect 5296 6500 5300 6556
rect 5236 6496 5300 6500
rect 4176 6012 4240 6016
rect 4176 5956 4180 6012
rect 4180 5956 4236 6012
rect 4236 5956 4240 6012
rect 4176 5952 4240 5956
rect 4256 6012 4320 6016
rect 4256 5956 4260 6012
rect 4260 5956 4316 6012
rect 4316 5956 4320 6012
rect 4256 5952 4320 5956
rect 4336 6012 4400 6016
rect 4336 5956 4340 6012
rect 4340 5956 4396 6012
rect 4396 5956 4400 6012
rect 4336 5952 4400 5956
rect 4416 6012 4480 6016
rect 4416 5956 4420 6012
rect 4420 5956 4476 6012
rect 4476 5956 4480 6012
rect 4416 5952 4480 5956
rect 4496 6012 4560 6016
rect 4496 5956 4500 6012
rect 4500 5956 4556 6012
rect 4556 5956 4560 6012
rect 4496 5952 4560 5956
rect 4916 5468 4980 5472
rect 4916 5412 4920 5468
rect 4920 5412 4976 5468
rect 4976 5412 4980 5468
rect 4916 5408 4980 5412
rect 4996 5468 5060 5472
rect 4996 5412 5000 5468
rect 5000 5412 5056 5468
rect 5056 5412 5060 5468
rect 4996 5408 5060 5412
rect 5076 5468 5140 5472
rect 5076 5412 5080 5468
rect 5080 5412 5136 5468
rect 5136 5412 5140 5468
rect 5076 5408 5140 5412
rect 5156 5468 5220 5472
rect 5156 5412 5160 5468
rect 5160 5412 5216 5468
rect 5216 5412 5220 5468
rect 5156 5408 5220 5412
rect 5236 5468 5300 5472
rect 5236 5412 5240 5468
rect 5240 5412 5296 5468
rect 5296 5412 5300 5468
rect 5236 5408 5300 5412
rect 4176 4924 4240 4928
rect 4176 4868 4180 4924
rect 4180 4868 4236 4924
rect 4236 4868 4240 4924
rect 4176 4864 4240 4868
rect 4256 4924 4320 4928
rect 4256 4868 4260 4924
rect 4260 4868 4316 4924
rect 4316 4868 4320 4924
rect 4256 4864 4320 4868
rect 4336 4924 4400 4928
rect 4336 4868 4340 4924
rect 4340 4868 4396 4924
rect 4396 4868 4400 4924
rect 4336 4864 4400 4868
rect 4416 4924 4480 4928
rect 4416 4868 4420 4924
rect 4420 4868 4476 4924
rect 4476 4868 4480 4924
rect 4416 4864 4480 4868
rect 4496 4924 4560 4928
rect 4496 4868 4500 4924
rect 4500 4868 4556 4924
rect 4556 4868 4560 4924
rect 4496 4864 4560 4868
rect 4916 4380 4980 4384
rect 4916 4324 4920 4380
rect 4920 4324 4976 4380
rect 4976 4324 4980 4380
rect 4916 4320 4980 4324
rect 4996 4380 5060 4384
rect 4996 4324 5000 4380
rect 5000 4324 5056 4380
rect 5056 4324 5060 4380
rect 4996 4320 5060 4324
rect 5076 4380 5140 4384
rect 5076 4324 5080 4380
rect 5080 4324 5136 4380
rect 5136 4324 5140 4380
rect 5076 4320 5140 4324
rect 5156 4380 5220 4384
rect 5156 4324 5160 4380
rect 5160 4324 5216 4380
rect 5216 4324 5220 4380
rect 5156 4320 5220 4324
rect 5236 4380 5300 4384
rect 5236 4324 5240 4380
rect 5240 4324 5296 4380
rect 5296 4324 5300 4380
rect 5236 4320 5300 4324
rect 4176 3836 4240 3840
rect 4176 3780 4180 3836
rect 4180 3780 4236 3836
rect 4236 3780 4240 3836
rect 4176 3776 4240 3780
rect 4256 3836 4320 3840
rect 4256 3780 4260 3836
rect 4260 3780 4316 3836
rect 4316 3780 4320 3836
rect 4256 3776 4320 3780
rect 4336 3836 4400 3840
rect 4336 3780 4340 3836
rect 4340 3780 4396 3836
rect 4396 3780 4400 3836
rect 4336 3776 4400 3780
rect 4416 3836 4480 3840
rect 4416 3780 4420 3836
rect 4420 3780 4476 3836
rect 4476 3780 4480 3836
rect 4416 3776 4480 3780
rect 4496 3836 4560 3840
rect 4496 3780 4500 3836
rect 4500 3780 4556 3836
rect 4556 3780 4560 3836
rect 4496 3776 4560 3780
rect 4916 3292 4980 3296
rect 4916 3236 4920 3292
rect 4920 3236 4976 3292
rect 4976 3236 4980 3292
rect 4916 3232 4980 3236
rect 4996 3292 5060 3296
rect 4996 3236 5000 3292
rect 5000 3236 5056 3292
rect 5056 3236 5060 3292
rect 4996 3232 5060 3236
rect 5076 3292 5140 3296
rect 5076 3236 5080 3292
rect 5080 3236 5136 3292
rect 5136 3236 5140 3292
rect 5076 3232 5140 3236
rect 5156 3292 5220 3296
rect 5156 3236 5160 3292
rect 5160 3236 5216 3292
rect 5216 3236 5220 3292
rect 5156 3232 5220 3236
rect 5236 3292 5300 3296
rect 5236 3236 5240 3292
rect 5240 3236 5296 3292
rect 5296 3236 5300 3292
rect 5236 3232 5300 3236
rect 4176 2748 4240 2752
rect 4176 2692 4180 2748
rect 4180 2692 4236 2748
rect 4236 2692 4240 2748
rect 4176 2688 4240 2692
rect 4256 2748 4320 2752
rect 4256 2692 4260 2748
rect 4260 2692 4316 2748
rect 4316 2692 4320 2748
rect 4256 2688 4320 2692
rect 4336 2748 4400 2752
rect 4336 2692 4340 2748
rect 4340 2692 4396 2748
rect 4396 2692 4400 2748
rect 4336 2688 4400 2692
rect 4416 2748 4480 2752
rect 4416 2692 4420 2748
rect 4420 2692 4476 2748
rect 4476 2692 4480 2748
rect 4416 2688 4480 2692
rect 4496 2748 4560 2752
rect 4496 2692 4500 2748
rect 4500 2692 4556 2748
rect 4556 2692 4560 2748
rect 4496 2688 4560 2692
rect 4916 2204 4980 2208
rect 4916 2148 4920 2204
rect 4920 2148 4976 2204
rect 4976 2148 4980 2204
rect 4916 2144 4980 2148
rect 4996 2204 5060 2208
rect 4996 2148 5000 2204
rect 5000 2148 5056 2204
rect 5056 2148 5060 2204
rect 4996 2144 5060 2148
rect 5076 2204 5140 2208
rect 5076 2148 5080 2204
rect 5080 2148 5136 2204
rect 5136 2148 5140 2204
rect 5076 2144 5140 2148
rect 5156 2204 5220 2208
rect 5156 2148 5160 2204
rect 5160 2148 5216 2204
rect 5216 2148 5220 2204
rect 5156 2144 5220 2148
rect 5236 2204 5300 2208
rect 5236 2148 5240 2204
rect 5240 2148 5296 2204
rect 5296 2148 5300 2204
rect 5236 2144 5300 2148
<< metal4 >>
rect 4168 8192 4568 8752
rect 4168 8128 4176 8192
rect 4240 8128 4256 8192
rect 4320 8128 4336 8192
rect 4400 8128 4416 8192
rect 4480 8128 4496 8192
rect 4560 8128 4568 8192
rect 4168 7104 4568 8128
rect 4168 7040 4176 7104
rect 4240 7040 4256 7104
rect 4320 7040 4336 7104
rect 4400 7040 4416 7104
rect 4480 7040 4496 7104
rect 4560 7040 4568 7104
rect 4168 6016 4568 7040
rect 4168 5952 4176 6016
rect 4240 5952 4256 6016
rect 4320 5952 4336 6016
rect 4400 5952 4416 6016
rect 4480 5952 4496 6016
rect 4560 5952 4568 6016
rect 4168 4928 4568 5952
rect 4168 4864 4176 4928
rect 4240 4864 4256 4928
rect 4320 4864 4336 4928
rect 4400 4864 4416 4928
rect 4480 4864 4496 4928
rect 4560 4864 4568 4928
rect 4168 3840 4568 4864
rect 4168 3776 4176 3840
rect 4240 3776 4256 3840
rect 4320 3776 4336 3840
rect 4400 3776 4416 3840
rect 4480 3776 4496 3840
rect 4560 3776 4568 3840
rect 4168 2752 4568 3776
rect 4168 2688 4176 2752
rect 4240 2688 4256 2752
rect 4320 2688 4336 2752
rect 4400 2688 4416 2752
rect 4480 2688 4496 2752
rect 4560 2688 4568 2752
rect 4168 2128 4568 2688
rect 4908 8736 5308 8752
rect 4908 8672 4916 8736
rect 4980 8672 4996 8736
rect 5060 8672 5076 8736
rect 5140 8672 5156 8736
rect 5220 8672 5236 8736
rect 5300 8672 5308 8736
rect 4908 7648 5308 8672
rect 4908 7584 4916 7648
rect 4980 7584 4996 7648
rect 5060 7584 5076 7648
rect 5140 7584 5156 7648
rect 5220 7584 5236 7648
rect 5300 7584 5308 7648
rect 4908 6560 5308 7584
rect 4908 6496 4916 6560
rect 4980 6496 4996 6560
rect 5060 6496 5076 6560
rect 5140 6496 5156 6560
rect 5220 6496 5236 6560
rect 5300 6496 5308 6560
rect 4908 5472 5308 6496
rect 4908 5408 4916 5472
rect 4980 5408 4996 5472
rect 5060 5408 5076 5472
rect 5140 5408 5156 5472
rect 5220 5408 5236 5472
rect 5300 5408 5308 5472
rect 4908 4384 5308 5408
rect 4908 4320 4916 4384
rect 4980 4320 4996 4384
rect 5060 4320 5076 4384
rect 5140 4320 5156 4384
rect 5220 4320 5236 4384
rect 5300 4320 5308 4384
rect 4908 3296 5308 4320
rect 4908 3232 4916 3296
rect 4980 3232 4996 3296
rect 5060 3232 5076 3296
rect 5140 3232 5156 3296
rect 5220 3232 5236 3296
rect 5300 3232 5308 3296
rect 4908 2208 5308 3232
rect 4908 2144 4916 2208
rect 4980 2144 4996 2208
rect 5060 2144 5076 2208
rect 5140 2144 5156 2208
rect 5220 2144 5236 2208
rect 5300 2144 5308 2208
rect 4908 2128 5308 2144
use sky130_fd_sc_hd__and3_1  _14_
timestamp -25199
transform -1 0 4232 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _15_
timestamp -25199
transform 1 0 3772 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _16_
timestamp -25199
transform -1 0 2392 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _17_
timestamp -25199
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _18_
timestamp -25199
transform -1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _19_
timestamp -25199
transform -1 0 2484 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _20_
timestamp -25199
transform 1 0 6348 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _21_
timestamp -25199
transform 1 0 6348 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _22_
timestamp -25199
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _23_
timestamp -25199
transform -1 0 7176 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _24_
timestamp -25199
transform 1 0 6348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _25_
timestamp -25199
transform 1 0 6072 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _26_
timestamp -25199
transform 1 0 6348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _27_
timestamp -25199
transform 1 0 1932 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _28_
timestamp -25199
transform 1 0 4232 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _29_
timestamp -25199
transform 1 0 1656 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _30_
timestamp -25199
transform 1 0 1840 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _31_
timestamp -25199
transform 1 0 1840 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _32_
timestamp -25199
transform -1 0 6256 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _33_
timestamp -25199
transform -1 0 6256 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _34_
timestamp -25199
transform -1 0 6256 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _35_
timestamp -25199
transform -1 0 7176 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _36_
timestamp -25199
transform 1 0 4416 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _37_
timestamp -25199
transform 1 0 5336 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _38_
timestamp -25199
transform 1 0 5244 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _39_
timestamp -25199
transform 1 0 1472 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp -25199
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp -25199
transform -1 0 1840 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp -25199
transform -1 0 1564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp -25199
transform -1 0 1840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -25199
transform 1 0 3864 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp -25199
transform -1 0 4324 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp -25199
transform 1 0 5796 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  fanout13
timestamp -25199
transform -1 0 7544 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout14
timestamp -25199
transform 1 0 2760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout15
timestamp -25199
transform -1 0 4968 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout16
timestamp -25199
transform 1 0 3496 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636943256
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15
timestamp -25199
transform 1 0 2484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21
timestamp -25199
transform 1 0 3036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp -25199
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66
timestamp -25199
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70
timestamp -25199
transform 1 0 7544 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636943256
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636943256
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_27
timestamp -25199
transform 1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_66
timestamp -25199
transform 1 0 7176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_70
timestamp -25199
transform 1 0 7544 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636943256
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636943256
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -25199
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp -25199
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_37
timestamp -25199
transform 1 0 4508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp -25199
transform 1 0 7176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_70
timestamp -25199
transform 1 0 7544 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_5
timestamp 1636943256
transform 1 0 1564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_17
timestamp 1636943256
transform 1 0 2668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_29
timestamp -25199
transform 1 0 3772 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_35
timestamp -25199
transform 1 0 4324 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_66
timestamp -25199
transform 1 0 7176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_70
timestamp -25199
transform 1 0 7544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_6
timestamp -25199
transform 1 0 1656 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_14
timestamp 1636943256
transform 1 0 2392 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp -25199
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_31
timestamp 1636943256
transform 1 0 3956 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_43
timestamp -25199
transform 1 0 5060 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp -25199
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_66
timestamp -25199
transform 1 0 7176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_70
timestamp -25199
transform 1 0 7544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp -25199
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp -25199
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_42
timestamp -25199
transform 1 0 4968 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_66
timestamp -25199
transform 1 0 7176 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_70
timestamp -25199
transform 1 0 7544 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp -25199
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_35
timestamp -25199
transform 1 0 4324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_66
timestamp -25199
transform 1 0 7176 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_70
timestamp -25199
transform 1 0 7544 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_34
timestamp -25199
transform 1 0 4232 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_42
timestamp -25199
transform 1 0 4968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp -25199
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_24
timestamp -25199
transform 1 0 3312 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_32
timestamp -25199
transform 1 0 4048 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp -25199
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_70
timestamp -25199
transform 1 0 7544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp -25199
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_22
timestamp -25199
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636943256
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636943256
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_53
timestamp -25199
transform 1 0 5980 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_63
timestamp -25199
transform 1 0 6900 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_8
timestamp 1636943256
transform 1 0 1840 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_20
timestamp -25199
transform 1 0 2944 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_29
timestamp 1636943256
transform 1 0 3772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_41
timestamp 1636943256
transform 1 0 4876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp -25199
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp -25199
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp -25199
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp -25199
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp -25199
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  output4
timestamp -25199
transform 1 0 6532 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output5
timestamp -25199
transform -1 0 3680 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output6
timestamp -25199
transform -1 0 4416 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output7
timestamp -25199
transform -1 0 4416 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output8
timestamp -25199
transform -1 0 5336 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output9
timestamp -25199
transform -1 0 6256 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output10
timestamp -25199
transform 1 0 7084 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output11
timestamp -25199
transform 1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output12
timestamp -25199
transform 1 0 7084 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -25199
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -25199
transform -1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -25199
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -25199
transform -1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -25199
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -25199
transform -1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -25199
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -25199
transform -1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -25199
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -25199
transform -1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -25199
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -25199
transform -1 0 7912 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -25199
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -25199
transform -1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -25199
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -25199
transform -1 0 7912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -25199
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -25199
transform -1 0 7912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -25199
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -25199
transform -1 0 7912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -25199
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -25199
transform -1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -25199
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -25199
transform -1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -25199
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -25199
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_26
timestamp -25199
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_27
timestamp -25199
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_28
timestamp -25199
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_29
timestamp -25199
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_30
timestamp -25199
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_31
timestamp -25199
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_32
timestamp -25199
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_33
timestamp -25199
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_34
timestamp -25199
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_35
timestamp -25199
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_36
timestamp -25199
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_37
timestamp -25199
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal3 s 8249 9800 9049 9920 0 FreeSans 480 0 0 0 byte_ready_o
port 0 nsew signal output
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 clk
port 1 nsew signal input
flabel metal3 s 8249 1096 9049 1216 0 FreeSans 480 0 0 0 data_parallel_o[0]
port 2 nsew signal output
flabel metal3 s 8249 2184 9049 2304 0 FreeSans 480 0 0 0 data_parallel_o[1]
port 3 nsew signal output
flabel metal3 s 8249 3272 9049 3392 0 FreeSans 480 0 0 0 data_parallel_o[2]
port 4 nsew signal output
flabel metal3 s 8249 4360 9049 4480 0 FreeSans 480 0 0 0 data_parallel_o[3]
port 5 nsew signal output
flabel metal3 s 8249 5448 9049 5568 0 FreeSans 480 0 0 0 data_parallel_o[4]
port 6 nsew signal output
flabel metal3 s 8249 6536 9049 6656 0 FreeSans 480 0 0 0 data_parallel_o[5]
port 7 nsew signal output
flabel metal3 s 8249 7624 9049 7744 0 FreeSans 480 0 0 0 data_parallel_o[6]
port 8 nsew signal output
flabel metal3 s 8249 8712 9049 8832 0 FreeSans 480 0 0 0 data_parallel_o[7]
port 9 nsew signal output
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 data_serial_i
port 10 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 rst_n
port 11 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 valid_serial_i
port 12 nsew signal input
flabel metal4 s 4168 2128 4568 8752 0 FreeSans 1920 90 0 0 vccd1
port 13 nsew power bidirectional
flabel metal4 s 4908 2128 5308 8752 0 FreeSans 1920 90 0 0 vssd1
port 14 nsew ground bidirectional
rlabel via1 4508 8160 4508 8160 0 vccd1
rlabel metal1 4508 8704 4508 8704 0 vssd1
rlabel metal1 4462 6970 4462 6970 0 _00_
rlabel metal1 1886 4794 1886 4794 0 _01_
rlabel metal1 1968 5882 1968 5882 0 _02_
rlabel metal2 1886 6460 1886 6460 0 _03_
rlabel metal1 6026 2482 6026 2482 0 _04_
rlabel metal1 6118 3162 6118 3162 0 _05_
rlabel metal2 5934 3502 5934 3502 0 _06_
rlabel metal2 6854 4284 6854 4284 0 _07_
rlabel metal1 5566 6222 5566 6222 0 _08_
rlabel metal1 5704 5610 5704 5610 0 _09_
rlabel metal1 5835 6970 5835 6970 0 _10_
rlabel metal2 1794 7582 1794 7582 0 _11_
rlabel metal1 3864 5814 3864 5814 0 _12_
rlabel metal1 1794 6222 1794 6222 0 _13_
rlabel metal2 6854 9197 6854 9197 0 byte_ready_o
rlabel metal2 3818 2941 3818 2941 0 clk
rlabel metal1 5014 5338 5014 5338 0 clknet_0_clk
rlabel metal1 3588 6290 3588 6290 0 clknet_1_0__leaf_clk
rlabel metal1 5290 6732 5290 6732 0 clknet_1_1__leaf_clk
rlabel metal2 3450 4794 3450 4794 0 count\[0\]
rlabel metal1 3818 5882 3818 5882 0 count\[1\]
rlabel metal1 2944 6630 2944 6630 0 count\[2\]
rlabel metal1 6026 2312 6026 2312 0 data_parallel_o[0]
rlabel metal1 6118 2924 6118 2924 0 data_parallel_o[1]
rlabel metal1 4508 2482 4508 2482 0 data_parallel_o[2]
rlabel metal1 5290 3570 5290 3570 0 data_parallel_o[3]
rlabel metal2 5934 5389 5934 5389 0 data_parallel_o[4]
rlabel metal2 7406 6647 7406 6647 0 data_parallel_o[5]
rlabel metal2 7406 7735 7406 7735 0 data_parallel_o[6]
rlabel metal2 7406 8653 7406 8653 0 data_parallel_o[7]
rlabel metal1 1380 6766 1380 6766 0 data_serial_i
rlabel metal2 1610 7378 1610 7378 0 net1
rlabel metal2 6854 6596 6854 6596 0 net10
rlabel metal2 6946 7174 6946 7174 0 net11
rlabel metal1 6762 7514 6762 7514 0 net12
rlabel metal2 6578 5678 6578 5678 0 net13
rlabel via1 3994 5610 3994 5610 0 net14
rlabel metal1 6033 6358 6033 6358 0 net15
rlabel metal1 3726 5304 3726 5304 0 net16
rlabel metal2 3634 6018 3634 6018 0 net2
rlabel metal2 2898 8092 2898 8092 0 net3
rlabel metal1 6302 7310 6302 7310 0 net4
rlabel metal2 4462 2312 4462 2312 0 net5
rlabel metal1 4508 3026 4508 3026 0 net6
rlabel metal1 6762 3162 6762 3162 0 net7
rlabel metal1 6808 4250 6808 4250 0 net8
rlabel metal1 6486 6426 6486 6426 0 net9
rlabel via2 1426 4165 1426 4165 0 rst_n
rlabel metal1 1380 8466 1380 8466 0 valid_serial_i
<< properties >>
string FIXED_BBOX 0 0 9049 11193
<< end >>
