VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pmu
  CLASS BLOCK ;
  FOREIGN pmu ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 150.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END clk
  PIN pm_current_s0_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 10.920 150.000 11.520 ;
    END
  END pm_current_s0_o[0]
  PIN pm_current_s0_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 15.000 150.000 15.600 ;
    END
  END pm_current_s0_o[1]
  PIN pm_current_s0_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 19.080 150.000 19.680 ;
    END
  END pm_current_s0_o[2]
  PIN pm_current_s0_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 23.160 150.000 23.760 ;
    END
  END pm_current_s0_o[3]
  PIN pm_current_s0_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 27.240 150.000 27.840 ;
    END
  END pm_current_s0_o[4]
  PIN pm_current_s0_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 31.320 150.000 31.920 ;
    END
  END pm_current_s0_o[5]
  PIN pm_current_s0_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 35.400 150.000 36.000 ;
    END
  END pm_current_s0_o[6]
  PIN pm_current_s0_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 39.480 150.000 40.080 ;
    END
  END pm_current_s0_o[7]
  PIN pm_current_s1_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 43.560 150.000 44.160 ;
    END
  END pm_current_s1_o[0]
  PIN pm_current_s1_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 47.640 150.000 48.240 ;
    END
  END pm_current_s1_o[1]
  PIN pm_current_s1_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 51.720 150.000 52.320 ;
    END
  END pm_current_s1_o[2]
  PIN pm_current_s1_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 55.800 150.000 56.400 ;
    END
  END pm_current_s1_o[3]
  PIN pm_current_s1_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 59.880 150.000 60.480 ;
    END
  END pm_current_s1_o[4]
  PIN pm_current_s1_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 63.960 150.000 64.560 ;
    END
  END pm_current_s1_o[5]
  PIN pm_current_s1_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 68.040 150.000 68.640 ;
    END
  END pm_current_s1_o[6]
  PIN pm_current_s1_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 72.120 150.000 72.720 ;
    END
  END pm_current_s1_o[7]
  PIN pm_current_s2_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 76.200 150.000 76.800 ;
    END
  END pm_current_s2_o[0]
  PIN pm_current_s2_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 80.280 150.000 80.880 ;
    END
  END pm_current_s2_o[1]
  PIN pm_current_s2_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 84.360 150.000 84.960 ;
    END
  END pm_current_s2_o[2]
  PIN pm_current_s2_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 88.440 150.000 89.040 ;
    END
  END pm_current_s2_o[3]
  PIN pm_current_s2_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 92.520 150.000 93.120 ;
    END
  END pm_current_s2_o[4]
  PIN pm_current_s2_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 96.600 150.000 97.200 ;
    END
  END pm_current_s2_o[5]
  PIN pm_current_s2_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 100.680 150.000 101.280 ;
    END
  END pm_current_s2_o[6]
  PIN pm_current_s2_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 104.760 150.000 105.360 ;
    END
  END pm_current_s2_o[7]
  PIN pm_current_s3_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 108.840 150.000 109.440 ;
    END
  END pm_current_s3_o[0]
  PIN pm_current_s3_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 112.920 150.000 113.520 ;
    END
  END pm_current_s3_o[1]
  PIN pm_current_s3_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 117.000 150.000 117.600 ;
    END
  END pm_current_s3_o[2]
  PIN pm_current_s3_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 121.080 150.000 121.680 ;
    END
  END pm_current_s3_o[3]
  PIN pm_current_s3_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 125.160 150.000 125.760 ;
    END
  END pm_current_s3_o[4]
  PIN pm_current_s3_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 129.240 150.000 129.840 ;
    END
  END pm_current_s3_o[5]
  PIN pm_current_s3_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 133.320 150.000 133.920 ;
    END
  END pm_current_s3_o[6]
  PIN pm_current_s3_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 137.400 150.000 138.000 ;
    END
  END pm_current_s3_o[7]
  PIN pm_new_s0_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END pm_new_s0_i[0]
  PIN pm_new_s0_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END pm_new_s0_i[1]
  PIN pm_new_s0_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END pm_new_s0_i[2]
  PIN pm_new_s0_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END pm_new_s0_i[3]
  PIN pm_new_s0_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END pm_new_s0_i[4]
  PIN pm_new_s0_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END pm_new_s0_i[5]
  PIN pm_new_s0_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END pm_new_s0_i[6]
  PIN pm_new_s0_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END pm_new_s0_i[7]
  PIN pm_new_s1_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END pm_new_s1_i[0]
  PIN pm_new_s1_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END pm_new_s1_i[1]
  PIN pm_new_s1_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END pm_new_s1_i[2]
  PIN pm_new_s1_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END pm_new_s1_i[3]
  PIN pm_new_s1_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END pm_new_s1_i[4]
  PIN pm_new_s1_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END pm_new_s1_i[5]
  PIN pm_new_s1_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END pm_new_s1_i[6]
  PIN pm_new_s1_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END pm_new_s1_i[7]
  PIN pm_new_s2_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END pm_new_s2_i[0]
  PIN pm_new_s2_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END pm_new_s2_i[1]
  PIN pm_new_s2_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END pm_new_s2_i[2]
  PIN pm_new_s2_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END pm_new_s2_i[3]
  PIN pm_new_s2_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END pm_new_s2_i[4]
  PIN pm_new_s2_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END pm_new_s2_i[5]
  PIN pm_new_s2_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END pm_new_s2_i[6]
  PIN pm_new_s2_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END pm_new_s2_i[7]
  PIN pm_new_s3_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END pm_new_s3_i[0]
  PIN pm_new_s3_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END pm_new_s3_i[1]
  PIN pm_new_s3_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END pm_new_s3_i[2]
  PIN pm_new_s3_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END pm_new_s3_i[3]
  PIN pm_new_s3_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END pm_new_s3_i[4]
  PIN pm_new_s3_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END pm_new_s3_i[5]
  PIN pm_new_s3_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END pm_new_s3_i[6]
  PIN pm_new_s3_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END pm_new_s3_i[7]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END rst_n
  PIN valid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END valid_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.520 10.640 16.520 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.520 10.640 56.520 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.520 10.640 96.520 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.520 10.640 136.520 138.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 18.220 10.640 20.220 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.220 10.640 60.220 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.220 10.640 100.220 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.220 10.640 140.220 138.960 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 144.630 138.910 ;
      LAYER li1 ;
        RECT 5.520 10.795 144.440 138.805 ;
      LAYER met1 ;
        RECT 0.530 10.640 144.440 138.960 ;
      LAYER met2 ;
        RECT 0.550 5.595 142.050 143.325 ;
      LAYER met3 ;
        RECT 4.400 142.440 146.000 143.305 ;
        RECT 0.525 139.760 146.000 142.440 ;
        RECT 4.400 138.400 146.000 139.760 ;
        RECT 4.400 138.360 145.600 138.400 ;
        RECT 0.525 137.000 145.600 138.360 ;
        RECT 0.525 135.680 146.000 137.000 ;
        RECT 4.400 134.320 146.000 135.680 ;
        RECT 4.400 134.280 145.600 134.320 ;
        RECT 0.525 132.920 145.600 134.280 ;
        RECT 0.525 131.600 146.000 132.920 ;
        RECT 4.400 130.240 146.000 131.600 ;
        RECT 4.400 130.200 145.600 130.240 ;
        RECT 0.525 128.840 145.600 130.200 ;
        RECT 0.525 127.520 146.000 128.840 ;
        RECT 4.400 126.160 146.000 127.520 ;
        RECT 4.400 126.120 145.600 126.160 ;
        RECT 0.525 124.760 145.600 126.120 ;
        RECT 0.525 123.440 146.000 124.760 ;
        RECT 4.400 122.080 146.000 123.440 ;
        RECT 4.400 122.040 145.600 122.080 ;
        RECT 0.525 120.680 145.600 122.040 ;
        RECT 0.525 119.360 146.000 120.680 ;
        RECT 4.400 118.000 146.000 119.360 ;
        RECT 4.400 117.960 145.600 118.000 ;
        RECT 0.525 116.600 145.600 117.960 ;
        RECT 0.525 115.280 146.000 116.600 ;
        RECT 4.400 113.920 146.000 115.280 ;
        RECT 4.400 113.880 145.600 113.920 ;
        RECT 0.525 112.520 145.600 113.880 ;
        RECT 0.525 111.200 146.000 112.520 ;
        RECT 4.400 109.840 146.000 111.200 ;
        RECT 4.400 109.800 145.600 109.840 ;
        RECT 0.525 108.440 145.600 109.800 ;
        RECT 0.525 107.120 146.000 108.440 ;
        RECT 4.400 105.760 146.000 107.120 ;
        RECT 4.400 105.720 145.600 105.760 ;
        RECT 0.525 104.360 145.600 105.720 ;
        RECT 0.525 103.040 146.000 104.360 ;
        RECT 4.400 101.680 146.000 103.040 ;
        RECT 4.400 101.640 145.600 101.680 ;
        RECT 0.525 100.280 145.600 101.640 ;
        RECT 0.525 98.960 146.000 100.280 ;
        RECT 4.400 97.600 146.000 98.960 ;
        RECT 4.400 97.560 145.600 97.600 ;
        RECT 0.525 96.200 145.600 97.560 ;
        RECT 0.525 94.880 146.000 96.200 ;
        RECT 4.400 93.520 146.000 94.880 ;
        RECT 4.400 93.480 145.600 93.520 ;
        RECT 0.525 92.120 145.600 93.480 ;
        RECT 0.525 90.800 146.000 92.120 ;
        RECT 4.400 89.440 146.000 90.800 ;
        RECT 4.400 89.400 145.600 89.440 ;
        RECT 0.525 88.040 145.600 89.400 ;
        RECT 0.525 86.720 146.000 88.040 ;
        RECT 4.400 85.360 146.000 86.720 ;
        RECT 4.400 85.320 145.600 85.360 ;
        RECT 0.525 83.960 145.600 85.320 ;
        RECT 0.525 82.640 146.000 83.960 ;
        RECT 4.400 81.280 146.000 82.640 ;
        RECT 4.400 81.240 145.600 81.280 ;
        RECT 0.525 79.880 145.600 81.240 ;
        RECT 0.525 78.560 146.000 79.880 ;
        RECT 4.400 77.200 146.000 78.560 ;
        RECT 4.400 77.160 145.600 77.200 ;
        RECT 0.525 75.800 145.600 77.160 ;
        RECT 0.525 74.480 146.000 75.800 ;
        RECT 4.400 73.120 146.000 74.480 ;
        RECT 4.400 73.080 145.600 73.120 ;
        RECT 0.525 71.720 145.600 73.080 ;
        RECT 0.525 70.400 146.000 71.720 ;
        RECT 4.400 69.040 146.000 70.400 ;
        RECT 4.400 69.000 145.600 69.040 ;
        RECT 0.525 67.640 145.600 69.000 ;
        RECT 0.525 66.320 146.000 67.640 ;
        RECT 4.400 64.960 146.000 66.320 ;
        RECT 4.400 64.920 145.600 64.960 ;
        RECT 0.525 63.560 145.600 64.920 ;
        RECT 0.525 62.240 146.000 63.560 ;
        RECT 4.400 60.880 146.000 62.240 ;
        RECT 4.400 60.840 145.600 60.880 ;
        RECT 0.525 59.480 145.600 60.840 ;
        RECT 0.525 58.160 146.000 59.480 ;
        RECT 4.400 56.800 146.000 58.160 ;
        RECT 4.400 56.760 145.600 56.800 ;
        RECT 0.525 55.400 145.600 56.760 ;
        RECT 0.525 54.080 146.000 55.400 ;
        RECT 4.400 52.720 146.000 54.080 ;
        RECT 4.400 52.680 145.600 52.720 ;
        RECT 0.525 51.320 145.600 52.680 ;
        RECT 0.525 50.000 146.000 51.320 ;
        RECT 4.400 48.640 146.000 50.000 ;
        RECT 4.400 48.600 145.600 48.640 ;
        RECT 0.525 47.240 145.600 48.600 ;
        RECT 0.525 45.920 146.000 47.240 ;
        RECT 4.400 44.560 146.000 45.920 ;
        RECT 4.400 44.520 145.600 44.560 ;
        RECT 0.525 43.160 145.600 44.520 ;
        RECT 0.525 41.840 146.000 43.160 ;
        RECT 4.400 40.480 146.000 41.840 ;
        RECT 4.400 40.440 145.600 40.480 ;
        RECT 0.525 39.080 145.600 40.440 ;
        RECT 0.525 37.760 146.000 39.080 ;
        RECT 4.400 36.400 146.000 37.760 ;
        RECT 4.400 36.360 145.600 36.400 ;
        RECT 0.525 35.000 145.600 36.360 ;
        RECT 0.525 33.680 146.000 35.000 ;
        RECT 4.400 32.320 146.000 33.680 ;
        RECT 4.400 32.280 145.600 32.320 ;
        RECT 0.525 30.920 145.600 32.280 ;
        RECT 0.525 29.600 146.000 30.920 ;
        RECT 4.400 28.240 146.000 29.600 ;
        RECT 4.400 28.200 145.600 28.240 ;
        RECT 0.525 26.840 145.600 28.200 ;
        RECT 0.525 25.520 146.000 26.840 ;
        RECT 4.400 24.160 146.000 25.520 ;
        RECT 4.400 24.120 145.600 24.160 ;
        RECT 0.525 22.760 145.600 24.120 ;
        RECT 0.525 21.440 146.000 22.760 ;
        RECT 4.400 20.080 146.000 21.440 ;
        RECT 4.400 20.040 145.600 20.080 ;
        RECT 0.525 18.680 145.600 20.040 ;
        RECT 0.525 17.360 146.000 18.680 ;
        RECT 4.400 16.000 146.000 17.360 ;
        RECT 4.400 15.960 145.600 16.000 ;
        RECT 0.525 14.600 145.600 15.960 ;
        RECT 0.525 13.280 146.000 14.600 ;
        RECT 4.400 11.920 146.000 13.280 ;
        RECT 4.400 11.880 145.600 11.920 ;
        RECT 0.525 10.520 145.600 11.880 ;
        RECT 0.525 9.200 146.000 10.520 ;
        RECT 4.400 7.800 146.000 9.200 ;
        RECT 0.525 5.120 146.000 7.800 ;
        RECT 4.400 4.270 146.000 5.120 ;
      LAYER met4 ;
        RECT 3.975 24.655 14.120 77.345 ;
        RECT 16.920 24.655 17.820 77.345 ;
        RECT 20.620 24.655 54.120 77.345 ;
        RECT 56.920 24.655 57.665 77.345 ;
  END
END pmu
END LIBRARY

