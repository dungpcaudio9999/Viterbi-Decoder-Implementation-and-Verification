magic
tech sky130A
magscale 1 2
timestamp 1769196404
<< viali >>
rect 2145 27557 2179 27591
rect 28365 27489 28399 27523
rect 1409 27421 1443 27455
rect 1685 27421 1719 27455
rect 1961 27421 1995 27455
rect 11713 27421 11747 27455
rect 28089 27421 28123 27455
rect 1593 27285 1627 27319
rect 1869 27285 1903 27319
rect 11529 27285 11563 27319
rect 11069 27081 11103 27115
rect 11989 27081 12023 27115
rect 10977 26945 11011 26979
rect 11897 26945 11931 26979
rect 12541 26945 12575 26979
rect 28089 26945 28123 26979
rect 11253 26877 11287 26911
rect 12173 26877 12207 26911
rect 28365 26877 28399 26911
rect 10609 26741 10643 26775
rect 11529 26741 11563 26775
rect 12357 26741 12391 26775
rect 9183 26537 9217 26571
rect 1593 26469 1627 26503
rect 10609 26401 10643 26435
rect 11437 26401 11471 26435
rect 13553 26401 13587 26435
rect 1409 26333 1443 26367
rect 10977 26333 11011 26367
rect 11069 26333 11103 26367
rect 12863 26333 12897 26367
rect 28089 26333 28123 26367
rect 13369 26265 13403 26299
rect 28365 26265 28399 26299
rect 13001 26197 13035 26231
rect 13461 26197 13495 26231
rect 10885 25993 10919 26027
rect 13507 25993 13541 26027
rect 1409 25857 1443 25891
rect 10977 25857 11011 25891
rect 10793 25789 10827 25823
rect 11713 25789 11747 25823
rect 12081 25789 12115 25823
rect 1593 25653 1627 25687
rect 11345 25653 11379 25687
rect 11437 25313 11471 25347
rect 11069 25245 11103 25279
rect 12863 25245 12897 25279
rect 28089 25245 28123 25279
rect 28365 25177 28399 25211
rect 1409 24769 1443 24803
rect 13875 24769 13909 24803
rect 28089 24769 28123 24803
rect 12081 24701 12115 24735
rect 12449 24701 12483 24735
rect 28365 24701 28399 24735
rect 1593 24565 1627 24599
rect 13001 24361 13035 24395
rect 13461 24225 13495 24259
rect 13553 24225 13587 24259
rect 1409 24157 1443 24191
rect 11069 24157 11103 24191
rect 11437 24157 11471 24191
rect 13369 24157 13403 24191
rect 12863 24089 12897 24123
rect 1593 24021 1627 24055
rect 11529 23817 11563 23851
rect 11897 23817 11931 23851
rect 11989 23749 12023 23783
rect 28089 23681 28123 23715
rect 12081 23613 12115 23647
rect 28365 23613 28399 23647
rect 11437 23205 11471 23239
rect 14565 23137 14599 23171
rect 14657 23137 14691 23171
rect 1409 23069 1443 23103
rect 11253 23069 11287 23103
rect 14473 23069 14507 23103
rect 28089 23069 28123 23103
rect 11529 23001 11563 23035
rect 28365 23001 28399 23035
rect 1593 22933 1627 22967
rect 13001 22933 13035 22967
rect 14105 22933 14139 22967
rect 11989 22729 12023 22763
rect 14887 22729 14921 22763
rect 11897 22661 11931 22695
rect 1409 22593 1443 22627
rect 12449 22593 12483 22627
rect 13461 22593 13495 22627
rect 12081 22525 12115 22559
rect 13093 22525 13127 22559
rect 12633 22457 12667 22491
rect 1593 22389 1627 22423
rect 11529 22389 11563 22423
rect 11069 22049 11103 22083
rect 14565 22049 14599 22083
rect 14749 22049 14783 22083
rect 11437 21981 11471 22015
rect 28089 21981 28123 22015
rect 12863 21913 12897 21947
rect 14473 21913 14507 21947
rect 28365 21913 28399 21947
rect 14105 21845 14139 21879
rect 14887 21641 14921 21675
rect 1409 21505 1443 21539
rect 13093 21505 13127 21539
rect 13461 21505 13495 21539
rect 28089 21505 28123 21539
rect 28365 21437 28399 21471
rect 1593 21301 1627 21335
rect 14565 20961 14599 20995
rect 14657 20961 14691 20995
rect 1409 20893 1443 20927
rect 14473 20825 14507 20859
rect 1593 20757 1627 20791
rect 14105 20757 14139 20791
rect 14887 20417 14921 20451
rect 28089 20417 28123 20451
rect 13093 20349 13127 20383
rect 13461 20349 13495 20383
rect 28365 20349 28399 20383
rect 1593 20009 1627 20043
rect 11069 19873 11103 19907
rect 13645 19873 13679 19907
rect 13829 19873 13863 19907
rect 1409 19805 1443 19839
rect 11437 19805 11471 19839
rect 12863 19805 12897 19839
rect 28089 19805 28123 19839
rect 28365 19737 28399 19771
rect 13185 19669 13219 19703
rect 13553 19669 13587 19703
rect 1593 19465 1627 19499
rect 11529 19465 11563 19499
rect 11897 19465 11931 19499
rect 11989 19397 12023 19431
rect 1409 19329 1443 19363
rect 12633 19329 12667 19363
rect 13001 19329 13035 19363
rect 14427 19329 14461 19363
rect 12081 19261 12115 19295
rect 14657 18785 14691 18819
rect 14565 18717 14599 18751
rect 28089 18717 28123 18751
rect 12265 18649 12299 18683
rect 28365 18649 28399 18683
rect 14105 18581 14139 18615
rect 14473 18581 14507 18615
rect 1593 18377 1627 18411
rect 1409 18241 1443 18275
rect 12725 18241 12759 18275
rect 14151 18241 14185 18275
rect 28089 18241 28123 18275
rect 12357 18173 12391 18207
rect 28365 18173 28399 18207
rect 13461 17833 13495 17867
rect 14565 17697 14599 17731
rect 14657 17697 14691 17731
rect 1409 17629 1443 17663
rect 12173 17629 12207 17663
rect 1593 17493 1627 17527
rect 14105 17493 14139 17527
rect 14473 17493 14507 17527
rect 12449 17153 12483 17187
rect 13875 17153 13909 17187
rect 28089 17153 28123 17187
rect 12081 17085 12115 17119
rect 28365 17085 28399 17119
rect 1409 16541 1443 16575
rect 11621 16541 11655 16575
rect 11989 16541 12023 16575
rect 28089 16541 28123 16575
rect 28365 16473 28399 16507
rect 1593 16405 1627 16439
rect 13415 16405 13449 16439
rect 10885 16201 10919 16235
rect 1409 16065 1443 16099
rect 10977 16065 11011 16099
rect 11529 16065 11563 16099
rect 10701 15997 10735 16031
rect 11897 15997 11931 16031
rect 11345 15929 11379 15963
rect 1593 15861 1627 15895
rect 13323 15861 13357 15895
rect 11713 15657 11747 15691
rect 12081 15657 12115 15691
rect 10793 15589 10827 15623
rect 12541 15521 12575 15555
rect 12725 15521 12759 15555
rect 10977 15453 11011 15487
rect 28089 15453 28123 15487
rect 11253 15385 11287 15419
rect 11621 15385 11655 15419
rect 12449 15385 12483 15419
rect 28365 15385 28399 15419
rect 11345 15317 11379 15351
rect 11069 15113 11103 15147
rect 11529 15045 11563 15079
rect 1409 14977 1443 15011
rect 10977 14977 11011 15011
rect 28089 14977 28123 15011
rect 11161 14909 11195 14943
rect 28365 14909 28399 14943
rect 1593 14841 1627 14875
rect 10609 14773 10643 14807
rect 12817 14773 12851 14807
rect 10977 14433 11011 14467
rect 1409 14365 1443 14399
rect 10609 14365 10643 14399
rect 12403 14365 12437 14399
rect 12541 14297 12575 14331
rect 12725 14297 12759 14331
rect 1593 14229 1627 14263
rect 11989 14025 12023 14059
rect 11897 13889 11931 13923
rect 28089 13889 28123 13923
rect 12081 13821 12115 13855
rect 28365 13821 28399 13855
rect 11529 13685 11563 13719
rect 12403 13481 12437 13515
rect 10977 13345 11011 13379
rect 13001 13345 13035 13379
rect 13093 13345 13127 13379
rect 1409 13277 1443 13311
rect 10609 13277 10643 13311
rect 12909 13277 12943 13311
rect 28089 13277 28123 13311
rect 28365 13209 28399 13243
rect 1593 13141 1627 13175
rect 12541 13141 12575 13175
rect 10885 12937 10919 12971
rect 13323 12937 13357 12971
rect 1409 12801 1443 12835
rect 10977 12801 11011 12835
rect 10793 12733 10827 12767
rect 11529 12733 11563 12767
rect 11897 12733 11931 12767
rect 1593 12597 1627 12631
rect 11345 12597 11379 12631
rect 11069 12257 11103 12291
rect 10517 12189 10551 12223
rect 10701 12189 10735 12223
rect 12495 12189 12529 12223
rect 28089 12189 28123 12223
rect 28365 12121 28399 12155
rect 1409 11713 1443 11747
rect 11345 11713 11379 11747
rect 13323 11713 13357 11747
rect 28089 11713 28123 11747
rect 11529 11645 11563 11679
rect 11897 11645 11931 11679
rect 28365 11645 28399 11679
rect 10057 11577 10091 11611
rect 1593 11509 1627 11543
rect 1593 11237 1627 11271
rect 1409 11101 1443 11135
rect 10701 11101 10735 11135
rect 11069 11101 11103 11135
rect 12495 11033 12529 11067
rect 10885 10761 10919 10795
rect 11529 10761 11563 10795
rect 11989 10761 12023 10795
rect 10333 10693 10367 10727
rect 10977 10693 11011 10727
rect 11897 10625 11931 10659
rect 28089 10625 28123 10659
rect 10517 10557 10551 10591
rect 10793 10557 10827 10591
rect 12081 10557 12115 10591
rect 28365 10557 28399 10591
rect 11345 10489 11379 10523
rect 12633 10149 12667 10183
rect 11069 10081 11103 10115
rect 13185 10081 13219 10115
rect 1409 10013 1443 10047
rect 10701 10013 10735 10047
rect 12495 10013 12529 10047
rect 13001 10013 13035 10047
rect 28089 10013 28123 10047
rect 28365 9945 28399 9979
rect 1593 9877 1627 9911
rect 13093 9877 13127 9911
rect 10885 9673 10919 9707
rect 1409 9537 1443 9571
rect 10977 9537 11011 9571
rect 11529 9537 11563 9571
rect 10793 9469 10827 9503
rect 11897 9469 11931 9503
rect 11345 9401 11379 9435
rect 1593 9333 1627 9367
rect 13323 9333 13357 9367
rect 11897 9129 11931 9163
rect 11989 8925 12023 8959
rect 28089 8925 28123 8959
rect 28365 8857 28399 8891
rect 10885 8585 10919 8619
rect 10977 8517 11011 8551
rect 1409 8449 1443 8483
rect 28089 8449 28123 8483
rect 10793 8381 10827 8415
rect 11529 8381 11563 8415
rect 11805 8381 11839 8415
rect 13277 8381 13311 8415
rect 28365 8381 28399 8415
rect 1593 8313 1627 8347
rect 11345 8245 11379 8279
rect 10701 7905 10735 7939
rect 1409 7837 1443 7871
rect 10977 7769 11011 7803
rect 1593 7701 1627 7735
rect 12449 7701 12483 7735
rect 11529 7497 11563 7531
rect 11897 7497 11931 7531
rect 11989 7429 12023 7463
rect 28089 7361 28123 7395
rect 12081 7293 12115 7327
rect 28365 7293 28399 7327
rect 11069 6817 11103 6851
rect 1409 6749 1443 6783
rect 10885 6749 10919 6783
rect 12817 6749 12851 6783
rect 28089 6749 28123 6783
rect 28365 6681 28399 6715
rect 1593 6613 1627 6647
rect 10057 6409 10091 6443
rect 10885 6409 10919 6443
rect 1409 6273 1443 6307
rect 10149 6273 10183 6307
rect 10977 6273 11011 6307
rect 11529 6273 11563 6307
rect 9965 6205 9999 6239
rect 10701 6205 10735 6239
rect 11805 6205 11839 6239
rect 11345 6137 11379 6171
rect 1593 6069 1627 6103
rect 10517 6069 10551 6103
rect 13277 6069 13311 6103
rect 10701 5729 10735 5763
rect 10977 5729 11011 5763
rect 12449 5729 12483 5763
rect 28089 5661 28123 5695
rect 28365 5593 28399 5627
rect 11989 5321 12023 5355
rect 1409 5185 1443 5219
rect 11897 5185 11931 5219
rect 28089 5185 28123 5219
rect 12081 5117 12115 5151
rect 28365 5117 28399 5151
rect 1593 4981 1627 5015
rect 11529 4981 11563 5015
rect 10609 4641 10643 4675
rect 10885 4641 10919 4675
rect 12909 4641 12943 4675
rect 13001 4641 13035 4675
rect 1409 4573 1443 4607
rect 1593 4437 1627 4471
rect 12357 4437 12391 4471
rect 12449 4437 12483 4471
rect 12817 4437 12851 4471
rect 11161 4165 11195 4199
rect 11345 4097 11379 4131
rect 28089 4097 28123 4131
rect 11529 4029 11563 4063
rect 11805 4029 11839 4063
rect 13277 4029 13311 4063
rect 28365 4029 28399 4063
rect 10333 3689 10367 3723
rect 12449 3689 12483 3723
rect 10609 3553 10643 3587
rect 10885 3553 10919 3587
rect 12357 3553 12391 3587
rect 12909 3553 12943 3587
rect 13001 3553 13035 3587
rect 1409 3485 1443 3519
rect 12817 3485 12851 3519
rect 28089 3485 28123 3519
rect 10425 3417 10459 3451
rect 13277 3417 13311 3451
rect 13461 3417 13495 3451
rect 28365 3417 28399 3451
rect 1593 3349 1627 3383
rect 10885 3145 10919 3179
rect 1409 3009 1443 3043
rect 10977 3009 11011 3043
rect 11529 3009 11563 3043
rect 10701 2941 10735 2975
rect 11805 2941 11839 2975
rect 11345 2873 11379 2907
rect 1593 2805 1627 2839
rect 13277 2805 13311 2839
rect 11897 2601 11931 2635
rect 1409 2397 1443 2431
rect 11989 2397 12023 2431
rect 28089 2397 28123 2431
rect 28365 2329 28399 2363
rect 1593 2261 1627 2295
<< metal1 >>
rect 1104 27770 28888 27792
rect 1104 27718 2918 27770
rect 2970 27718 2982 27770
rect 3034 27718 3046 27770
rect 3098 27718 3110 27770
rect 3162 27718 3174 27770
rect 3226 27718 3238 27770
rect 3290 27718 10918 27770
rect 10970 27718 10982 27770
rect 11034 27718 11046 27770
rect 11098 27718 11110 27770
rect 11162 27718 11174 27770
rect 11226 27718 11238 27770
rect 11290 27718 18918 27770
rect 18970 27718 18982 27770
rect 19034 27718 19046 27770
rect 19098 27718 19110 27770
rect 19162 27718 19174 27770
rect 19226 27718 19238 27770
rect 19290 27718 26918 27770
rect 26970 27718 26982 27770
rect 27034 27718 27046 27770
rect 27098 27718 27110 27770
rect 27162 27718 27174 27770
rect 27226 27718 27238 27770
rect 27290 27718 28888 27770
rect 1104 27696 28888 27718
rect 1026 27548 1032 27600
rect 1084 27588 1090 27600
rect 2133 27591 2191 27597
rect 1084 27560 1992 27588
rect 1084 27548 1090 27560
rect 934 27480 940 27532
rect 992 27520 998 27532
rect 992 27492 1716 27520
rect 992 27480 998 27492
rect 842 27412 848 27464
rect 900 27452 906 27464
rect 1688 27461 1716 27492
rect 1964 27461 1992 27560
rect 2133 27557 2145 27591
rect 2179 27588 2191 27591
rect 10962 27588 10968 27600
rect 2179 27560 10968 27588
rect 2179 27557 2191 27560
rect 2133 27551 2191 27557
rect 10962 27548 10968 27560
rect 11020 27548 11026 27600
rect 28350 27480 28356 27532
rect 28408 27480 28414 27532
rect 1397 27455 1455 27461
rect 1397 27452 1409 27455
rect 900 27424 1409 27452
rect 900 27412 906 27424
rect 1397 27421 1409 27424
rect 1443 27421 1455 27455
rect 1397 27415 1455 27421
rect 1673 27455 1731 27461
rect 1673 27421 1685 27455
rect 1719 27421 1731 27455
rect 1673 27415 1731 27421
rect 1949 27455 2007 27461
rect 1949 27421 1961 27455
rect 1995 27421 2007 27455
rect 1949 27415 2007 27421
rect 11701 27455 11759 27461
rect 11701 27421 11713 27455
rect 11747 27452 11759 27455
rect 12342 27452 12348 27464
rect 11747 27424 12348 27452
rect 11747 27421 11759 27424
rect 11701 27415 11759 27421
rect 12342 27412 12348 27424
rect 12400 27412 12406 27464
rect 21266 27412 21272 27464
rect 21324 27452 21330 27464
rect 28077 27455 28135 27461
rect 28077 27452 28089 27455
rect 21324 27424 28089 27452
rect 21324 27412 21330 27424
rect 28077 27421 28089 27424
rect 28123 27421 28135 27455
rect 28077 27415 28135 27421
rect 11422 27384 11428 27396
rect 1872 27356 11428 27384
rect 1578 27276 1584 27328
rect 1636 27276 1642 27328
rect 1872 27325 1900 27356
rect 11422 27344 11428 27356
rect 11480 27344 11486 27396
rect 1857 27319 1915 27325
rect 1857 27285 1869 27319
rect 1903 27285 1915 27319
rect 1857 27279 1915 27285
rect 11517 27319 11575 27325
rect 11517 27285 11529 27319
rect 11563 27316 11575 27319
rect 12158 27316 12164 27328
rect 11563 27288 12164 27316
rect 11563 27285 11575 27288
rect 11517 27279 11575 27285
rect 12158 27276 12164 27288
rect 12216 27276 12222 27328
rect 1104 27226 28888 27248
rect 1104 27174 3658 27226
rect 3710 27174 3722 27226
rect 3774 27174 3786 27226
rect 3838 27174 3850 27226
rect 3902 27174 3914 27226
rect 3966 27174 3978 27226
rect 4030 27174 11658 27226
rect 11710 27174 11722 27226
rect 11774 27174 11786 27226
rect 11838 27174 11850 27226
rect 11902 27174 11914 27226
rect 11966 27174 11978 27226
rect 12030 27174 19658 27226
rect 19710 27174 19722 27226
rect 19774 27174 19786 27226
rect 19838 27174 19850 27226
rect 19902 27174 19914 27226
rect 19966 27174 19978 27226
rect 20030 27174 27658 27226
rect 27710 27174 27722 27226
rect 27774 27174 27786 27226
rect 27838 27174 27850 27226
rect 27902 27174 27914 27226
rect 27966 27174 27978 27226
rect 28030 27174 28888 27226
rect 1104 27152 28888 27174
rect 1578 27072 1584 27124
rect 1636 27112 1642 27124
rect 1636 27084 6914 27112
rect 1636 27072 1642 27084
rect 6886 27044 6914 27084
rect 10962 27072 10968 27124
rect 11020 27112 11026 27124
rect 11057 27115 11115 27121
rect 11057 27112 11069 27115
rect 11020 27084 11069 27112
rect 11020 27072 11026 27084
rect 11057 27081 11069 27084
rect 11103 27081 11115 27115
rect 11057 27075 11115 27081
rect 11422 27072 11428 27124
rect 11480 27112 11486 27124
rect 11977 27115 12035 27121
rect 11977 27112 11989 27115
rect 11480 27084 11989 27112
rect 11480 27072 11486 27084
rect 11977 27081 11989 27084
rect 12023 27081 12035 27115
rect 11977 27075 12035 27081
rect 13262 27044 13268 27056
rect 6886 27016 13268 27044
rect 13262 27004 13268 27016
rect 13320 27004 13326 27056
rect 10965 26979 11023 26985
rect 10965 26945 10977 26979
rect 11011 26945 11023 26979
rect 10965 26939 11023 26945
rect 11885 26979 11943 26985
rect 11885 26945 11897 26979
rect 11931 26976 11943 26979
rect 12250 26976 12256 26988
rect 11931 26948 12256 26976
rect 11931 26945 11943 26948
rect 11885 26939 11943 26945
rect 9214 26800 9220 26852
rect 9272 26840 9278 26852
rect 10980 26840 11008 26939
rect 12250 26936 12256 26948
rect 12308 26936 12314 26988
rect 12434 26936 12440 26988
rect 12492 26976 12498 26988
rect 12529 26979 12587 26985
rect 12529 26976 12541 26979
rect 12492 26948 12541 26976
rect 12492 26936 12498 26948
rect 12529 26945 12541 26948
rect 12575 26945 12587 26979
rect 12529 26939 12587 26945
rect 21358 26936 21364 26988
rect 21416 26976 21422 26988
rect 28077 26979 28135 26985
rect 28077 26976 28089 26979
rect 21416 26948 28089 26976
rect 21416 26936 21422 26948
rect 28077 26945 28089 26948
rect 28123 26945 28135 26979
rect 28077 26939 28135 26945
rect 11241 26911 11299 26917
rect 11241 26877 11253 26911
rect 11287 26908 11299 26911
rect 12158 26908 12164 26920
rect 11287 26880 12164 26908
rect 11287 26877 11299 26880
rect 11241 26871 11299 26877
rect 12158 26868 12164 26880
rect 12216 26868 12222 26920
rect 28350 26868 28356 26920
rect 28408 26868 28414 26920
rect 21266 26840 21272 26852
rect 9272 26812 21272 26840
rect 9272 26800 9278 26812
rect 21266 26800 21272 26812
rect 21324 26800 21330 26852
rect 10594 26732 10600 26784
rect 10652 26732 10658 26784
rect 11422 26732 11428 26784
rect 11480 26772 11486 26784
rect 11517 26775 11575 26781
rect 11517 26772 11529 26775
rect 11480 26744 11529 26772
rect 11480 26732 11486 26744
rect 11517 26741 11529 26744
rect 11563 26741 11575 26775
rect 11517 26735 11575 26741
rect 12066 26732 12072 26784
rect 12124 26772 12130 26784
rect 12345 26775 12403 26781
rect 12345 26772 12357 26775
rect 12124 26744 12357 26772
rect 12124 26732 12130 26744
rect 12345 26741 12357 26744
rect 12391 26741 12403 26775
rect 12345 26735 12403 26741
rect 1104 26682 28888 26704
rect 1104 26630 2918 26682
rect 2970 26630 2982 26682
rect 3034 26630 3046 26682
rect 3098 26630 3110 26682
rect 3162 26630 3174 26682
rect 3226 26630 3238 26682
rect 3290 26630 10918 26682
rect 10970 26630 10982 26682
rect 11034 26630 11046 26682
rect 11098 26630 11110 26682
rect 11162 26630 11174 26682
rect 11226 26630 11238 26682
rect 11290 26630 18918 26682
rect 18970 26630 18982 26682
rect 19034 26630 19046 26682
rect 19098 26630 19110 26682
rect 19162 26630 19174 26682
rect 19226 26630 19238 26682
rect 19290 26630 26918 26682
rect 26970 26630 26982 26682
rect 27034 26630 27046 26682
rect 27098 26630 27110 26682
rect 27162 26630 27174 26682
rect 27226 26630 27238 26682
rect 27290 26630 28888 26682
rect 1104 26608 28888 26630
rect 9214 26577 9220 26580
rect 9171 26571 9220 26577
rect 9171 26537 9183 26571
rect 9217 26537 9220 26571
rect 9171 26531 9220 26537
rect 9214 26528 9220 26531
rect 9272 26528 9278 26580
rect 1581 26503 1639 26509
rect 1581 26469 1593 26503
rect 1627 26500 1639 26503
rect 1627 26472 6914 26500
rect 1627 26469 1639 26472
rect 1581 26463 1639 26469
rect 6886 26432 6914 26472
rect 10410 26432 10416 26444
rect 6886 26404 10416 26432
rect 10410 26392 10416 26404
rect 10468 26392 10474 26444
rect 10594 26392 10600 26444
rect 10652 26392 10658 26444
rect 11422 26392 11428 26444
rect 11480 26392 11486 26444
rect 12158 26392 12164 26444
rect 12216 26432 12222 26444
rect 13541 26435 13599 26441
rect 13541 26432 13553 26435
rect 12216 26404 13553 26432
rect 12216 26392 12222 26404
rect 13541 26401 13553 26404
rect 13587 26401 13599 26435
rect 13541 26395 13599 26401
rect 842 26324 848 26376
rect 900 26364 906 26376
rect 1397 26367 1455 26373
rect 1397 26364 1409 26367
rect 900 26336 1409 26364
rect 900 26324 906 26336
rect 1397 26333 1409 26336
rect 1443 26333 1455 26367
rect 1397 26327 1455 26333
rect 10965 26367 11023 26373
rect 10965 26333 10977 26367
rect 11011 26364 11023 26367
rect 11057 26367 11115 26373
rect 11057 26364 11069 26367
rect 11011 26336 11069 26364
rect 11011 26333 11023 26336
rect 10965 26327 11023 26333
rect 11057 26333 11069 26336
rect 11103 26364 11115 26367
rect 11330 26364 11336 26376
rect 11103 26336 11336 26364
rect 11103 26333 11115 26336
rect 11057 26327 11115 26333
rect 11330 26324 11336 26336
rect 11388 26324 11394 26376
rect 12250 26324 12256 26376
rect 12308 26364 12314 26376
rect 12851 26367 12909 26373
rect 12851 26364 12863 26367
rect 12308 26336 12863 26364
rect 12308 26324 12314 26336
rect 12851 26333 12863 26336
rect 12897 26364 12909 26367
rect 21358 26364 21364 26376
rect 12897 26336 21364 26364
rect 12897 26333 12909 26336
rect 12851 26327 12909 26333
rect 21358 26324 21364 26336
rect 21416 26324 21422 26376
rect 28077 26367 28135 26373
rect 28077 26364 28089 26367
rect 26206 26336 28089 26364
rect 10258 26268 10364 26296
rect 10336 26228 10364 26268
rect 11716 26268 11822 26296
rect 11716 26228 11744 26268
rect 13262 26256 13268 26308
rect 13320 26256 13326 26308
rect 13357 26299 13415 26305
rect 13357 26265 13369 26299
rect 13403 26296 13415 26299
rect 13538 26296 13544 26308
rect 13403 26268 13544 26296
rect 13403 26265 13415 26268
rect 13357 26259 13415 26265
rect 13538 26256 13544 26268
rect 13596 26296 13602 26308
rect 26206 26296 26234 26336
rect 28077 26333 28089 26336
rect 28123 26333 28135 26367
rect 28077 26327 28135 26333
rect 13596 26268 26234 26296
rect 13596 26256 13602 26268
rect 28350 26256 28356 26308
rect 28408 26256 28414 26308
rect 12066 26228 12072 26240
rect 10336 26200 12072 26228
rect 12066 26188 12072 26200
rect 12124 26188 12130 26240
rect 12986 26188 12992 26240
rect 13044 26188 13050 26240
rect 13280 26228 13308 26256
rect 13449 26231 13507 26237
rect 13449 26228 13461 26231
rect 13280 26200 13461 26228
rect 13449 26197 13461 26200
rect 13495 26197 13507 26231
rect 13449 26191 13507 26197
rect 1104 26138 28888 26160
rect 1104 26086 3658 26138
rect 3710 26086 3722 26138
rect 3774 26086 3786 26138
rect 3838 26086 3850 26138
rect 3902 26086 3914 26138
rect 3966 26086 3978 26138
rect 4030 26086 11658 26138
rect 11710 26086 11722 26138
rect 11774 26086 11786 26138
rect 11838 26086 11850 26138
rect 11902 26086 11914 26138
rect 11966 26086 11978 26138
rect 12030 26086 19658 26138
rect 19710 26086 19722 26138
rect 19774 26086 19786 26138
rect 19838 26086 19850 26138
rect 19902 26086 19914 26138
rect 19966 26086 19978 26138
rect 20030 26086 27658 26138
rect 27710 26086 27722 26138
rect 27774 26086 27786 26138
rect 27838 26086 27850 26138
rect 27902 26086 27914 26138
rect 27966 26086 27978 26138
rect 28030 26086 28888 26138
rect 1104 26064 28888 26086
rect 10410 25984 10416 26036
rect 10468 26024 10474 26036
rect 10873 26027 10931 26033
rect 10873 26024 10885 26027
rect 10468 25996 10885 26024
rect 10468 25984 10474 25996
rect 10873 25993 10885 25996
rect 10919 25993 10931 26027
rect 10873 25987 10931 25993
rect 12066 25984 12072 26036
rect 12124 26024 12130 26036
rect 13538 26033 13544 26036
rect 13495 26027 13544 26033
rect 12124 25996 12388 26024
rect 12124 25984 12130 25996
rect 12360 25956 12388 25996
rect 13495 25993 13507 26027
rect 13541 25993 13544 26027
rect 13495 25987 13544 25993
rect 13538 25984 13544 25987
rect 13596 25984 13602 26036
rect 12360 25928 12466 25956
rect 842 25848 848 25900
rect 900 25888 906 25900
rect 1397 25891 1455 25897
rect 1397 25888 1409 25891
rect 900 25860 1409 25888
rect 900 25848 906 25860
rect 1397 25857 1409 25860
rect 1443 25857 1455 25891
rect 1397 25851 1455 25857
rect 10965 25891 11023 25897
rect 10965 25857 10977 25891
rect 11011 25888 11023 25891
rect 11606 25888 11612 25900
rect 11011 25860 11612 25888
rect 11011 25857 11023 25860
rect 10965 25851 11023 25857
rect 11606 25848 11612 25860
rect 11664 25848 11670 25900
rect 10781 25823 10839 25829
rect 10781 25789 10793 25823
rect 10827 25789 10839 25823
rect 10781 25783 10839 25789
rect 10796 25752 10824 25783
rect 11330 25780 11336 25832
rect 11388 25820 11394 25832
rect 11701 25823 11759 25829
rect 11701 25820 11713 25823
rect 11388 25792 11713 25820
rect 11388 25780 11394 25792
rect 11701 25789 11713 25792
rect 11747 25789 11759 25823
rect 11701 25783 11759 25789
rect 12069 25823 12127 25829
rect 12069 25789 12081 25823
rect 12115 25820 12127 25823
rect 12986 25820 12992 25832
rect 12115 25792 12992 25820
rect 12115 25789 12127 25792
rect 12069 25783 12127 25789
rect 12986 25780 12992 25792
rect 13044 25780 13050 25832
rect 10796 25724 11744 25752
rect 1581 25687 1639 25693
rect 1581 25653 1593 25687
rect 1627 25684 1639 25687
rect 10594 25684 10600 25696
rect 1627 25656 10600 25684
rect 1627 25653 1639 25656
rect 1581 25647 1639 25653
rect 10594 25644 10600 25656
rect 10652 25644 10658 25696
rect 11333 25687 11391 25693
rect 11333 25653 11345 25687
rect 11379 25684 11391 25687
rect 11422 25684 11428 25696
rect 11379 25656 11428 25684
rect 11379 25653 11391 25656
rect 11333 25647 11391 25653
rect 11422 25644 11428 25656
rect 11480 25644 11486 25696
rect 11716 25684 11744 25724
rect 12066 25684 12072 25696
rect 11716 25656 12072 25684
rect 12066 25644 12072 25656
rect 12124 25644 12130 25696
rect 1104 25594 28888 25616
rect 1104 25542 2918 25594
rect 2970 25542 2982 25594
rect 3034 25542 3046 25594
rect 3098 25542 3110 25594
rect 3162 25542 3174 25594
rect 3226 25542 3238 25594
rect 3290 25542 10918 25594
rect 10970 25542 10982 25594
rect 11034 25542 11046 25594
rect 11098 25542 11110 25594
rect 11162 25542 11174 25594
rect 11226 25542 11238 25594
rect 11290 25542 18918 25594
rect 18970 25542 18982 25594
rect 19034 25542 19046 25594
rect 19098 25542 19110 25594
rect 19162 25542 19174 25594
rect 19226 25542 19238 25594
rect 19290 25542 26918 25594
rect 26970 25542 26982 25594
rect 27034 25542 27046 25594
rect 27098 25542 27110 25594
rect 27162 25542 27174 25594
rect 27226 25542 27238 25594
rect 27290 25542 28888 25594
rect 1104 25520 28888 25542
rect 11422 25304 11428 25356
rect 11480 25304 11486 25356
rect 11606 25304 11612 25356
rect 11664 25344 11670 25356
rect 11664 25316 12894 25344
rect 11664 25304 11670 25316
rect 11057 25279 11115 25285
rect 11057 25245 11069 25279
rect 11103 25276 11115 25279
rect 11330 25276 11336 25288
rect 11103 25248 11336 25276
rect 11103 25245 11115 25248
rect 11057 25239 11115 25245
rect 11330 25236 11336 25248
rect 11388 25236 11394 25288
rect 12866 25285 12894 25316
rect 12851 25279 12909 25285
rect 12851 25245 12863 25279
rect 12897 25276 12909 25279
rect 28077 25279 28135 25285
rect 28077 25276 28089 25279
rect 12897 25248 28089 25276
rect 12897 25245 12909 25248
rect 12851 25239 12909 25245
rect 28077 25245 28089 25248
rect 28123 25245 28135 25279
rect 28077 25239 28135 25245
rect 12466 25180 12848 25208
rect 12820 25152 12848 25180
rect 28350 25168 28356 25220
rect 28408 25168 28414 25220
rect 12802 25100 12808 25152
rect 12860 25100 12866 25152
rect 1104 25050 28888 25072
rect 1104 24998 3658 25050
rect 3710 24998 3722 25050
rect 3774 24998 3786 25050
rect 3838 24998 3850 25050
rect 3902 24998 3914 25050
rect 3966 24998 3978 25050
rect 4030 24998 11658 25050
rect 11710 24998 11722 25050
rect 11774 24998 11786 25050
rect 11838 24998 11850 25050
rect 11902 24998 11914 25050
rect 11966 24998 11978 25050
rect 12030 24998 19658 25050
rect 19710 24998 19722 25050
rect 19774 24998 19786 25050
rect 19838 24998 19850 25050
rect 19902 24998 19914 25050
rect 19966 24998 19978 25050
rect 20030 24998 27658 25050
rect 27710 24998 27722 25050
rect 27774 24998 27786 25050
rect 27838 24998 27850 25050
rect 27902 24998 27914 25050
rect 27966 24998 27978 25050
rect 28030 24998 28888 25050
rect 1104 24976 28888 24998
rect 12802 24828 12808 24880
rect 12860 24828 12866 24880
rect 842 24760 848 24812
rect 900 24800 906 24812
rect 1397 24803 1455 24809
rect 1397 24800 1409 24803
rect 900 24772 1409 24800
rect 900 24760 906 24772
rect 1397 24769 1409 24772
rect 1443 24769 1455 24803
rect 1397 24763 1455 24769
rect 13354 24760 13360 24812
rect 13412 24800 13418 24812
rect 13863 24803 13921 24809
rect 13863 24800 13875 24803
rect 13412 24772 13875 24800
rect 13412 24760 13418 24772
rect 13863 24769 13875 24772
rect 13909 24800 13921 24803
rect 28077 24803 28135 24809
rect 28077 24800 28089 24803
rect 13909 24772 28089 24800
rect 13909 24769 13921 24772
rect 13863 24763 13921 24769
rect 28077 24769 28089 24772
rect 28123 24769 28135 24803
rect 28077 24763 28135 24769
rect 11330 24692 11336 24744
rect 11388 24732 11394 24744
rect 12069 24735 12127 24741
rect 12069 24732 12081 24735
rect 11388 24704 12081 24732
rect 11388 24692 11394 24704
rect 12069 24701 12081 24704
rect 12115 24701 12127 24735
rect 12069 24695 12127 24701
rect 12437 24735 12495 24741
rect 12437 24701 12449 24735
rect 12483 24732 12495 24735
rect 12986 24732 12992 24744
rect 12483 24704 12992 24732
rect 12483 24701 12495 24704
rect 12437 24695 12495 24701
rect 12986 24692 12992 24704
rect 13044 24692 13050 24744
rect 28350 24692 28356 24744
rect 28408 24692 28414 24744
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24596 1639 24599
rect 11422 24596 11428 24608
rect 1627 24568 11428 24596
rect 1627 24565 1639 24568
rect 1581 24559 1639 24565
rect 11422 24556 11428 24568
rect 11480 24556 11486 24608
rect 1104 24506 28888 24528
rect 1104 24454 2918 24506
rect 2970 24454 2982 24506
rect 3034 24454 3046 24506
rect 3098 24454 3110 24506
rect 3162 24454 3174 24506
rect 3226 24454 3238 24506
rect 3290 24454 10918 24506
rect 10970 24454 10982 24506
rect 11034 24454 11046 24506
rect 11098 24454 11110 24506
rect 11162 24454 11174 24506
rect 11226 24454 11238 24506
rect 11290 24454 18918 24506
rect 18970 24454 18982 24506
rect 19034 24454 19046 24506
rect 19098 24454 19110 24506
rect 19162 24454 19174 24506
rect 19226 24454 19238 24506
rect 19290 24454 26918 24506
rect 26970 24454 26982 24506
rect 27034 24454 27046 24506
rect 27098 24454 27110 24506
rect 27162 24454 27174 24506
rect 27226 24454 27238 24506
rect 27290 24454 28888 24506
rect 1104 24432 28888 24454
rect 12986 24352 12992 24404
rect 13044 24352 13050 24404
rect 12250 24284 12256 24336
rect 12308 24324 12314 24336
rect 12308 24296 13584 24324
rect 12308 24284 12314 24296
rect 10594 24216 10600 24268
rect 10652 24256 10658 24268
rect 13556 24265 13584 24296
rect 13449 24259 13507 24265
rect 13449 24256 13461 24259
rect 10652 24228 13461 24256
rect 10652 24216 10658 24228
rect 13449 24225 13461 24228
rect 13495 24225 13507 24259
rect 13449 24219 13507 24225
rect 13541 24259 13599 24265
rect 13541 24225 13553 24259
rect 13587 24225 13599 24259
rect 13541 24219 13599 24225
rect 842 24148 848 24200
rect 900 24188 906 24200
rect 1397 24191 1455 24197
rect 1397 24188 1409 24191
rect 900 24160 1409 24188
rect 900 24148 906 24160
rect 1397 24157 1409 24160
rect 1443 24157 1455 24191
rect 1397 24151 1455 24157
rect 11057 24191 11115 24197
rect 11057 24157 11069 24191
rect 11103 24188 11115 24191
rect 11330 24188 11336 24200
rect 11103 24160 11336 24188
rect 11103 24157 11115 24160
rect 11057 24151 11115 24157
rect 11330 24148 11336 24160
rect 11388 24148 11394 24200
rect 11425 24191 11483 24197
rect 11425 24157 11437 24191
rect 11471 24188 11483 24191
rect 11514 24188 11520 24200
rect 11471 24160 11520 24188
rect 11471 24157 11483 24160
rect 11425 24151 11483 24157
rect 11514 24148 11520 24160
rect 11572 24148 11578 24200
rect 13354 24148 13360 24200
rect 13412 24148 13418 24200
rect 12466 24092 12572 24120
rect 1578 24012 1584 24064
rect 1636 24012 1642 24064
rect 12544 24052 12572 24092
rect 12618 24080 12624 24132
rect 12676 24120 12682 24132
rect 12851 24123 12909 24129
rect 12851 24120 12863 24123
rect 12676 24092 12863 24120
rect 12676 24080 12682 24092
rect 12851 24089 12863 24092
rect 12897 24120 12909 24123
rect 28074 24120 28080 24132
rect 12897 24092 28080 24120
rect 12897 24089 12909 24092
rect 12851 24083 12909 24089
rect 28074 24080 28080 24092
rect 28132 24080 28138 24132
rect 12710 24052 12716 24064
rect 12544 24024 12716 24052
rect 12710 24012 12716 24024
rect 12768 24012 12774 24064
rect 1104 23962 28888 23984
rect 1104 23910 3658 23962
rect 3710 23910 3722 23962
rect 3774 23910 3786 23962
rect 3838 23910 3850 23962
rect 3902 23910 3914 23962
rect 3966 23910 3978 23962
rect 4030 23910 11658 23962
rect 11710 23910 11722 23962
rect 11774 23910 11786 23962
rect 11838 23910 11850 23962
rect 11902 23910 11914 23962
rect 11966 23910 11978 23962
rect 12030 23910 19658 23962
rect 19710 23910 19722 23962
rect 19774 23910 19786 23962
rect 19838 23910 19850 23962
rect 19902 23910 19914 23962
rect 19966 23910 19978 23962
rect 20030 23910 27658 23962
rect 27710 23910 27722 23962
rect 27774 23910 27786 23962
rect 27838 23910 27850 23962
rect 27902 23910 27914 23962
rect 27966 23910 27978 23962
rect 28030 23910 28888 23962
rect 1104 23888 28888 23910
rect 1578 23808 1584 23860
rect 1636 23848 1642 23860
rect 1636 23820 6914 23848
rect 1636 23808 1642 23820
rect 6886 23712 6914 23820
rect 11514 23808 11520 23860
rect 11572 23808 11578 23860
rect 11885 23851 11943 23857
rect 11885 23817 11897 23851
rect 11931 23848 11943 23851
rect 12618 23848 12624 23860
rect 11931 23820 12624 23848
rect 11931 23817 11943 23820
rect 11885 23811 11943 23817
rect 12618 23808 12624 23820
rect 12676 23808 12682 23860
rect 11422 23740 11428 23792
rect 11480 23780 11486 23792
rect 11977 23783 12035 23789
rect 11977 23780 11989 23783
rect 11480 23752 11989 23780
rect 11480 23740 11486 23752
rect 11977 23749 11989 23752
rect 12023 23749 12035 23783
rect 11977 23743 12035 23749
rect 14550 23712 14556 23724
rect 6886 23684 14556 23712
rect 14550 23672 14556 23684
rect 14608 23672 14614 23724
rect 28074 23672 28080 23724
rect 28132 23672 28138 23724
rect 12066 23604 12072 23656
rect 12124 23604 12130 23656
rect 28350 23604 28356 23656
rect 28408 23604 28414 23656
rect 1104 23418 28888 23440
rect 1104 23366 2918 23418
rect 2970 23366 2982 23418
rect 3034 23366 3046 23418
rect 3098 23366 3110 23418
rect 3162 23366 3174 23418
rect 3226 23366 3238 23418
rect 3290 23366 10918 23418
rect 10970 23366 10982 23418
rect 11034 23366 11046 23418
rect 11098 23366 11110 23418
rect 11162 23366 11174 23418
rect 11226 23366 11238 23418
rect 11290 23366 18918 23418
rect 18970 23366 18982 23418
rect 19034 23366 19046 23418
rect 19098 23366 19110 23418
rect 19162 23366 19174 23418
rect 19226 23366 19238 23418
rect 19290 23366 26918 23418
rect 26970 23366 26982 23418
rect 27034 23366 27046 23418
rect 27098 23366 27110 23418
rect 27162 23366 27174 23418
rect 27226 23366 27238 23418
rect 27290 23366 28888 23418
rect 1104 23344 28888 23366
rect 11425 23239 11483 23245
rect 11425 23205 11437 23239
rect 11471 23236 11483 23239
rect 12066 23236 12072 23248
rect 11471 23208 12072 23236
rect 11471 23205 11483 23208
rect 11425 23199 11483 23205
rect 12066 23196 12072 23208
rect 12124 23236 12130 23248
rect 12124 23208 14688 23236
rect 12124 23196 12130 23208
rect 14660 23180 14688 23208
rect 14550 23128 14556 23180
rect 14608 23128 14614 23180
rect 14642 23128 14648 23180
rect 14700 23128 14706 23180
rect 842 23060 848 23112
rect 900 23100 906 23112
rect 1397 23103 1455 23109
rect 1397 23100 1409 23103
rect 900 23072 1409 23100
rect 900 23060 906 23072
rect 1397 23069 1409 23072
rect 1443 23069 1455 23103
rect 1397 23063 1455 23069
rect 11241 23103 11299 23109
rect 11241 23069 11253 23103
rect 11287 23100 11299 23103
rect 12158 23100 12164 23112
rect 11287 23072 12164 23100
rect 11287 23069 11299 23072
rect 11241 23063 11299 23069
rect 12158 23060 12164 23072
rect 12216 23060 12222 23112
rect 14461 23103 14519 23109
rect 14461 23069 14473 23103
rect 14507 23100 14519 23103
rect 14918 23100 14924 23112
rect 14507 23072 14924 23100
rect 14507 23069 14519 23072
rect 14461 23063 14519 23069
rect 14918 23060 14924 23072
rect 14976 23100 14982 23112
rect 28077 23103 28135 23109
rect 28077 23100 28089 23103
rect 14976 23072 28089 23100
rect 14976 23060 14982 23072
rect 28077 23069 28089 23072
rect 28123 23069 28135 23103
rect 28077 23063 28135 23069
rect 11514 22992 11520 23044
rect 11572 22992 11578 23044
rect 28350 22992 28356 23044
rect 28408 22992 28414 23044
rect 1581 22967 1639 22973
rect 1581 22933 1593 22967
rect 1627 22964 1639 22967
rect 11146 22964 11152 22976
rect 1627 22936 11152 22964
rect 1627 22933 1639 22936
rect 1581 22927 1639 22933
rect 11146 22924 11152 22936
rect 11204 22924 11210 22976
rect 12989 22967 13047 22973
rect 12989 22933 13001 22967
rect 13035 22964 13047 22967
rect 13078 22964 13084 22976
rect 13035 22936 13084 22964
rect 13035 22933 13047 22936
rect 12989 22927 13047 22933
rect 13078 22924 13084 22936
rect 13136 22924 13142 22976
rect 13446 22924 13452 22976
rect 13504 22964 13510 22976
rect 14093 22967 14151 22973
rect 14093 22964 14105 22967
rect 13504 22936 14105 22964
rect 13504 22924 13510 22936
rect 14093 22933 14105 22936
rect 14139 22933 14151 22967
rect 14093 22927 14151 22933
rect 1104 22874 28888 22896
rect 1104 22822 3658 22874
rect 3710 22822 3722 22874
rect 3774 22822 3786 22874
rect 3838 22822 3850 22874
rect 3902 22822 3914 22874
rect 3966 22822 3978 22874
rect 4030 22822 11658 22874
rect 11710 22822 11722 22874
rect 11774 22822 11786 22874
rect 11838 22822 11850 22874
rect 11902 22822 11914 22874
rect 11966 22822 11978 22874
rect 12030 22822 19658 22874
rect 19710 22822 19722 22874
rect 19774 22822 19786 22874
rect 19838 22822 19850 22874
rect 19902 22822 19914 22874
rect 19966 22822 19978 22874
rect 20030 22822 27658 22874
rect 27710 22822 27722 22874
rect 27774 22822 27786 22874
rect 27838 22822 27850 22874
rect 27902 22822 27914 22874
rect 27966 22822 27978 22874
rect 28030 22822 28888 22874
rect 1104 22800 28888 22822
rect 11146 22720 11152 22772
rect 11204 22760 11210 22772
rect 14918 22769 14924 22772
rect 11977 22763 12035 22769
rect 11977 22760 11989 22763
rect 11204 22732 11989 22760
rect 11204 22720 11210 22732
rect 11977 22729 11989 22732
rect 12023 22729 12035 22763
rect 11977 22723 12035 22729
rect 14875 22763 14924 22769
rect 14875 22729 14887 22763
rect 14921 22729 14924 22763
rect 14875 22723 14924 22729
rect 14918 22720 14924 22723
rect 14976 22720 14982 22772
rect 11885 22695 11943 22701
rect 11885 22661 11897 22695
rect 11931 22692 11943 22695
rect 12618 22692 12624 22704
rect 11931 22664 12624 22692
rect 11931 22661 11943 22664
rect 11885 22655 11943 22661
rect 12618 22652 12624 22664
rect 12676 22652 12682 22704
rect 13814 22652 13820 22704
rect 13872 22652 13878 22704
rect 842 22584 848 22636
rect 900 22624 906 22636
rect 1397 22627 1455 22633
rect 1397 22624 1409 22627
rect 900 22596 1409 22624
rect 900 22584 906 22596
rect 1397 22593 1409 22596
rect 1443 22593 1455 22627
rect 1397 22587 1455 22593
rect 12434 22584 12440 22636
rect 12492 22584 12498 22636
rect 13446 22584 13452 22636
rect 13504 22584 13510 22636
rect 12066 22516 12072 22568
rect 12124 22516 12130 22568
rect 13078 22516 13084 22568
rect 13136 22516 13142 22568
rect 12621 22491 12679 22497
rect 12621 22457 12633 22491
rect 12667 22488 12679 22491
rect 12710 22488 12716 22500
rect 12667 22460 12716 22488
rect 12667 22457 12679 22460
rect 12621 22451 12679 22457
rect 12710 22448 12716 22460
rect 12768 22448 12774 22500
rect 1578 22380 1584 22432
rect 1636 22380 1642 22432
rect 11422 22380 11428 22432
rect 11480 22420 11486 22432
rect 11517 22423 11575 22429
rect 11517 22420 11529 22423
rect 11480 22392 11529 22420
rect 11480 22380 11486 22392
rect 11517 22389 11529 22392
rect 11563 22389 11575 22423
rect 11517 22383 11575 22389
rect 1104 22330 28888 22352
rect 1104 22278 2918 22330
rect 2970 22278 2982 22330
rect 3034 22278 3046 22330
rect 3098 22278 3110 22330
rect 3162 22278 3174 22330
rect 3226 22278 3238 22330
rect 3290 22278 10918 22330
rect 10970 22278 10982 22330
rect 11034 22278 11046 22330
rect 11098 22278 11110 22330
rect 11162 22278 11174 22330
rect 11226 22278 11238 22330
rect 11290 22278 18918 22330
rect 18970 22278 18982 22330
rect 19034 22278 19046 22330
rect 19098 22278 19110 22330
rect 19162 22278 19174 22330
rect 19226 22278 19238 22330
rect 19290 22278 26918 22330
rect 26970 22278 26982 22330
rect 27034 22278 27046 22330
rect 27098 22278 27110 22330
rect 27162 22278 27174 22330
rect 27226 22278 27238 22330
rect 27290 22278 28888 22330
rect 1104 22256 28888 22278
rect 1578 22176 1584 22228
rect 1636 22216 1642 22228
rect 1636 22188 14596 22216
rect 1636 22176 1642 22188
rect 11057 22083 11115 22089
rect 11057 22049 11069 22083
rect 11103 22080 11115 22083
rect 11330 22080 11336 22092
rect 11103 22052 11336 22080
rect 11103 22049 11115 22052
rect 11057 22043 11115 22049
rect 11330 22040 11336 22052
rect 11388 22080 11394 22092
rect 13078 22080 13084 22092
rect 11388 22052 13084 22080
rect 11388 22040 11394 22052
rect 13078 22040 13084 22052
rect 13136 22040 13142 22092
rect 14568 22089 14596 22188
rect 14642 22108 14648 22160
rect 14700 22148 14706 22160
rect 14700 22120 14780 22148
rect 14700 22108 14706 22120
rect 14752 22089 14780 22120
rect 14553 22083 14611 22089
rect 14553 22049 14565 22083
rect 14599 22049 14611 22083
rect 14553 22043 14611 22049
rect 14737 22083 14795 22089
rect 14737 22049 14749 22083
rect 14783 22049 14795 22083
rect 14737 22043 14795 22049
rect 11422 21972 11428 22024
rect 11480 21972 11486 22024
rect 12710 22012 12716 22024
rect 12452 21984 12716 22012
rect 12452 21930 12480 21984
rect 12710 21972 12716 21984
rect 12768 22012 12774 22024
rect 13722 22012 13728 22024
rect 12768 21984 13728 22012
rect 12768 21972 12774 21984
rect 13722 21972 13728 21984
rect 13780 21972 13786 22024
rect 28077 22015 28135 22021
rect 28077 22012 28089 22015
rect 26206 21984 28089 22012
rect 12618 21904 12624 21956
rect 12676 21944 12682 21956
rect 12851 21947 12909 21953
rect 12851 21944 12863 21947
rect 12676 21916 12863 21944
rect 12676 21904 12682 21916
rect 12851 21913 12863 21916
rect 12897 21944 12909 21947
rect 14461 21947 14519 21953
rect 12897 21916 14228 21944
rect 12897 21913 12909 21916
rect 12851 21907 12909 21913
rect 13446 21836 13452 21888
rect 13504 21876 13510 21888
rect 14093 21879 14151 21885
rect 14093 21876 14105 21879
rect 13504 21848 14105 21876
rect 13504 21836 13510 21848
rect 14093 21845 14105 21848
rect 14139 21845 14151 21879
rect 14200 21876 14228 21916
rect 14461 21913 14473 21947
rect 14507 21944 14519 21947
rect 14826 21944 14832 21956
rect 14507 21916 14832 21944
rect 14507 21913 14519 21916
rect 14461 21907 14519 21913
rect 14826 21904 14832 21916
rect 14884 21944 14890 21956
rect 17862 21944 17868 21956
rect 14884 21916 17868 21944
rect 14884 21904 14890 21916
rect 17862 21904 17868 21916
rect 17920 21904 17926 21956
rect 26206 21876 26234 21984
rect 28077 21981 28089 21984
rect 28123 21981 28135 22015
rect 28077 21975 28135 21981
rect 28350 21904 28356 21956
rect 28408 21904 28414 21956
rect 14200 21848 26234 21876
rect 14093 21839 14151 21845
rect 1104 21786 28888 21808
rect 1104 21734 3658 21786
rect 3710 21734 3722 21786
rect 3774 21734 3786 21786
rect 3838 21734 3850 21786
rect 3902 21734 3914 21786
rect 3966 21734 3978 21786
rect 4030 21734 11658 21786
rect 11710 21734 11722 21786
rect 11774 21734 11786 21786
rect 11838 21734 11850 21786
rect 11902 21734 11914 21786
rect 11966 21734 11978 21786
rect 12030 21734 19658 21786
rect 19710 21734 19722 21786
rect 19774 21734 19786 21786
rect 19838 21734 19850 21786
rect 19902 21734 19914 21786
rect 19966 21734 19978 21786
rect 20030 21734 27658 21786
rect 27710 21734 27722 21786
rect 27774 21734 27786 21786
rect 27838 21734 27850 21786
rect 27902 21734 27914 21786
rect 27966 21734 27978 21786
rect 28030 21734 28888 21786
rect 1104 21712 28888 21734
rect 13722 21632 13728 21684
rect 13780 21632 13786 21684
rect 14826 21632 14832 21684
rect 14884 21681 14890 21684
rect 14884 21675 14933 21681
rect 14884 21641 14887 21675
rect 14921 21641 14933 21675
rect 14884 21635 14933 21641
rect 14884 21632 14890 21635
rect 13740 21604 13768 21632
rect 13740 21576 13846 21604
rect 1394 21496 1400 21548
rect 1452 21496 1458 21548
rect 13078 21496 13084 21548
rect 13136 21496 13142 21548
rect 13446 21496 13452 21548
rect 13504 21496 13510 21548
rect 17862 21496 17868 21548
rect 17920 21536 17926 21548
rect 28077 21539 28135 21545
rect 28077 21536 28089 21539
rect 17920 21508 28089 21536
rect 17920 21496 17926 21508
rect 28077 21505 28089 21508
rect 28123 21505 28135 21539
rect 28077 21499 28135 21505
rect 28350 21428 28356 21480
rect 28408 21428 28414 21480
rect 1581 21335 1639 21341
rect 1581 21301 1593 21335
rect 1627 21332 1639 21335
rect 14550 21332 14556 21344
rect 1627 21304 14556 21332
rect 1627 21301 1639 21304
rect 1581 21295 1639 21301
rect 14550 21292 14556 21304
rect 14608 21292 14614 21344
rect 1104 21242 28888 21264
rect 1104 21190 2918 21242
rect 2970 21190 2982 21242
rect 3034 21190 3046 21242
rect 3098 21190 3110 21242
rect 3162 21190 3174 21242
rect 3226 21190 3238 21242
rect 3290 21190 10918 21242
rect 10970 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 11238 21242
rect 11290 21190 18918 21242
rect 18970 21190 18982 21242
rect 19034 21190 19046 21242
rect 19098 21190 19110 21242
rect 19162 21190 19174 21242
rect 19226 21190 19238 21242
rect 19290 21190 26918 21242
rect 26970 21190 26982 21242
rect 27034 21190 27046 21242
rect 27098 21190 27110 21242
rect 27162 21190 27174 21242
rect 27226 21190 27238 21242
rect 27290 21190 28888 21242
rect 1104 21168 28888 21190
rect 12158 21020 12164 21072
rect 12216 21060 12222 21072
rect 12216 21032 14688 21060
rect 12216 21020 12222 21032
rect 14550 20952 14556 21004
rect 14608 20952 14614 21004
rect 14660 21001 14688 21032
rect 14645 20995 14703 21001
rect 14645 20961 14657 20995
rect 14691 20961 14703 20995
rect 14645 20955 14703 20961
rect 1394 20884 1400 20936
rect 1452 20884 1458 20936
rect 14461 20859 14519 20865
rect 14461 20825 14473 20859
rect 14507 20856 14519 20859
rect 14642 20856 14648 20868
rect 14507 20828 14648 20856
rect 14507 20825 14519 20828
rect 14461 20819 14519 20825
rect 14642 20816 14648 20828
rect 14700 20816 14706 20868
rect 1581 20791 1639 20797
rect 1581 20757 1593 20791
rect 1627 20788 1639 20791
rect 11330 20788 11336 20800
rect 1627 20760 11336 20788
rect 1627 20757 1639 20760
rect 1581 20751 1639 20757
rect 11330 20748 11336 20760
rect 11388 20748 11394 20800
rect 13906 20748 13912 20800
rect 13964 20788 13970 20800
rect 14093 20791 14151 20797
rect 14093 20788 14105 20791
rect 13964 20760 14105 20788
rect 13964 20748 13970 20760
rect 14093 20757 14105 20760
rect 14139 20757 14151 20791
rect 14093 20751 14151 20757
rect 1104 20698 28888 20720
rect 1104 20646 3658 20698
rect 3710 20646 3722 20698
rect 3774 20646 3786 20698
rect 3838 20646 3850 20698
rect 3902 20646 3914 20698
rect 3966 20646 3978 20698
rect 4030 20646 11658 20698
rect 11710 20646 11722 20698
rect 11774 20646 11786 20698
rect 11838 20646 11850 20698
rect 11902 20646 11914 20698
rect 11966 20646 11978 20698
rect 12030 20646 19658 20698
rect 19710 20646 19722 20698
rect 19774 20646 19786 20698
rect 19838 20646 19850 20698
rect 19902 20646 19914 20698
rect 19966 20646 19978 20698
rect 20030 20646 27658 20698
rect 27710 20646 27722 20698
rect 27774 20646 27786 20698
rect 27838 20646 27850 20698
rect 27902 20646 27914 20698
rect 27966 20646 27978 20698
rect 28030 20646 28888 20698
rect 1104 20624 28888 20646
rect 12434 20544 12440 20596
rect 12492 20584 12498 20596
rect 12492 20556 13768 20584
rect 12492 20544 12498 20556
rect 13740 20516 13768 20556
rect 13740 20488 13846 20516
rect 14642 20408 14648 20460
rect 14700 20448 14706 20460
rect 14875 20451 14933 20457
rect 14875 20448 14887 20451
rect 14700 20420 14887 20448
rect 14700 20408 14706 20420
rect 14875 20417 14887 20420
rect 14921 20448 14933 20451
rect 28077 20451 28135 20457
rect 28077 20448 28089 20451
rect 14921 20420 28089 20448
rect 14921 20417 14933 20420
rect 14875 20411 14933 20417
rect 28077 20417 28089 20420
rect 28123 20417 28135 20451
rect 28077 20411 28135 20417
rect 12342 20340 12348 20392
rect 12400 20380 12406 20392
rect 13081 20383 13139 20389
rect 13081 20380 13093 20383
rect 12400 20352 13093 20380
rect 12400 20340 12406 20352
rect 13081 20349 13093 20352
rect 13127 20349 13139 20383
rect 13081 20343 13139 20349
rect 13449 20383 13507 20389
rect 13449 20349 13461 20383
rect 13495 20380 13507 20383
rect 13906 20380 13912 20392
rect 13495 20352 13912 20380
rect 13495 20349 13507 20352
rect 13449 20343 13507 20349
rect 13906 20340 13912 20352
rect 13964 20340 13970 20392
rect 28350 20340 28356 20392
rect 28408 20340 28414 20392
rect 1104 20154 28888 20176
rect 1104 20102 2918 20154
rect 2970 20102 2982 20154
rect 3034 20102 3046 20154
rect 3098 20102 3110 20154
rect 3162 20102 3174 20154
rect 3226 20102 3238 20154
rect 3290 20102 10918 20154
rect 10970 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 11238 20154
rect 11290 20102 18918 20154
rect 18970 20102 18982 20154
rect 19034 20102 19046 20154
rect 19098 20102 19110 20154
rect 19162 20102 19174 20154
rect 19226 20102 19238 20154
rect 19290 20102 26918 20154
rect 26970 20102 26982 20154
rect 27034 20102 27046 20154
rect 27098 20102 27110 20154
rect 27162 20102 27174 20154
rect 27226 20102 27238 20154
rect 27290 20102 28888 20154
rect 1104 20080 28888 20102
rect 1581 20043 1639 20049
rect 1581 20009 1593 20043
rect 1627 20040 1639 20043
rect 1627 20012 13676 20040
rect 1627 20009 1639 20012
rect 1581 20003 1639 20009
rect 11057 19907 11115 19913
rect 11057 19873 11069 19907
rect 11103 19904 11115 19907
rect 12342 19904 12348 19916
rect 11103 19876 12348 19904
rect 11103 19873 11115 19876
rect 11057 19867 11115 19873
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 13648 19913 13676 20012
rect 13633 19907 13691 19913
rect 13633 19873 13645 19907
rect 13679 19873 13691 19907
rect 13633 19867 13691 19873
rect 13814 19864 13820 19916
rect 13872 19864 13878 19916
rect 1394 19796 1400 19848
rect 1452 19796 1458 19848
rect 11422 19796 11428 19848
rect 11480 19796 11486 19848
rect 12250 19796 12256 19848
rect 12308 19836 12314 19848
rect 12851 19839 12909 19845
rect 12851 19836 12863 19839
rect 12308 19808 12863 19836
rect 12308 19796 12314 19808
rect 12851 19805 12863 19808
rect 12897 19836 12909 19839
rect 28077 19839 28135 19845
rect 28077 19836 28089 19839
rect 12897 19808 28089 19836
rect 12897 19805 12909 19808
rect 12851 19799 12909 19805
rect 28077 19805 28089 19808
rect 28123 19805 28135 19839
rect 28077 19799 28135 19805
rect 12434 19728 12440 19780
rect 12492 19728 12498 19780
rect 28350 19728 28356 19780
rect 28408 19728 28414 19780
rect 12986 19660 12992 19712
rect 13044 19700 13050 19712
rect 13173 19703 13231 19709
rect 13173 19700 13185 19703
rect 13044 19672 13185 19700
rect 13044 19660 13050 19672
rect 13173 19669 13185 19672
rect 13219 19669 13231 19703
rect 13173 19663 13231 19669
rect 13538 19660 13544 19712
rect 13596 19660 13602 19712
rect 1104 19610 28888 19632
rect 1104 19558 3658 19610
rect 3710 19558 3722 19610
rect 3774 19558 3786 19610
rect 3838 19558 3850 19610
rect 3902 19558 3914 19610
rect 3966 19558 3978 19610
rect 4030 19558 11658 19610
rect 11710 19558 11722 19610
rect 11774 19558 11786 19610
rect 11838 19558 11850 19610
rect 11902 19558 11914 19610
rect 11966 19558 11978 19610
rect 12030 19558 19658 19610
rect 19710 19558 19722 19610
rect 19774 19558 19786 19610
rect 19838 19558 19850 19610
rect 19902 19558 19914 19610
rect 19966 19558 19978 19610
rect 20030 19558 27658 19610
rect 27710 19558 27722 19610
rect 27774 19558 27786 19610
rect 27838 19558 27850 19610
rect 27902 19558 27914 19610
rect 27966 19558 27978 19610
rect 28030 19558 28888 19610
rect 1104 19536 28888 19558
rect 1581 19499 1639 19505
rect 1581 19465 1593 19499
rect 1627 19496 1639 19499
rect 1627 19468 6914 19496
rect 1627 19465 1639 19468
rect 1581 19459 1639 19465
rect 842 19320 848 19372
rect 900 19360 906 19372
rect 1397 19363 1455 19369
rect 1397 19360 1409 19363
rect 900 19332 1409 19360
rect 900 19320 906 19332
rect 1397 19329 1409 19332
rect 1443 19329 1455 19363
rect 6886 19360 6914 19468
rect 11422 19456 11428 19508
rect 11480 19496 11486 19508
rect 11517 19499 11575 19505
rect 11517 19496 11529 19499
rect 11480 19468 11529 19496
rect 11480 19456 11486 19468
rect 11517 19465 11529 19468
rect 11563 19465 11575 19499
rect 11517 19459 11575 19465
rect 11885 19499 11943 19505
rect 11885 19465 11897 19499
rect 11931 19496 11943 19499
rect 12250 19496 12256 19508
rect 11931 19468 12256 19496
rect 11931 19465 11943 19468
rect 11885 19459 11943 19465
rect 12250 19456 12256 19468
rect 12308 19456 12314 19508
rect 13538 19456 13544 19508
rect 13596 19496 13602 19508
rect 13596 19468 14136 19496
rect 13596 19456 13602 19468
rect 11330 19388 11336 19440
rect 11388 19428 11394 19440
rect 11977 19431 12035 19437
rect 11977 19428 11989 19431
rect 11388 19400 11989 19428
rect 11388 19388 11394 19400
rect 11977 19397 11989 19400
rect 12023 19397 12035 19431
rect 11977 19391 12035 19397
rect 12268 19400 12756 19428
rect 12268 19360 12296 19400
rect 6886 19332 12296 19360
rect 1397 19323 1455 19329
rect 12342 19320 12348 19372
rect 12400 19360 12406 19372
rect 12621 19363 12679 19369
rect 12621 19360 12633 19363
rect 12400 19332 12633 19360
rect 12400 19320 12406 19332
rect 12621 19329 12633 19332
rect 12667 19329 12679 19363
rect 12728 19360 12756 19400
rect 13722 19388 13728 19440
rect 13780 19388 13786 19440
rect 12728 19332 12940 19360
rect 12621 19323 12679 19329
rect 11422 19252 11428 19304
rect 11480 19292 11486 19304
rect 12069 19295 12127 19301
rect 12069 19292 12081 19295
rect 11480 19264 12081 19292
rect 11480 19252 11486 19264
rect 12069 19261 12081 19264
rect 12115 19292 12127 19295
rect 12158 19292 12164 19304
rect 12115 19264 12164 19292
rect 12115 19261 12127 19264
rect 12069 19255 12127 19261
rect 12158 19252 12164 19264
rect 12216 19252 12222 19304
rect 12912 19292 12940 19332
rect 12986 19320 12992 19372
rect 13044 19320 13050 19372
rect 14108 19360 14136 19468
rect 14415 19363 14473 19369
rect 14415 19360 14427 19363
rect 14108 19332 14427 19360
rect 14415 19329 14427 19332
rect 14461 19360 14473 19363
rect 23474 19360 23480 19372
rect 14461 19332 23480 19360
rect 14461 19329 14473 19332
rect 14415 19323 14473 19329
rect 23474 19320 23480 19332
rect 23532 19320 23538 19372
rect 14550 19292 14556 19304
rect 12912 19264 14556 19292
rect 14550 19252 14556 19264
rect 14608 19252 14614 19304
rect 1104 19066 28888 19088
rect 1104 19014 2918 19066
rect 2970 19014 2982 19066
rect 3034 19014 3046 19066
rect 3098 19014 3110 19066
rect 3162 19014 3174 19066
rect 3226 19014 3238 19066
rect 3290 19014 10918 19066
rect 10970 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 11238 19066
rect 11290 19014 18918 19066
rect 18970 19014 18982 19066
rect 19034 19014 19046 19066
rect 19098 19014 19110 19066
rect 19162 19014 19174 19066
rect 19226 19014 19238 19066
rect 19290 19014 26918 19066
rect 26970 19014 26982 19066
rect 27034 19014 27046 19066
rect 27098 19014 27110 19066
rect 27162 19014 27174 19066
rect 27226 19014 27238 19066
rect 27290 19014 28888 19066
rect 1104 18992 28888 19014
rect 13814 18776 13820 18828
rect 13872 18816 13878 18828
rect 14642 18816 14648 18828
rect 13872 18788 14648 18816
rect 13872 18776 13878 18788
rect 14642 18776 14648 18788
rect 14700 18776 14706 18828
rect 14550 18708 14556 18760
rect 14608 18708 14614 18760
rect 23474 18708 23480 18760
rect 23532 18748 23538 18760
rect 28077 18751 28135 18757
rect 28077 18748 28089 18751
rect 23532 18720 28089 18748
rect 23532 18708 23538 18720
rect 28077 18717 28089 18720
rect 28123 18717 28135 18751
rect 28077 18711 28135 18717
rect 12253 18683 12311 18689
rect 12253 18649 12265 18683
rect 12299 18680 12311 18683
rect 12342 18680 12348 18692
rect 12299 18652 12348 18680
rect 12299 18649 12311 18652
rect 12253 18643 12311 18649
rect 12342 18640 12348 18652
rect 12400 18640 12406 18692
rect 28350 18640 28356 18692
rect 28408 18640 28414 18692
rect 12710 18572 12716 18624
rect 12768 18612 12774 18624
rect 14093 18615 14151 18621
rect 14093 18612 14105 18615
rect 12768 18584 14105 18612
rect 12768 18572 12774 18584
rect 14093 18581 14105 18584
rect 14139 18581 14151 18615
rect 14093 18575 14151 18581
rect 14458 18572 14464 18624
rect 14516 18572 14522 18624
rect 1104 18522 28888 18544
rect 1104 18470 3658 18522
rect 3710 18470 3722 18522
rect 3774 18470 3786 18522
rect 3838 18470 3850 18522
rect 3902 18470 3914 18522
rect 3966 18470 3978 18522
rect 4030 18470 11658 18522
rect 11710 18470 11722 18522
rect 11774 18470 11786 18522
rect 11838 18470 11850 18522
rect 11902 18470 11914 18522
rect 11966 18470 11978 18522
rect 12030 18470 19658 18522
rect 19710 18470 19722 18522
rect 19774 18470 19786 18522
rect 19838 18470 19850 18522
rect 19902 18470 19914 18522
rect 19966 18470 19978 18522
rect 20030 18470 27658 18522
rect 27710 18470 27722 18522
rect 27774 18470 27786 18522
rect 27838 18470 27850 18522
rect 27902 18470 27914 18522
rect 27966 18470 27978 18522
rect 28030 18470 28888 18522
rect 1104 18448 28888 18470
rect 1581 18411 1639 18417
rect 1581 18377 1593 18411
rect 1627 18408 1639 18411
rect 14550 18408 14556 18420
rect 1627 18380 14556 18408
rect 1627 18377 1639 18380
rect 1581 18371 1639 18377
rect 14550 18368 14556 18380
rect 14608 18368 14614 18420
rect 13722 18300 13728 18352
rect 13780 18300 13786 18352
rect 1394 18232 1400 18284
rect 1452 18232 1458 18284
rect 12710 18232 12716 18284
rect 12768 18232 12774 18284
rect 14139 18275 14197 18281
rect 14139 18241 14151 18275
rect 14185 18272 14197 18275
rect 14458 18272 14464 18284
rect 14185 18244 14464 18272
rect 14185 18241 14197 18244
rect 14139 18235 14197 18241
rect 14458 18232 14464 18244
rect 14516 18272 14522 18284
rect 28077 18275 28135 18281
rect 28077 18272 28089 18275
rect 14516 18244 28089 18272
rect 14516 18232 14522 18244
rect 28077 18241 28089 18244
rect 28123 18241 28135 18275
rect 28077 18235 28135 18241
rect 12342 18164 12348 18216
rect 12400 18164 12406 18216
rect 28350 18164 28356 18216
rect 28408 18164 28414 18216
rect 1104 17978 28888 18000
rect 1104 17926 2918 17978
rect 2970 17926 2982 17978
rect 3034 17926 3046 17978
rect 3098 17926 3110 17978
rect 3162 17926 3174 17978
rect 3226 17926 3238 17978
rect 3290 17926 10918 17978
rect 10970 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 11238 17978
rect 11290 17926 18918 17978
rect 18970 17926 18982 17978
rect 19034 17926 19046 17978
rect 19098 17926 19110 17978
rect 19162 17926 19174 17978
rect 19226 17926 19238 17978
rect 19290 17926 26918 17978
rect 26970 17926 26982 17978
rect 27034 17926 27046 17978
rect 27098 17926 27110 17978
rect 27162 17926 27174 17978
rect 27226 17926 27238 17978
rect 27290 17926 28888 17978
rect 1104 17904 28888 17926
rect 12342 17824 12348 17876
rect 12400 17864 12406 17876
rect 13449 17867 13507 17873
rect 13449 17864 13461 17867
rect 12400 17836 13461 17864
rect 12400 17824 12406 17836
rect 13449 17833 13461 17836
rect 13495 17833 13507 17867
rect 13449 17827 13507 17833
rect 14550 17688 14556 17740
rect 14608 17688 14614 17740
rect 14642 17688 14648 17740
rect 14700 17688 14706 17740
rect 1394 17620 1400 17672
rect 1452 17620 1458 17672
rect 11514 17620 11520 17672
rect 11572 17660 11578 17672
rect 12158 17660 12164 17672
rect 11572 17632 12164 17660
rect 11572 17620 11578 17632
rect 12158 17620 12164 17632
rect 12216 17620 12222 17672
rect 1581 17527 1639 17533
rect 1581 17493 1593 17527
rect 1627 17524 1639 17527
rect 11330 17524 11336 17536
rect 1627 17496 11336 17524
rect 1627 17493 1639 17496
rect 1581 17487 1639 17493
rect 11330 17484 11336 17496
rect 11388 17484 11394 17536
rect 12434 17484 12440 17536
rect 12492 17524 12498 17536
rect 14093 17527 14151 17533
rect 14093 17524 14105 17527
rect 12492 17496 14105 17524
rect 12492 17484 12498 17496
rect 14093 17493 14105 17496
rect 14139 17493 14151 17527
rect 14093 17487 14151 17493
rect 14458 17484 14464 17536
rect 14516 17484 14522 17536
rect 1104 17434 28888 17456
rect 1104 17382 3658 17434
rect 3710 17382 3722 17434
rect 3774 17382 3786 17434
rect 3838 17382 3850 17434
rect 3902 17382 3914 17434
rect 3966 17382 3978 17434
rect 4030 17382 11658 17434
rect 11710 17382 11722 17434
rect 11774 17382 11786 17434
rect 11838 17382 11850 17434
rect 11902 17382 11914 17434
rect 11966 17382 11978 17434
rect 12030 17382 19658 17434
rect 19710 17382 19722 17434
rect 19774 17382 19786 17434
rect 19838 17382 19850 17434
rect 19902 17382 19914 17434
rect 19966 17382 19978 17434
rect 20030 17382 27658 17434
rect 27710 17382 27722 17434
rect 27774 17382 27786 17434
rect 27838 17382 27850 17434
rect 27902 17382 27914 17434
rect 27966 17382 27978 17434
rect 28030 17382 28888 17434
rect 1104 17360 28888 17382
rect 13722 17252 13728 17264
rect 13478 17238 13728 17252
rect 13464 17224 13728 17238
rect 12434 17144 12440 17196
rect 12492 17144 12498 17196
rect 11514 17076 11520 17128
rect 11572 17116 11578 17128
rect 12069 17119 12127 17125
rect 12069 17116 12081 17119
rect 11572 17088 12081 17116
rect 11572 17076 11578 17088
rect 12069 17085 12081 17088
rect 12115 17116 12127 17119
rect 12342 17116 12348 17128
rect 12115 17088 12348 17116
rect 12115 17085 12127 17088
rect 12069 17079 12127 17085
rect 12342 17076 12348 17088
rect 12400 17076 12406 17128
rect 12986 17076 12992 17128
rect 13044 17116 13050 17128
rect 13464 17116 13492 17224
rect 13722 17212 13728 17224
rect 13780 17212 13786 17264
rect 13863 17187 13921 17193
rect 13863 17153 13875 17187
rect 13909 17184 13921 17187
rect 14458 17184 14464 17196
rect 13909 17156 14464 17184
rect 13909 17153 13921 17156
rect 13863 17147 13921 17153
rect 14458 17144 14464 17156
rect 14516 17184 14522 17196
rect 28077 17187 28135 17193
rect 28077 17184 28089 17187
rect 14516 17156 28089 17184
rect 14516 17144 14522 17156
rect 28077 17153 28089 17156
rect 28123 17153 28135 17187
rect 28077 17147 28135 17153
rect 13044 17088 13492 17116
rect 13044 17076 13050 17088
rect 28350 17076 28356 17128
rect 28408 17076 28414 17128
rect 1104 16890 28888 16912
rect 1104 16838 2918 16890
rect 2970 16838 2982 16890
rect 3034 16838 3046 16890
rect 3098 16838 3110 16890
rect 3162 16838 3174 16890
rect 3226 16838 3238 16890
rect 3290 16838 10918 16890
rect 10970 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 11238 16890
rect 11290 16838 18918 16890
rect 18970 16838 18982 16890
rect 19034 16838 19046 16890
rect 19098 16838 19110 16890
rect 19162 16838 19174 16890
rect 19226 16838 19238 16890
rect 19290 16838 26918 16890
rect 26970 16838 26982 16890
rect 27034 16838 27046 16890
rect 27098 16838 27110 16890
rect 27162 16838 27174 16890
rect 27226 16838 27238 16890
rect 27290 16838 28888 16890
rect 1104 16816 28888 16838
rect 1394 16532 1400 16584
rect 1452 16532 1458 16584
rect 11514 16532 11520 16584
rect 11572 16572 11578 16584
rect 11609 16575 11667 16581
rect 11609 16572 11621 16575
rect 11572 16544 11621 16572
rect 11572 16532 11578 16544
rect 11609 16541 11621 16544
rect 11655 16541 11667 16575
rect 11609 16535 11667 16541
rect 11977 16575 12035 16581
rect 11977 16541 11989 16575
rect 12023 16572 12035 16575
rect 12066 16572 12072 16584
rect 12023 16544 12072 16572
rect 12023 16541 12035 16544
rect 11977 16535 12035 16541
rect 12066 16532 12072 16544
rect 12124 16532 12130 16584
rect 21358 16532 21364 16584
rect 21416 16572 21422 16584
rect 28077 16575 28135 16581
rect 28077 16572 28089 16575
rect 21416 16544 28089 16572
rect 21416 16532 21422 16544
rect 28077 16541 28089 16544
rect 28123 16541 28135 16575
rect 28077 16535 28135 16541
rect 12268 16476 12374 16504
rect 1581 16439 1639 16445
rect 1581 16405 1593 16439
rect 1627 16436 1639 16439
rect 10870 16436 10876 16448
rect 1627 16408 10876 16436
rect 1627 16405 1639 16408
rect 1581 16399 1639 16405
rect 10870 16396 10876 16408
rect 10928 16396 10934 16448
rect 12268 16436 12296 16476
rect 28350 16464 28356 16516
rect 28408 16464 28414 16516
rect 12434 16436 12440 16448
rect 12268 16408 12440 16436
rect 12434 16396 12440 16408
rect 12492 16436 12498 16448
rect 12894 16436 12900 16448
rect 12492 16408 12900 16436
rect 12492 16396 12498 16408
rect 12894 16396 12900 16408
rect 12952 16396 12958 16448
rect 13446 16445 13452 16448
rect 13403 16439 13452 16445
rect 13403 16405 13415 16439
rect 13449 16405 13452 16439
rect 13403 16399 13452 16405
rect 13446 16396 13452 16399
rect 13504 16396 13510 16448
rect 1104 16346 28888 16368
rect 1104 16294 3658 16346
rect 3710 16294 3722 16346
rect 3774 16294 3786 16346
rect 3838 16294 3850 16346
rect 3902 16294 3914 16346
rect 3966 16294 3978 16346
rect 4030 16294 11658 16346
rect 11710 16294 11722 16346
rect 11774 16294 11786 16346
rect 11838 16294 11850 16346
rect 11902 16294 11914 16346
rect 11966 16294 11978 16346
rect 12030 16294 19658 16346
rect 19710 16294 19722 16346
rect 19774 16294 19786 16346
rect 19838 16294 19850 16346
rect 19902 16294 19914 16346
rect 19966 16294 19978 16346
rect 20030 16294 27658 16346
rect 27710 16294 27722 16346
rect 27774 16294 27786 16346
rect 27838 16294 27850 16346
rect 27902 16294 27914 16346
rect 27966 16294 27978 16346
rect 28030 16294 28888 16346
rect 1104 16272 28888 16294
rect 10870 16192 10876 16244
rect 10928 16192 10934 16244
rect 12434 16124 12440 16176
rect 12492 16124 12498 16176
rect 1394 16056 1400 16108
rect 1452 16056 1458 16108
rect 10965 16099 11023 16105
rect 10965 16065 10977 16099
rect 11011 16096 11023 16099
rect 11011 16068 11284 16096
rect 11011 16065 11023 16068
rect 10965 16059 11023 16065
rect 10686 15988 10692 16040
rect 10744 15988 10750 16040
rect 1581 15895 1639 15901
rect 1581 15861 1593 15895
rect 1627 15892 1639 15895
rect 10778 15892 10784 15904
rect 1627 15864 10784 15892
rect 1627 15861 1639 15864
rect 1581 15855 1639 15861
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 11256 15892 11284 16068
rect 11514 16056 11520 16108
rect 11572 16056 11578 16108
rect 11885 16031 11943 16037
rect 11885 16028 11897 16031
rect 11348 16000 11897 16028
rect 11348 15969 11376 16000
rect 11885 15997 11897 16000
rect 11931 15997 11943 16031
rect 11885 15991 11943 15997
rect 11333 15963 11391 15969
rect 11333 15929 11345 15963
rect 11379 15929 11391 15963
rect 11333 15923 11391 15929
rect 13311 15895 13369 15901
rect 13311 15892 13323 15895
rect 11256 15864 13323 15892
rect 13311 15861 13323 15864
rect 13357 15892 13369 15895
rect 28074 15892 28080 15904
rect 13357 15864 28080 15892
rect 13357 15861 13369 15864
rect 13311 15855 13369 15861
rect 28074 15852 28080 15864
rect 28132 15852 28138 15904
rect 1104 15802 28888 15824
rect 1104 15750 2918 15802
rect 2970 15750 2982 15802
rect 3034 15750 3046 15802
rect 3098 15750 3110 15802
rect 3162 15750 3174 15802
rect 3226 15750 3238 15802
rect 3290 15750 10918 15802
rect 10970 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 11238 15802
rect 11290 15750 18918 15802
rect 18970 15750 18982 15802
rect 19034 15750 19046 15802
rect 19098 15750 19110 15802
rect 19162 15750 19174 15802
rect 19226 15750 19238 15802
rect 19290 15750 26918 15802
rect 26970 15750 26982 15802
rect 27034 15750 27046 15802
rect 27098 15750 27110 15802
rect 27162 15750 27174 15802
rect 27226 15750 27238 15802
rect 27290 15750 28888 15802
rect 1104 15728 28888 15750
rect 11422 15648 11428 15700
rect 11480 15688 11486 15700
rect 11701 15691 11759 15697
rect 11701 15688 11713 15691
rect 11480 15660 11713 15688
rect 11480 15648 11486 15660
rect 11701 15657 11713 15660
rect 11747 15657 11759 15691
rect 11701 15651 11759 15657
rect 12066 15648 12072 15700
rect 12124 15648 12130 15700
rect 10686 15580 10692 15632
rect 10744 15620 10750 15632
rect 10781 15623 10839 15629
rect 10781 15620 10793 15623
rect 10744 15592 10793 15620
rect 10744 15580 10750 15592
rect 10781 15589 10793 15592
rect 10827 15620 10839 15623
rect 10827 15592 12756 15620
rect 10827 15589 10839 15592
rect 10781 15583 10839 15589
rect 11330 15512 11336 15564
rect 11388 15552 11394 15564
rect 12728 15561 12756 15592
rect 12529 15555 12587 15561
rect 12529 15552 12541 15555
rect 11388 15524 12541 15552
rect 11388 15512 11394 15524
rect 12529 15521 12541 15524
rect 12575 15521 12587 15555
rect 12529 15515 12587 15521
rect 12713 15555 12771 15561
rect 12713 15521 12725 15555
rect 12759 15552 12771 15555
rect 14642 15552 14648 15564
rect 12759 15524 14648 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 14642 15512 14648 15524
rect 14700 15512 14706 15564
rect 10965 15487 11023 15493
rect 10965 15453 10977 15487
rect 11011 15484 11023 15487
rect 11422 15484 11428 15496
rect 11011 15456 11428 15484
rect 11011 15453 11023 15456
rect 10965 15447 11023 15453
rect 11422 15444 11428 15456
rect 11480 15444 11486 15496
rect 12250 15484 12256 15496
rect 11532 15456 12256 15484
rect 11241 15419 11299 15425
rect 11241 15385 11253 15419
rect 11287 15416 11299 15419
rect 11532 15416 11560 15456
rect 12250 15444 12256 15456
rect 12308 15444 12314 15496
rect 28074 15444 28080 15496
rect 28132 15444 28138 15496
rect 11287 15388 11560 15416
rect 11287 15385 11299 15388
rect 11241 15379 11299 15385
rect 11606 15376 11612 15428
rect 11664 15376 11670 15428
rect 12437 15419 12495 15425
rect 12437 15385 12449 15419
rect 12483 15416 12495 15419
rect 13446 15416 13452 15428
rect 12483 15388 13452 15416
rect 12483 15385 12495 15388
rect 12437 15379 12495 15385
rect 13446 15376 13452 15388
rect 13504 15416 13510 15428
rect 21358 15416 21364 15428
rect 13504 15388 21364 15416
rect 13504 15376 13510 15388
rect 21358 15376 21364 15388
rect 21416 15376 21422 15428
rect 28350 15376 28356 15428
rect 28408 15376 28414 15428
rect 11333 15351 11391 15357
rect 11333 15317 11345 15351
rect 11379 15348 11391 15351
rect 12618 15348 12624 15360
rect 11379 15320 12624 15348
rect 11379 15317 11391 15320
rect 11333 15311 11391 15317
rect 12618 15308 12624 15320
rect 12676 15308 12682 15360
rect 1104 15258 28888 15280
rect 1104 15206 3658 15258
rect 3710 15206 3722 15258
rect 3774 15206 3786 15258
rect 3838 15206 3850 15258
rect 3902 15206 3914 15258
rect 3966 15206 3978 15258
rect 4030 15206 11658 15258
rect 11710 15206 11722 15258
rect 11774 15206 11786 15258
rect 11838 15206 11850 15258
rect 11902 15206 11914 15258
rect 11966 15206 11978 15258
rect 12030 15206 19658 15258
rect 19710 15206 19722 15258
rect 19774 15206 19786 15258
rect 19838 15206 19850 15258
rect 19902 15206 19914 15258
rect 19966 15206 19978 15258
rect 20030 15206 27658 15258
rect 27710 15206 27722 15258
rect 27774 15206 27786 15258
rect 27838 15206 27850 15258
rect 27902 15206 27914 15258
rect 27966 15206 27978 15258
rect 28030 15206 28888 15258
rect 1104 15184 28888 15206
rect 10778 15104 10784 15156
rect 10836 15144 10842 15156
rect 11057 15147 11115 15153
rect 11057 15144 11069 15147
rect 10836 15116 11069 15144
rect 10836 15104 10842 15116
rect 11057 15113 11069 15116
rect 11103 15113 11115 15147
rect 11057 15107 11115 15113
rect 11517 15079 11575 15085
rect 11517 15076 11529 15079
rect 6886 15048 11529 15076
rect 1394 14968 1400 15020
rect 1452 14968 1458 15020
rect 106 14900 112 14952
rect 164 14940 170 14952
rect 6886 14940 6914 15048
rect 11517 15045 11529 15048
rect 11563 15045 11575 15079
rect 11517 15039 11575 15045
rect 10965 15011 11023 15017
rect 10965 14977 10977 15011
rect 11011 15008 11023 15011
rect 11790 15008 11796 15020
rect 11011 14980 11796 15008
rect 11011 14977 11023 14980
rect 10965 14971 11023 14977
rect 11790 14968 11796 14980
rect 11848 14968 11854 15020
rect 28074 14968 28080 15020
rect 28132 14968 28138 15020
rect 164 14912 6914 14940
rect 164 14900 170 14912
rect 10686 14900 10692 14952
rect 10744 14940 10750 14952
rect 11149 14943 11207 14949
rect 11149 14940 11161 14943
rect 10744 14912 11161 14940
rect 10744 14900 10750 14912
rect 11149 14909 11161 14912
rect 11195 14909 11207 14943
rect 11149 14903 11207 14909
rect 28350 14900 28356 14952
rect 28408 14900 28414 14952
rect 1581 14875 1639 14881
rect 1581 14841 1593 14875
rect 1627 14872 1639 14875
rect 11514 14872 11520 14884
rect 1627 14844 11520 14872
rect 1627 14841 1639 14844
rect 1581 14835 1639 14841
rect 11514 14832 11520 14844
rect 11572 14832 11578 14884
rect 10597 14807 10655 14813
rect 10597 14773 10609 14807
rect 10643 14804 10655 14807
rect 10778 14804 10784 14816
rect 10643 14776 10784 14804
rect 10643 14773 10655 14776
rect 10597 14767 10655 14773
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 12158 14764 12164 14816
rect 12216 14804 12222 14816
rect 12802 14804 12808 14816
rect 12216 14776 12808 14804
rect 12216 14764 12222 14776
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 1104 14714 28888 14736
rect 1104 14662 2918 14714
rect 2970 14662 2982 14714
rect 3034 14662 3046 14714
rect 3098 14662 3110 14714
rect 3162 14662 3174 14714
rect 3226 14662 3238 14714
rect 3290 14662 10918 14714
rect 10970 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 11238 14714
rect 11290 14662 18918 14714
rect 18970 14662 18982 14714
rect 19034 14662 19046 14714
rect 19098 14662 19110 14714
rect 19162 14662 19174 14714
rect 19226 14662 19238 14714
rect 19290 14662 26918 14714
rect 26970 14662 26982 14714
rect 27034 14662 27046 14714
rect 27098 14662 27110 14714
rect 27162 14662 27174 14714
rect 27226 14662 27238 14714
rect 27290 14662 28888 14714
rect 1104 14640 28888 14662
rect 10778 14424 10784 14476
rect 10836 14464 10842 14476
rect 10965 14467 11023 14473
rect 10965 14464 10977 14467
rect 10836 14436 10977 14464
rect 10836 14424 10842 14436
rect 10965 14433 10977 14436
rect 11011 14433 11023 14467
rect 10965 14427 11023 14433
rect 1394 14356 1400 14408
rect 1452 14356 1458 14408
rect 10597 14399 10655 14405
rect 10597 14365 10609 14399
rect 10643 14396 10655 14399
rect 10686 14396 10692 14408
rect 10643 14368 10692 14396
rect 10643 14365 10655 14368
rect 10597 14359 10655 14365
rect 10686 14356 10692 14368
rect 10744 14356 10750 14408
rect 11790 14356 11796 14408
rect 11848 14396 11854 14408
rect 12391 14399 12449 14405
rect 12391 14396 12403 14399
rect 11848 14368 12403 14396
rect 11848 14356 11854 14368
rect 12391 14365 12403 14368
rect 12437 14396 12449 14399
rect 12437 14368 16574 14396
rect 12437 14365 12449 14368
rect 12391 14359 12449 14365
rect 12529 14331 12587 14337
rect 12529 14328 12541 14331
rect 12006 14300 12541 14328
rect 12452 14272 12480 14300
rect 12529 14297 12541 14300
rect 12575 14297 12587 14331
rect 12529 14291 12587 14297
rect 12710 14288 12716 14340
rect 12768 14288 12774 14340
rect 1581 14263 1639 14269
rect 1581 14229 1593 14263
rect 1627 14260 1639 14263
rect 12158 14260 12164 14272
rect 1627 14232 12164 14260
rect 1627 14229 1639 14232
rect 1581 14223 1639 14229
rect 12158 14220 12164 14232
rect 12216 14220 12222 14272
rect 12434 14220 12440 14272
rect 12492 14220 12498 14272
rect 16546 14260 16574 14368
rect 28074 14260 28080 14272
rect 16546 14232 28080 14260
rect 28074 14220 28080 14232
rect 28132 14220 28138 14272
rect 1104 14170 28888 14192
rect 1104 14118 3658 14170
rect 3710 14118 3722 14170
rect 3774 14118 3786 14170
rect 3838 14118 3850 14170
rect 3902 14118 3914 14170
rect 3966 14118 3978 14170
rect 4030 14118 11658 14170
rect 11710 14118 11722 14170
rect 11774 14118 11786 14170
rect 11838 14118 11850 14170
rect 11902 14118 11914 14170
rect 11966 14118 11978 14170
rect 12030 14118 19658 14170
rect 19710 14118 19722 14170
rect 19774 14118 19786 14170
rect 19838 14118 19850 14170
rect 19902 14118 19914 14170
rect 19966 14118 19978 14170
rect 20030 14118 27658 14170
rect 27710 14118 27722 14170
rect 27774 14118 27786 14170
rect 27838 14118 27850 14170
rect 27902 14118 27914 14170
rect 27966 14118 27978 14170
rect 28030 14118 28888 14170
rect 1104 14096 28888 14118
rect 11514 14016 11520 14068
rect 11572 14056 11578 14068
rect 11977 14059 12035 14065
rect 11977 14056 11989 14059
rect 11572 14028 11989 14056
rect 11572 14016 11578 14028
rect 11977 14025 11989 14028
rect 12023 14025 12035 14059
rect 11977 14019 12035 14025
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 12342 13920 12348 13932
rect 11931 13892 12348 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 12342 13880 12348 13892
rect 12400 13920 12406 13932
rect 28077 13923 28135 13929
rect 28077 13920 28089 13923
rect 12400 13892 28089 13920
rect 12400 13880 12406 13892
rect 28077 13889 28089 13892
rect 28123 13889 28135 13923
rect 28077 13883 28135 13889
rect 10318 13812 10324 13864
rect 10376 13852 10382 13864
rect 12069 13855 12127 13861
rect 12069 13852 12081 13855
rect 10376 13824 12081 13852
rect 10376 13812 10382 13824
rect 12069 13821 12081 13824
rect 12115 13821 12127 13855
rect 12069 13815 12127 13821
rect 28350 13812 28356 13864
rect 28408 13812 28414 13864
rect 11514 13676 11520 13728
rect 11572 13676 11578 13728
rect 1104 13626 28888 13648
rect 1104 13574 2918 13626
rect 2970 13574 2982 13626
rect 3034 13574 3046 13626
rect 3098 13574 3110 13626
rect 3162 13574 3174 13626
rect 3226 13574 3238 13626
rect 3290 13574 10918 13626
rect 10970 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 11238 13626
rect 11290 13574 18918 13626
rect 18970 13574 18982 13626
rect 19034 13574 19046 13626
rect 19098 13574 19110 13626
rect 19162 13574 19174 13626
rect 19226 13574 19238 13626
rect 19290 13574 26918 13626
rect 26970 13574 26982 13626
rect 27034 13574 27046 13626
rect 27098 13574 27110 13626
rect 27162 13574 27174 13626
rect 27226 13574 27238 13626
rect 27290 13574 28888 13626
rect 1104 13552 28888 13574
rect 10778 13472 10784 13524
rect 10836 13512 10842 13524
rect 10836 13484 11744 13512
rect 10836 13472 10842 13484
rect 11716 13444 11744 13484
rect 12342 13472 12348 13524
rect 12400 13521 12406 13524
rect 12400 13515 12449 13521
rect 12400 13481 12403 13515
rect 12437 13481 12449 13515
rect 12400 13475 12449 13481
rect 12400 13472 12406 13475
rect 11716 13416 13124 13444
rect 10965 13379 11023 13385
rect 10965 13345 10977 13379
rect 11011 13376 11023 13379
rect 11514 13376 11520 13388
rect 11011 13348 11520 13376
rect 11011 13345 11023 13348
rect 10965 13339 11023 13345
rect 11514 13336 11520 13348
rect 11572 13336 11578 13388
rect 12158 13336 12164 13388
rect 12216 13376 12222 13388
rect 13096 13385 13124 13416
rect 12989 13379 13047 13385
rect 12989 13376 13001 13379
rect 12216 13348 13001 13376
rect 12216 13336 12222 13348
rect 12989 13345 13001 13348
rect 13035 13345 13047 13379
rect 12989 13339 13047 13345
rect 13081 13379 13139 13385
rect 13081 13345 13093 13379
rect 13127 13345 13139 13379
rect 13081 13339 13139 13345
rect 1394 13268 1400 13320
rect 1452 13268 1458 13320
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13308 10655 13311
rect 10686 13308 10692 13320
rect 10643 13280 10692 13308
rect 10643 13277 10655 13280
rect 10597 13271 10655 13277
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 12897 13311 12955 13317
rect 12897 13277 12909 13311
rect 12943 13308 12955 13311
rect 13354 13308 13360 13320
rect 12943 13280 13360 13308
rect 12943 13277 12955 13280
rect 12897 13271 12955 13277
rect 13354 13268 13360 13280
rect 13412 13308 13418 13320
rect 28077 13311 28135 13317
rect 28077 13308 28089 13311
rect 13412 13280 28089 13308
rect 13412 13268 13418 13280
rect 28077 13277 28089 13280
rect 28123 13277 28135 13311
rect 28077 13271 28135 13277
rect 12342 13240 12348 13252
rect 12006 13212 12348 13240
rect 12342 13200 12348 13212
rect 12400 13200 12406 13252
rect 28350 13200 28356 13252
rect 28408 13200 28414 13252
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 10870 13172 10876 13184
rect 1627 13144 10876 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 12529 13175 12587 13181
rect 12529 13141 12541 13175
rect 12575 13172 12587 13175
rect 12618 13172 12624 13184
rect 12575 13144 12624 13172
rect 12575 13141 12587 13144
rect 12529 13135 12587 13141
rect 12618 13132 12624 13144
rect 12676 13132 12682 13184
rect 1104 13082 28888 13104
rect 1104 13030 3658 13082
rect 3710 13030 3722 13082
rect 3774 13030 3786 13082
rect 3838 13030 3850 13082
rect 3902 13030 3914 13082
rect 3966 13030 3978 13082
rect 4030 13030 11658 13082
rect 11710 13030 11722 13082
rect 11774 13030 11786 13082
rect 11838 13030 11850 13082
rect 11902 13030 11914 13082
rect 11966 13030 11978 13082
rect 12030 13030 19658 13082
rect 19710 13030 19722 13082
rect 19774 13030 19786 13082
rect 19838 13030 19850 13082
rect 19902 13030 19914 13082
rect 19966 13030 19978 13082
rect 20030 13030 27658 13082
rect 27710 13030 27722 13082
rect 27774 13030 27786 13082
rect 27838 13030 27850 13082
rect 27902 13030 27914 13082
rect 27966 13030 27978 13082
rect 28030 13030 28888 13082
rect 1104 13008 28888 13030
rect 10870 12928 10876 12980
rect 10928 12928 10934 12980
rect 13354 12977 13360 12980
rect 13311 12971 13360 12977
rect 13311 12937 13323 12971
rect 13357 12937 13360 12971
rect 13311 12931 13360 12937
rect 13354 12928 13360 12931
rect 13412 12928 13418 12980
rect 12434 12860 12440 12912
rect 12492 12860 12498 12912
rect 1394 12792 1400 12844
rect 1452 12792 1458 12844
rect 10965 12835 11023 12841
rect 10965 12801 10977 12835
rect 11011 12832 11023 12835
rect 11974 12832 11980 12844
rect 11011 12804 11980 12832
rect 11011 12801 11023 12804
rect 10965 12795 11023 12801
rect 11974 12792 11980 12804
rect 12032 12792 12038 12844
rect 10778 12724 10784 12776
rect 10836 12724 10842 12776
rect 11517 12767 11575 12773
rect 11517 12733 11529 12767
rect 11563 12733 11575 12767
rect 11517 12727 11575 12733
rect 11885 12767 11943 12773
rect 11885 12733 11897 12767
rect 11931 12764 11943 12767
rect 12618 12764 12624 12776
rect 11931 12736 12624 12764
rect 11931 12733 11943 12736
rect 11885 12727 11943 12733
rect 11532 12696 11560 12727
rect 12618 12724 12624 12736
rect 12676 12724 12682 12776
rect 10704 12668 11560 12696
rect 10704 12640 10732 12668
rect 1581 12631 1639 12637
rect 1581 12597 1593 12631
rect 1627 12628 1639 12631
rect 10594 12628 10600 12640
rect 1627 12600 10600 12628
rect 1627 12597 1639 12600
rect 1581 12591 1639 12597
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 10686 12588 10692 12640
rect 10744 12588 10750 12640
rect 11330 12588 11336 12640
rect 11388 12588 11394 12640
rect 1104 12538 28888 12560
rect 1104 12486 2918 12538
rect 2970 12486 2982 12538
rect 3034 12486 3046 12538
rect 3098 12486 3110 12538
rect 3162 12486 3174 12538
rect 3226 12486 3238 12538
rect 3290 12486 10918 12538
rect 10970 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 11238 12538
rect 11290 12486 18918 12538
rect 18970 12486 18982 12538
rect 19034 12486 19046 12538
rect 19098 12486 19110 12538
rect 19162 12486 19174 12538
rect 19226 12486 19238 12538
rect 19290 12486 26918 12538
rect 26970 12486 26982 12538
rect 27034 12486 27046 12538
rect 27098 12486 27110 12538
rect 27162 12486 27174 12538
rect 27226 12486 27238 12538
rect 27290 12486 28888 12538
rect 1104 12464 28888 12486
rect 11057 12291 11115 12297
rect 11057 12257 11069 12291
rect 11103 12288 11115 12291
rect 11330 12288 11336 12300
rect 11103 12260 11336 12288
rect 11103 12257 11115 12260
rect 11057 12251 11115 12257
rect 11330 12248 11336 12260
rect 11388 12248 11394 12300
rect 10505 12223 10563 12229
rect 10505 12189 10517 12223
rect 10551 12220 10563 12223
rect 10686 12220 10692 12232
rect 10551 12192 10692 12220
rect 10551 12189 10563 12192
rect 10505 12183 10563 12189
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 11974 12180 11980 12232
rect 12032 12220 12038 12232
rect 12483 12223 12541 12229
rect 12483 12220 12495 12223
rect 12032 12192 12495 12220
rect 12032 12180 12038 12192
rect 12483 12189 12495 12192
rect 12529 12220 12541 12223
rect 28077 12223 28135 12229
rect 28077 12220 28089 12223
rect 12529 12192 28089 12220
rect 12529 12189 12541 12192
rect 12483 12183 12541 12189
rect 28077 12189 28089 12192
rect 28123 12189 28135 12223
rect 28077 12183 28135 12189
rect 12342 12152 12348 12164
rect 12098 12124 12348 12152
rect 12342 12112 12348 12124
rect 12400 12112 12406 12164
rect 28350 12112 28356 12164
rect 28408 12112 28414 12164
rect 1104 11994 28888 12016
rect 1104 11942 3658 11994
rect 3710 11942 3722 11994
rect 3774 11942 3786 11994
rect 3838 11942 3850 11994
rect 3902 11942 3914 11994
rect 3966 11942 3978 11994
rect 4030 11942 11658 11994
rect 11710 11942 11722 11994
rect 11774 11942 11786 11994
rect 11838 11942 11850 11994
rect 11902 11942 11914 11994
rect 11966 11942 11978 11994
rect 12030 11942 19658 11994
rect 19710 11942 19722 11994
rect 19774 11942 19786 11994
rect 19838 11942 19850 11994
rect 19902 11942 19914 11994
rect 19966 11942 19978 11994
rect 20030 11942 27658 11994
rect 27710 11942 27722 11994
rect 27774 11942 27786 11994
rect 27838 11942 27850 11994
rect 27902 11942 27914 11994
rect 27966 11942 27978 11994
rect 28030 11942 28888 11994
rect 1104 11920 28888 11942
rect 12434 11772 12440 11824
rect 12492 11772 12498 11824
rect 1394 11704 1400 11756
rect 1452 11704 1458 11756
rect 11333 11747 11391 11753
rect 11333 11713 11345 11747
rect 11379 11744 11391 11747
rect 13311 11747 13369 11753
rect 13311 11744 13323 11747
rect 11379 11716 12020 11744
rect 11379 11713 11391 11716
rect 11333 11707 11391 11713
rect 10686 11676 10692 11688
rect 10060 11648 10692 11676
rect 10060 11617 10088 11648
rect 10686 11636 10692 11648
rect 10744 11676 10750 11688
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 10744 11648 11529 11676
rect 10744 11636 10750 11648
rect 11517 11645 11529 11648
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 11698 11636 11704 11688
rect 11756 11676 11762 11688
rect 11885 11679 11943 11685
rect 11885 11676 11897 11679
rect 11756 11648 11897 11676
rect 11756 11636 11762 11648
rect 11885 11645 11897 11648
rect 11931 11645 11943 11679
rect 11992 11676 12020 11716
rect 12912 11716 13323 11744
rect 12802 11676 12808 11688
rect 11992 11648 12808 11676
rect 11885 11639 11943 11645
rect 12802 11636 12808 11648
rect 12860 11636 12866 11688
rect 10045 11611 10103 11617
rect 10045 11577 10057 11611
rect 10091 11577 10103 11611
rect 11422 11608 11428 11620
rect 10045 11571 10103 11577
rect 11256 11580 11428 11608
rect 1581 11543 1639 11549
rect 1581 11509 1593 11543
rect 1627 11540 1639 11543
rect 11256 11540 11284 11580
rect 11422 11568 11428 11580
rect 11480 11568 11486 11620
rect 1627 11512 11284 11540
rect 1627 11509 1639 11512
rect 1581 11503 1639 11509
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 12912 11540 12940 11716
rect 13311 11713 13323 11716
rect 13357 11744 13369 11747
rect 28077 11747 28135 11753
rect 28077 11744 28089 11747
rect 13357 11716 28089 11744
rect 13357 11713 13369 11716
rect 13311 11707 13369 11713
rect 28077 11713 28089 11716
rect 28123 11713 28135 11747
rect 28077 11707 28135 11713
rect 28350 11636 28356 11688
rect 28408 11636 28414 11688
rect 11388 11512 12940 11540
rect 11388 11500 11394 11512
rect 1104 11450 28888 11472
rect 1104 11398 2918 11450
rect 2970 11398 2982 11450
rect 3034 11398 3046 11450
rect 3098 11398 3110 11450
rect 3162 11398 3174 11450
rect 3226 11398 3238 11450
rect 3290 11398 10918 11450
rect 10970 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 11238 11450
rect 11290 11398 18918 11450
rect 18970 11398 18982 11450
rect 19034 11398 19046 11450
rect 19098 11398 19110 11450
rect 19162 11398 19174 11450
rect 19226 11398 19238 11450
rect 19290 11398 26918 11450
rect 26970 11398 26982 11450
rect 27034 11398 27046 11450
rect 27098 11398 27110 11450
rect 27162 11398 27174 11450
rect 27226 11398 27238 11450
rect 27290 11398 28888 11450
rect 1104 11376 28888 11398
rect 1581 11271 1639 11277
rect 1581 11237 1593 11271
rect 1627 11268 1639 11271
rect 1627 11240 2774 11268
rect 1627 11237 1639 11240
rect 1581 11231 1639 11237
rect 2746 11200 2774 11240
rect 11238 11200 11244 11212
rect 2746 11172 11244 11200
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 11422 11160 11428 11212
rect 11480 11200 11486 11212
rect 12066 11200 12072 11212
rect 11480 11172 12072 11200
rect 11480 11160 11486 11172
rect 12066 11160 12072 11172
rect 12124 11160 12130 11212
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 10686 11092 10692 11144
rect 10744 11092 10750 11144
rect 11054 11092 11060 11144
rect 11112 11092 11118 11144
rect 12342 11064 12348 11076
rect 12098 11036 12348 11064
rect 12342 11024 12348 11036
rect 12400 11024 12406 11076
rect 12434 11024 12440 11076
rect 12492 11073 12498 11076
rect 12492 11067 12541 11073
rect 12492 11033 12495 11067
rect 12529 11033 12541 11067
rect 12492 11027 12541 11033
rect 12492 11024 12498 11027
rect 1104 10906 28888 10928
rect 1104 10854 3658 10906
rect 3710 10854 3722 10906
rect 3774 10854 3786 10906
rect 3838 10854 3850 10906
rect 3902 10854 3914 10906
rect 3966 10854 3978 10906
rect 4030 10854 11658 10906
rect 11710 10854 11722 10906
rect 11774 10854 11786 10906
rect 11838 10854 11850 10906
rect 11902 10854 11914 10906
rect 11966 10854 11978 10906
rect 12030 10854 19658 10906
rect 19710 10854 19722 10906
rect 19774 10854 19786 10906
rect 19838 10854 19850 10906
rect 19902 10854 19914 10906
rect 19966 10854 19978 10906
rect 20030 10854 27658 10906
rect 27710 10854 27722 10906
rect 27774 10854 27786 10906
rect 27838 10854 27850 10906
rect 27902 10854 27914 10906
rect 27966 10854 27978 10906
rect 28030 10854 28888 10906
rect 1104 10832 28888 10854
rect 10594 10752 10600 10804
rect 10652 10792 10658 10804
rect 10873 10795 10931 10801
rect 10873 10792 10885 10795
rect 10652 10764 10885 10792
rect 10652 10752 10658 10764
rect 10873 10761 10885 10764
rect 10919 10761 10931 10795
rect 10873 10755 10931 10761
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 11112 10764 11529 10792
rect 11112 10752 11118 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 11977 10795 12035 10801
rect 11977 10761 11989 10795
rect 12023 10792 12035 10795
rect 12066 10792 12072 10804
rect 12023 10764 12072 10792
rect 12023 10761 12035 10764
rect 11977 10755 12035 10761
rect 12066 10752 12072 10764
rect 12124 10752 12130 10804
rect 10318 10684 10324 10736
rect 10376 10684 10382 10736
rect 10965 10727 11023 10733
rect 10965 10693 10977 10727
rect 11011 10724 11023 10727
rect 11330 10724 11336 10736
rect 11011 10696 11336 10724
rect 11011 10693 11023 10696
rect 10965 10687 11023 10693
rect 11330 10684 11336 10696
rect 11388 10684 11394 10736
rect 10336 10656 10364 10684
rect 11422 10656 11428 10668
rect 10336 10628 11428 10656
rect 11422 10616 11428 10628
rect 11480 10616 11486 10668
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10656 11943 10659
rect 12434 10656 12440 10668
rect 11931 10628 12440 10656
rect 11931 10625 11943 10628
rect 11885 10619 11943 10625
rect 12434 10616 12440 10628
rect 12492 10656 12498 10668
rect 28077 10659 28135 10665
rect 28077 10656 28089 10659
rect 12492 10628 28089 10656
rect 12492 10616 12498 10628
rect 28077 10625 28089 10628
rect 28123 10625 28135 10659
rect 28077 10619 28135 10625
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10588 10563 10591
rect 10778 10588 10784 10600
rect 10551 10560 10784 10588
rect 10551 10557 10563 10560
rect 10505 10551 10563 10557
rect 10778 10548 10784 10560
rect 10836 10588 10842 10600
rect 12069 10591 12127 10597
rect 12069 10588 12081 10591
rect 10836 10560 12081 10588
rect 10836 10548 10842 10560
rect 12069 10557 12081 10560
rect 12115 10588 12127 10591
rect 13170 10588 13176 10600
rect 12115 10560 13176 10588
rect 12115 10557 12127 10560
rect 12069 10551 12127 10557
rect 13170 10548 13176 10560
rect 13228 10548 13234 10600
rect 28350 10548 28356 10600
rect 28408 10548 28414 10600
rect 11333 10523 11391 10529
rect 11333 10489 11345 10523
rect 11379 10520 11391 10523
rect 11514 10520 11520 10532
rect 11379 10492 11520 10520
rect 11379 10489 11391 10492
rect 11333 10483 11391 10489
rect 11514 10480 11520 10492
rect 11572 10480 11578 10532
rect 12066 10412 12072 10464
rect 12124 10452 12130 10464
rect 12250 10452 12256 10464
rect 12124 10424 12256 10452
rect 12124 10412 12130 10424
rect 12250 10412 12256 10424
rect 12308 10412 12314 10464
rect 1104 10362 28888 10384
rect 1104 10310 2918 10362
rect 2970 10310 2982 10362
rect 3034 10310 3046 10362
rect 3098 10310 3110 10362
rect 3162 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 10918 10362
rect 10970 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 11238 10362
rect 11290 10310 18918 10362
rect 18970 10310 18982 10362
rect 19034 10310 19046 10362
rect 19098 10310 19110 10362
rect 19162 10310 19174 10362
rect 19226 10310 19238 10362
rect 19290 10310 26918 10362
rect 26970 10310 26982 10362
rect 27034 10310 27046 10362
rect 27098 10310 27110 10362
rect 27162 10310 27174 10362
rect 27226 10310 27238 10362
rect 27290 10310 28888 10362
rect 1104 10288 28888 10310
rect 12621 10183 12679 10189
rect 12621 10149 12633 10183
rect 12667 10149 12679 10183
rect 12621 10143 12679 10149
rect 11057 10115 11115 10121
rect 11057 10081 11069 10115
rect 11103 10112 11115 10115
rect 12636 10112 12664 10143
rect 11103 10084 12664 10112
rect 11103 10081 11115 10084
rect 11057 10075 11115 10081
rect 13170 10072 13176 10124
rect 13228 10072 13234 10124
rect 1394 10004 1400 10056
rect 1452 10004 1458 10056
rect 10686 10004 10692 10056
rect 10744 10004 10750 10056
rect 12483 10047 12541 10053
rect 12483 10013 12495 10047
rect 12529 10044 12541 10047
rect 12989 10047 13047 10053
rect 12989 10044 13001 10047
rect 12529 10016 13001 10044
rect 12529 10013 12541 10016
rect 12483 10007 12541 10013
rect 12989 10013 13001 10016
rect 13035 10044 13047 10047
rect 28077 10047 28135 10053
rect 28077 10044 28089 10047
rect 13035 10016 28089 10044
rect 13035 10013 13047 10016
rect 12989 10007 13047 10013
rect 28077 10013 28089 10016
rect 28123 10013 28135 10047
rect 28077 10007 28135 10013
rect 12342 9976 12348 9988
rect 12098 9948 12348 9976
rect 12342 9936 12348 9948
rect 12400 9936 12406 9988
rect 28350 9936 28356 9988
rect 28408 9936 28414 9988
rect 1578 9868 1584 9920
rect 1636 9868 1642 9920
rect 11330 9868 11336 9920
rect 11388 9908 11394 9920
rect 13081 9911 13139 9917
rect 13081 9908 13093 9911
rect 11388 9880 13093 9908
rect 11388 9868 11394 9880
rect 13081 9877 13093 9880
rect 13127 9877 13139 9911
rect 13081 9871 13139 9877
rect 1104 9818 28888 9840
rect 1104 9766 3658 9818
rect 3710 9766 3722 9818
rect 3774 9766 3786 9818
rect 3838 9766 3850 9818
rect 3902 9766 3914 9818
rect 3966 9766 3978 9818
rect 4030 9766 11658 9818
rect 11710 9766 11722 9818
rect 11774 9766 11786 9818
rect 11838 9766 11850 9818
rect 11902 9766 11914 9818
rect 11966 9766 11978 9818
rect 12030 9766 19658 9818
rect 19710 9766 19722 9818
rect 19774 9766 19786 9818
rect 19838 9766 19850 9818
rect 19902 9766 19914 9818
rect 19966 9766 19978 9818
rect 20030 9766 27658 9818
rect 27710 9766 27722 9818
rect 27774 9766 27786 9818
rect 27838 9766 27850 9818
rect 27902 9766 27914 9818
rect 27966 9766 27978 9818
rect 28030 9766 28888 9818
rect 1104 9744 28888 9766
rect 1578 9664 1584 9716
rect 1636 9704 1642 9716
rect 10873 9707 10931 9713
rect 10873 9704 10885 9707
rect 1636 9676 10885 9704
rect 1636 9664 1642 9676
rect 10873 9673 10885 9676
rect 10919 9673 10931 9707
rect 10873 9667 10931 9673
rect 10686 9596 10692 9648
rect 10744 9636 10750 9648
rect 10744 9608 11560 9636
rect 10744 9596 10750 9608
rect 1394 9528 1400 9580
rect 1452 9528 1458 9580
rect 11532 9577 11560 9608
rect 12250 9596 12256 9648
rect 12308 9596 12314 9648
rect 10965 9571 11023 9577
rect 10965 9537 10977 9571
rect 11011 9537 11023 9571
rect 10965 9531 11023 9537
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 10778 9460 10784 9512
rect 10836 9460 10842 9512
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 10778 9364 10784 9376
rect 1627 9336 10784 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 10980 9364 11008 9531
rect 11885 9503 11943 9509
rect 11885 9500 11897 9503
rect 11348 9472 11897 9500
rect 11348 9441 11376 9472
rect 11885 9469 11897 9472
rect 11931 9469 11943 9503
rect 11885 9463 11943 9469
rect 11333 9435 11391 9441
rect 11333 9401 11345 9435
rect 11379 9401 11391 9435
rect 11333 9395 11391 9401
rect 13311 9367 13369 9373
rect 13311 9364 13323 9367
rect 10980 9336 13323 9364
rect 13311 9333 13323 9336
rect 13357 9364 13369 9367
rect 28074 9364 28080 9376
rect 13357 9336 28080 9364
rect 13357 9333 13369 9336
rect 13311 9327 13369 9333
rect 28074 9324 28080 9336
rect 28132 9324 28138 9376
rect 1104 9274 28888 9296
rect 1104 9222 2918 9274
rect 2970 9222 2982 9274
rect 3034 9222 3046 9274
rect 3098 9222 3110 9274
rect 3162 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 10918 9274
rect 10970 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 11238 9274
rect 11290 9222 18918 9274
rect 18970 9222 18982 9274
rect 19034 9222 19046 9274
rect 19098 9222 19110 9274
rect 19162 9222 19174 9274
rect 19226 9222 19238 9274
rect 19290 9222 26918 9274
rect 26970 9222 26982 9274
rect 27034 9222 27046 9274
rect 27098 9222 27110 9274
rect 27162 9222 27174 9274
rect 27226 9222 27238 9274
rect 27290 9222 28888 9274
rect 1104 9200 28888 9222
rect 11885 9163 11943 9169
rect 11885 9129 11897 9163
rect 11931 9160 11943 9163
rect 12250 9160 12256 9172
rect 11931 9132 12256 9160
rect 11931 9129 11943 9132
rect 11885 9123 11943 9129
rect 12250 9120 12256 9132
rect 12308 9120 12314 9172
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8956 12035 8959
rect 12066 8956 12072 8968
rect 12023 8928 12072 8956
rect 12023 8925 12035 8928
rect 11977 8919 12035 8925
rect 12066 8916 12072 8928
rect 12124 8916 12130 8968
rect 28074 8916 28080 8968
rect 28132 8916 28138 8968
rect 28350 8848 28356 8900
rect 28408 8848 28414 8900
rect 1104 8730 28888 8752
rect 1104 8678 3658 8730
rect 3710 8678 3722 8730
rect 3774 8678 3786 8730
rect 3838 8678 3850 8730
rect 3902 8678 3914 8730
rect 3966 8678 3978 8730
rect 4030 8678 11658 8730
rect 11710 8678 11722 8730
rect 11774 8678 11786 8730
rect 11838 8678 11850 8730
rect 11902 8678 11914 8730
rect 11966 8678 11978 8730
rect 12030 8678 19658 8730
rect 19710 8678 19722 8730
rect 19774 8678 19786 8730
rect 19838 8678 19850 8730
rect 19902 8678 19914 8730
rect 19966 8678 19978 8730
rect 20030 8678 27658 8730
rect 27710 8678 27722 8730
rect 27774 8678 27786 8730
rect 27838 8678 27850 8730
rect 27902 8678 27914 8730
rect 27966 8678 27978 8730
rect 28030 8678 28888 8730
rect 1104 8656 28888 8678
rect 10778 8576 10784 8628
rect 10836 8616 10842 8628
rect 10873 8619 10931 8625
rect 10873 8616 10885 8619
rect 10836 8588 10885 8616
rect 10836 8576 10842 8588
rect 10873 8585 10885 8588
rect 10919 8585 10931 8619
rect 10873 8579 10931 8585
rect 11900 8588 13308 8616
rect 10965 8551 11023 8557
rect 10965 8517 10977 8551
rect 11011 8548 11023 8551
rect 11900 8548 11928 8588
rect 11011 8520 11928 8548
rect 11011 8517 11023 8520
rect 10965 8511 11023 8517
rect 12066 8508 12072 8560
rect 12124 8548 12130 8560
rect 12124 8520 12282 8548
rect 12124 8508 12130 8520
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 11330 8480 11336 8492
rect 2746 8452 11336 8480
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 2746 8344 2774 8452
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 13280 8480 13308 8588
rect 28077 8483 28135 8489
rect 28077 8480 28089 8483
rect 13280 8452 28089 8480
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8412 10839 8415
rect 11422 8412 11428 8424
rect 10827 8384 11428 8412
rect 10827 8381 10839 8384
rect 10781 8375 10839 8381
rect 11422 8372 11428 8384
rect 11480 8372 11486 8424
rect 13280 8421 13308 8452
rect 28077 8449 28089 8452
rect 28123 8449 28135 8483
rect 28077 8443 28135 8449
rect 11517 8415 11575 8421
rect 11517 8381 11529 8415
rect 11563 8381 11575 8415
rect 11793 8415 11851 8421
rect 11793 8412 11805 8415
rect 11517 8375 11575 8381
rect 11624 8384 11805 8412
rect 11532 8344 11560 8375
rect 1627 8316 2774 8344
rect 10704 8316 11560 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 10704 8288 10732 8316
rect 10686 8236 10692 8288
rect 10744 8236 10750 8288
rect 11333 8279 11391 8285
rect 11333 8245 11345 8279
rect 11379 8276 11391 8279
rect 11624 8276 11652 8384
rect 11793 8381 11805 8384
rect 11839 8381 11851 8415
rect 11793 8375 11851 8381
rect 13265 8415 13323 8421
rect 13265 8381 13277 8415
rect 13311 8381 13323 8415
rect 13265 8375 13323 8381
rect 28350 8372 28356 8424
rect 28408 8372 28414 8424
rect 11379 8248 11652 8276
rect 11379 8245 11391 8248
rect 11333 8239 11391 8245
rect 1104 8186 28888 8208
rect 1104 8134 2918 8186
rect 2970 8134 2982 8186
rect 3034 8134 3046 8186
rect 3098 8134 3110 8186
rect 3162 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 10918 8186
rect 10970 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 11238 8186
rect 11290 8134 18918 8186
rect 18970 8134 18982 8186
rect 19034 8134 19046 8186
rect 19098 8134 19110 8186
rect 19162 8134 19174 8186
rect 19226 8134 19238 8186
rect 19290 8134 26918 8186
rect 26970 8134 26982 8186
rect 27034 8134 27046 8186
rect 27098 8134 27110 8186
rect 27162 8134 27174 8186
rect 27226 8134 27238 8186
rect 27290 8134 28888 8186
rect 1104 8112 28888 8134
rect 10686 7896 10692 7948
rect 10744 7896 10750 7948
rect 1394 7828 1400 7880
rect 1452 7828 1458 7880
rect 12066 7828 12072 7880
rect 12124 7868 12130 7880
rect 12342 7868 12348 7880
rect 12124 7840 12348 7868
rect 12124 7828 12130 7840
rect 12342 7828 12348 7840
rect 12400 7828 12406 7880
rect 10962 7760 10968 7812
rect 11020 7760 11026 7812
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 10134 7732 10140 7744
rect 1627 7704 10140 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 10134 7692 10140 7704
rect 10192 7692 10198 7744
rect 12434 7692 12440 7744
rect 12492 7732 12498 7744
rect 28074 7732 28080 7744
rect 12492 7704 28080 7732
rect 12492 7692 12498 7704
rect 28074 7692 28080 7704
rect 28132 7692 28138 7744
rect 1104 7642 28888 7664
rect 1104 7590 3658 7642
rect 3710 7590 3722 7642
rect 3774 7590 3786 7642
rect 3838 7590 3850 7642
rect 3902 7590 3914 7642
rect 3966 7590 3978 7642
rect 4030 7590 11658 7642
rect 11710 7590 11722 7642
rect 11774 7590 11786 7642
rect 11838 7590 11850 7642
rect 11902 7590 11914 7642
rect 11966 7590 11978 7642
rect 12030 7590 19658 7642
rect 19710 7590 19722 7642
rect 19774 7590 19786 7642
rect 19838 7590 19850 7642
rect 19902 7590 19914 7642
rect 19966 7590 19978 7642
rect 20030 7590 27658 7642
rect 27710 7590 27722 7642
rect 27774 7590 27786 7642
rect 27838 7590 27850 7642
rect 27902 7590 27914 7642
rect 27966 7590 27978 7642
rect 28030 7590 28888 7642
rect 1104 7568 28888 7590
rect 10962 7488 10968 7540
rect 11020 7528 11026 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 11020 7500 11529 7528
rect 11020 7488 11026 7500
rect 11517 7497 11529 7500
rect 11563 7497 11575 7531
rect 11517 7491 11575 7497
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 12434 7528 12440 7540
rect 11931 7500 12440 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 11330 7420 11336 7472
rect 11388 7460 11394 7472
rect 11977 7463 12035 7469
rect 11977 7460 11989 7463
rect 11388 7432 11989 7460
rect 11388 7420 11394 7432
rect 11977 7429 11989 7432
rect 12023 7429 12035 7463
rect 11977 7423 12035 7429
rect 28074 7352 28080 7404
rect 28132 7352 28138 7404
rect 11422 7284 11428 7336
rect 11480 7324 11486 7336
rect 12069 7327 12127 7333
rect 12069 7324 12081 7327
rect 11480 7296 12081 7324
rect 11480 7284 11486 7296
rect 12069 7293 12081 7296
rect 12115 7293 12127 7327
rect 12069 7287 12127 7293
rect 28350 7284 28356 7336
rect 28408 7284 28414 7336
rect 1104 7098 28888 7120
rect 1104 7046 2918 7098
rect 2970 7046 2982 7098
rect 3034 7046 3046 7098
rect 3098 7046 3110 7098
rect 3162 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 10918 7098
rect 10970 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 11238 7098
rect 11290 7046 18918 7098
rect 18970 7046 18982 7098
rect 19034 7046 19046 7098
rect 19098 7046 19110 7098
rect 19162 7046 19174 7098
rect 19226 7046 19238 7098
rect 19290 7046 26918 7098
rect 26970 7046 26982 7098
rect 27034 7046 27046 7098
rect 27098 7046 27110 7098
rect 27162 7046 27174 7098
rect 27226 7046 27238 7098
rect 27290 7046 28888 7098
rect 1104 7024 28888 7046
rect 10686 6808 10692 6860
rect 10744 6848 10750 6860
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 10744 6820 11069 6848
rect 10744 6808 10750 6820
rect 1394 6740 1400 6792
rect 1452 6740 1458 6792
rect 10888 6789 10916 6820
rect 11057 6817 11069 6820
rect 11103 6817 11115 6851
rect 11057 6811 11115 6817
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6780 10931 6783
rect 10919 6752 10953 6780
rect 10919 6749 10931 6752
rect 10873 6743 10931 6749
rect 12802 6740 12808 6792
rect 12860 6740 12866 6792
rect 28074 6740 28080 6792
rect 28132 6740 28138 6792
rect 28350 6672 28356 6724
rect 28408 6672 28414 6724
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 10042 6644 10048 6656
rect 1627 6616 10048 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 1104 6554 28888 6576
rect 1104 6502 3658 6554
rect 3710 6502 3722 6554
rect 3774 6502 3786 6554
rect 3838 6502 3850 6554
rect 3902 6502 3914 6554
rect 3966 6502 3978 6554
rect 4030 6502 11658 6554
rect 11710 6502 11722 6554
rect 11774 6502 11786 6554
rect 11838 6502 11850 6554
rect 11902 6502 11914 6554
rect 11966 6502 11978 6554
rect 12030 6502 19658 6554
rect 19710 6502 19722 6554
rect 19774 6502 19786 6554
rect 19838 6502 19850 6554
rect 19902 6502 19914 6554
rect 19966 6502 19978 6554
rect 20030 6502 27658 6554
rect 27710 6502 27722 6554
rect 27774 6502 27786 6554
rect 27838 6502 27850 6554
rect 27902 6502 27914 6554
rect 27966 6502 27978 6554
rect 28030 6502 28888 6554
rect 1104 6480 28888 6502
rect 10042 6400 10048 6452
rect 10100 6400 10106 6452
rect 10134 6400 10140 6452
rect 10192 6440 10198 6452
rect 10873 6443 10931 6449
rect 10873 6440 10885 6443
rect 10192 6412 10885 6440
rect 10192 6400 10198 6412
rect 10873 6409 10885 6412
rect 10919 6409 10931 6443
rect 10873 6403 10931 6409
rect 10686 6332 10692 6384
rect 10744 6372 10750 6384
rect 10744 6344 11560 6372
rect 10744 6332 10750 6344
rect 1394 6264 1400 6316
rect 1452 6264 1458 6316
rect 10134 6264 10140 6316
rect 10192 6264 10198 6316
rect 11532 6313 11560 6344
rect 12250 6332 12256 6384
rect 12308 6332 12314 6384
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6304 11023 6307
rect 11517 6307 11575 6313
rect 11011 6276 11284 6304
rect 11011 6273 11023 6276
rect 10965 6267 11023 6273
rect 9953 6239 10011 6245
rect 9953 6205 9965 6239
rect 9999 6236 10011 6239
rect 10689 6239 10747 6245
rect 10689 6236 10701 6239
rect 9999 6208 10701 6236
rect 9999 6205 10011 6208
rect 9953 6199 10011 6205
rect 10689 6205 10701 6208
rect 10735 6236 10747 6239
rect 10778 6236 10784 6248
rect 10735 6208 10784 6236
rect 10735 6205 10747 6208
rect 10689 6199 10747 6205
rect 10778 6196 10784 6208
rect 10836 6196 10842 6248
rect 10410 6168 10416 6180
rect 2746 6140 10416 6168
rect 1581 6103 1639 6109
rect 1581 6069 1593 6103
rect 1627 6100 1639 6103
rect 2746 6100 2774 6140
rect 10410 6128 10416 6140
rect 10468 6128 10474 6180
rect 1627 6072 2774 6100
rect 1627 6069 1639 6072
rect 1581 6063 1639 6069
rect 10502 6060 10508 6112
rect 10560 6060 10566 6112
rect 11256 6100 11284 6276
rect 11517 6273 11529 6307
rect 11563 6273 11575 6307
rect 11517 6267 11575 6273
rect 11793 6239 11851 6245
rect 11793 6236 11805 6239
rect 11348 6208 11805 6236
rect 11348 6177 11376 6208
rect 11793 6205 11805 6208
rect 11839 6205 11851 6239
rect 11793 6199 11851 6205
rect 11333 6171 11391 6177
rect 11333 6137 11345 6171
rect 11379 6137 11391 6171
rect 11333 6131 11391 6137
rect 13265 6103 13323 6109
rect 13265 6100 13277 6103
rect 11256 6072 13277 6100
rect 13265 6069 13277 6072
rect 13311 6100 13323 6103
rect 28074 6100 28080 6112
rect 13311 6072 28080 6100
rect 13311 6069 13323 6072
rect 13265 6063 13323 6069
rect 28074 6060 28080 6072
rect 28132 6060 28138 6112
rect 1104 6010 28888 6032
rect 1104 5958 2918 6010
rect 2970 5958 2982 6010
rect 3034 5958 3046 6010
rect 3098 5958 3110 6010
rect 3162 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 10918 6010
rect 10970 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 11238 6010
rect 11290 5958 18918 6010
rect 18970 5958 18982 6010
rect 19034 5958 19046 6010
rect 19098 5958 19110 6010
rect 19162 5958 19174 6010
rect 19226 5958 19238 6010
rect 19290 5958 26918 6010
rect 26970 5958 26982 6010
rect 27034 5958 27046 6010
rect 27098 5958 27110 6010
rect 27162 5958 27174 6010
rect 27226 5958 27238 6010
rect 27290 5958 28888 6010
rect 1104 5936 28888 5958
rect 10134 5856 10140 5908
rect 10192 5896 10198 5908
rect 10192 5868 12480 5896
rect 10192 5856 10198 5868
rect 10502 5788 10508 5840
rect 10560 5828 10566 5840
rect 10560 5800 10824 5828
rect 10560 5788 10566 5800
rect 10686 5720 10692 5772
rect 10744 5720 10750 5772
rect 10796 5760 10824 5800
rect 12452 5769 12480 5868
rect 10965 5763 11023 5769
rect 10965 5760 10977 5763
rect 10796 5732 10977 5760
rect 10965 5729 10977 5732
rect 11011 5729 11023 5763
rect 10965 5723 11023 5729
rect 12437 5763 12495 5769
rect 12437 5729 12449 5763
rect 12483 5729 12495 5763
rect 12437 5723 12495 5729
rect 12452 5692 12480 5723
rect 28077 5695 28135 5701
rect 28077 5692 28089 5695
rect 12452 5664 28089 5692
rect 28077 5661 28089 5664
rect 28123 5661 28135 5695
rect 28077 5655 28135 5661
rect 12250 5624 12256 5636
rect 12190 5596 12256 5624
rect 12250 5584 12256 5596
rect 12308 5584 12314 5636
rect 28350 5584 28356 5636
rect 28408 5584 28414 5636
rect 1104 5466 28888 5488
rect 1104 5414 3658 5466
rect 3710 5414 3722 5466
rect 3774 5414 3786 5466
rect 3838 5414 3850 5466
rect 3902 5414 3914 5466
rect 3966 5414 3978 5466
rect 4030 5414 11658 5466
rect 11710 5414 11722 5466
rect 11774 5414 11786 5466
rect 11838 5414 11850 5466
rect 11902 5414 11914 5466
rect 11966 5414 11978 5466
rect 12030 5414 19658 5466
rect 19710 5414 19722 5466
rect 19774 5414 19786 5466
rect 19838 5414 19850 5466
rect 19902 5414 19914 5466
rect 19966 5414 19978 5466
rect 20030 5414 27658 5466
rect 27710 5414 27722 5466
rect 27774 5414 27786 5466
rect 27838 5414 27850 5466
rect 27902 5414 27914 5466
rect 27966 5414 27978 5466
rect 28030 5414 28888 5466
rect 1104 5392 28888 5414
rect 10410 5312 10416 5364
rect 10468 5352 10474 5364
rect 11977 5355 12035 5361
rect 11977 5352 11989 5355
rect 10468 5324 11989 5352
rect 10468 5312 10474 5324
rect 11977 5321 11989 5324
rect 12023 5321 12035 5355
rect 11977 5315 12035 5321
rect 1394 5176 1400 5228
rect 1452 5176 1458 5228
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5216 11943 5219
rect 12526 5216 12532 5228
rect 11931 5188 12532 5216
rect 11931 5185 11943 5188
rect 11885 5179 11943 5185
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 28074 5176 28080 5228
rect 28132 5176 28138 5228
rect 10778 5108 10784 5160
rect 10836 5148 10842 5160
rect 12069 5151 12127 5157
rect 12069 5148 12081 5151
rect 10836 5120 12081 5148
rect 10836 5108 10842 5120
rect 12069 5117 12081 5120
rect 12115 5148 12127 5151
rect 12986 5148 12992 5160
rect 12115 5120 12992 5148
rect 12115 5117 12127 5120
rect 12069 5111 12127 5117
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 28350 5108 28356 5160
rect 28408 5108 28414 5160
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 7558 5012 7564 5024
rect 1627 4984 7564 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 7558 4972 7564 4984
rect 7616 4972 7622 5024
rect 11514 4972 11520 5024
rect 11572 4972 11578 5024
rect 1104 4922 28888 4944
rect 1104 4870 2918 4922
rect 2970 4870 2982 4922
rect 3034 4870 3046 4922
rect 3098 4870 3110 4922
rect 3162 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 10918 4922
rect 10970 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 11238 4922
rect 11290 4870 18918 4922
rect 18970 4870 18982 4922
rect 19034 4870 19046 4922
rect 19098 4870 19110 4922
rect 19162 4870 19174 4922
rect 19226 4870 19238 4922
rect 19290 4870 26918 4922
rect 26970 4870 26982 4922
rect 27034 4870 27046 4922
rect 27098 4870 27110 4922
rect 27162 4870 27174 4922
rect 27226 4870 27238 4922
rect 27290 4870 28888 4922
rect 1104 4848 28888 4870
rect 7558 4768 7564 4820
rect 7616 4808 7622 4820
rect 7616 4780 12940 4808
rect 7616 4768 7622 4780
rect 10594 4632 10600 4684
rect 10652 4632 10658 4684
rect 10873 4675 10931 4681
rect 10873 4641 10885 4675
rect 10919 4672 10931 4675
rect 11514 4672 11520 4684
rect 10919 4644 11520 4672
rect 10919 4641 10931 4644
rect 10873 4635 10931 4641
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 12250 4672 12256 4684
rect 11992 4644 12256 4672
rect 1394 4564 1400 4616
rect 1452 4564 1458 4616
rect 11992 4590 12020 4644
rect 12250 4632 12256 4644
rect 12308 4632 12314 4684
rect 12912 4681 12940 4780
rect 12897 4675 12955 4681
rect 12897 4641 12909 4675
rect 12943 4641 12955 4675
rect 12897 4635 12955 4641
rect 12986 4632 12992 4684
rect 13044 4632 13050 4684
rect 12710 4604 12716 4616
rect 12176 4576 12716 4604
rect 1581 4471 1639 4477
rect 1581 4437 1593 4471
rect 1627 4468 1639 4471
rect 12176 4468 12204 4576
rect 12710 4564 12716 4576
rect 12768 4564 12774 4616
rect 12526 4536 12532 4548
rect 12360 4508 12532 4536
rect 12360 4477 12388 4508
rect 12526 4496 12532 4508
rect 12584 4496 12590 4548
rect 1627 4440 12204 4468
rect 12345 4471 12403 4477
rect 1627 4437 1639 4440
rect 1581 4431 1639 4437
rect 12345 4437 12357 4471
rect 12391 4437 12403 4471
rect 12345 4431 12403 4437
rect 12434 4428 12440 4480
rect 12492 4428 12498 4480
rect 12802 4428 12808 4480
rect 12860 4428 12866 4480
rect 1104 4378 28888 4400
rect 1104 4326 3658 4378
rect 3710 4326 3722 4378
rect 3774 4326 3786 4378
rect 3838 4326 3850 4378
rect 3902 4326 3914 4378
rect 3966 4326 3978 4378
rect 4030 4326 11658 4378
rect 11710 4326 11722 4378
rect 11774 4326 11786 4378
rect 11838 4326 11850 4378
rect 11902 4326 11914 4378
rect 11966 4326 11978 4378
rect 12030 4326 19658 4378
rect 19710 4326 19722 4378
rect 19774 4326 19786 4378
rect 19838 4326 19850 4378
rect 19902 4326 19914 4378
rect 19966 4326 19978 4378
rect 20030 4326 27658 4378
rect 27710 4326 27722 4378
rect 27774 4326 27786 4378
rect 27838 4326 27850 4378
rect 27902 4326 27914 4378
rect 27966 4326 27978 4378
rect 28030 4326 28888 4378
rect 1104 4304 28888 4326
rect 12526 4224 12532 4276
rect 12584 4264 12590 4276
rect 28074 4264 28080 4276
rect 12584 4236 28080 4264
rect 12584 4224 12590 4236
rect 28074 4224 28080 4236
rect 28132 4224 28138 4276
rect 11149 4199 11207 4205
rect 11149 4165 11161 4199
rect 11195 4196 11207 4199
rect 11514 4196 11520 4208
rect 11195 4168 11520 4196
rect 11195 4165 11207 4168
rect 11149 4159 11207 4165
rect 11514 4156 11520 4168
rect 11572 4156 11578 4208
rect 12250 4156 12256 4208
rect 12308 4156 12314 4208
rect 11333 4131 11391 4137
rect 11333 4097 11345 4131
rect 11379 4128 11391 4131
rect 11422 4128 11428 4140
rect 11379 4100 11428 4128
rect 11379 4097 11391 4100
rect 11333 4091 11391 4097
rect 11422 4088 11428 4100
rect 11480 4088 11486 4140
rect 28077 4131 28135 4137
rect 28077 4128 28089 4131
rect 13280 4100 28089 4128
rect 10594 4020 10600 4072
rect 10652 4060 10658 4072
rect 11517 4063 11575 4069
rect 11517 4060 11529 4063
rect 10652 4032 11529 4060
rect 10652 4020 10658 4032
rect 11517 4029 11529 4032
rect 11563 4029 11575 4063
rect 11517 4023 11575 4029
rect 11793 4063 11851 4069
rect 11793 4029 11805 4063
rect 11839 4060 11851 4063
rect 12434 4060 12440 4072
rect 11839 4032 12440 4060
rect 11839 4029 11851 4032
rect 11793 4023 11851 4029
rect 12434 4020 12440 4032
rect 12492 4020 12498 4072
rect 12802 4020 12808 4072
rect 12860 4060 12866 4072
rect 13280 4069 13308 4100
rect 28077 4097 28089 4100
rect 28123 4097 28135 4131
rect 28077 4091 28135 4097
rect 13265 4063 13323 4069
rect 13265 4060 13277 4063
rect 12860 4032 13277 4060
rect 12860 4020 12866 4032
rect 13265 4029 13277 4032
rect 13311 4029 13323 4063
rect 13265 4023 13323 4029
rect 28350 4020 28356 4072
rect 28408 4020 28414 4072
rect 1104 3834 28888 3856
rect 1104 3782 2918 3834
rect 2970 3782 2982 3834
rect 3034 3782 3046 3834
rect 3098 3782 3110 3834
rect 3162 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 10918 3834
rect 10970 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 11238 3834
rect 11290 3782 18918 3834
rect 18970 3782 18982 3834
rect 19034 3782 19046 3834
rect 19098 3782 19110 3834
rect 19162 3782 19174 3834
rect 19226 3782 19238 3834
rect 19290 3782 26918 3834
rect 26970 3782 26982 3834
rect 27034 3782 27046 3834
rect 27098 3782 27110 3834
rect 27162 3782 27174 3834
rect 27226 3782 27238 3834
rect 27290 3782 28888 3834
rect 1104 3760 28888 3782
rect 10321 3723 10379 3729
rect 10321 3689 10333 3723
rect 10367 3720 10379 3723
rect 10686 3720 10692 3732
rect 10367 3692 10692 3720
rect 10367 3689 10379 3692
rect 10321 3683 10379 3689
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 12437 3723 12495 3729
rect 12437 3720 12449 3723
rect 11900 3692 12449 3720
rect 10594 3544 10600 3596
rect 10652 3544 10658 3596
rect 10873 3587 10931 3593
rect 10873 3553 10885 3587
rect 10919 3584 10931 3587
rect 11900 3584 11928 3692
rect 12437 3689 12449 3692
rect 12483 3689 12495 3723
rect 12437 3683 12495 3689
rect 10919 3556 11928 3584
rect 12345 3587 12403 3593
rect 10919 3553 10931 3556
rect 10873 3547 10931 3553
rect 12345 3553 12357 3587
rect 12391 3553 12403 3587
rect 12345 3547 12403 3553
rect 1394 3476 1400 3528
rect 1452 3476 1458 3528
rect 12360 3516 12388 3547
rect 12710 3544 12716 3596
rect 12768 3584 12774 3596
rect 12897 3587 12955 3593
rect 12897 3584 12909 3587
rect 12768 3556 12909 3584
rect 12768 3544 12774 3556
rect 12897 3553 12909 3556
rect 12943 3553 12955 3587
rect 12897 3547 12955 3553
rect 12986 3544 12992 3596
rect 13044 3544 13050 3596
rect 12805 3519 12863 3525
rect 12805 3516 12817 3519
rect 12360 3488 12817 3516
rect 12805 3485 12817 3488
rect 12851 3516 12863 3519
rect 28077 3519 28135 3525
rect 28077 3516 28089 3519
rect 12851 3488 28089 3516
rect 12851 3485 12863 3488
rect 12805 3479 12863 3485
rect 28077 3485 28089 3488
rect 28123 3485 28135 3519
rect 28077 3479 28135 3485
rect 10413 3451 10471 3457
rect 10413 3417 10425 3451
rect 10459 3448 10471 3451
rect 11146 3448 11152 3460
rect 10459 3420 11152 3448
rect 10459 3417 10471 3420
rect 10413 3411 10471 3417
rect 11146 3408 11152 3420
rect 11204 3408 11210 3460
rect 12250 3448 12256 3460
rect 12098 3420 12256 3448
rect 12250 3408 12256 3420
rect 12308 3408 12314 3460
rect 12342 3408 12348 3460
rect 12400 3448 12406 3460
rect 13265 3451 13323 3457
rect 13265 3448 13277 3451
rect 12400 3420 13277 3448
rect 12400 3408 12406 3420
rect 13265 3417 13277 3420
rect 13311 3417 13323 3451
rect 13265 3411 13323 3417
rect 13449 3451 13507 3457
rect 13449 3417 13461 3451
rect 13495 3417 13507 3451
rect 13449 3411 13507 3417
rect 1581 3383 1639 3389
rect 1581 3349 1593 3383
rect 1627 3380 1639 3383
rect 10226 3380 10232 3392
rect 1627 3352 10232 3380
rect 1627 3349 1639 3352
rect 1581 3343 1639 3349
rect 10226 3340 10232 3352
rect 10284 3340 10290 3392
rect 12158 3340 12164 3392
rect 12216 3380 12222 3392
rect 13464 3380 13492 3411
rect 28350 3408 28356 3460
rect 28408 3408 28414 3460
rect 12216 3352 13492 3380
rect 12216 3340 12222 3352
rect 1104 3290 28888 3312
rect 1104 3238 3658 3290
rect 3710 3238 3722 3290
rect 3774 3238 3786 3290
rect 3838 3238 3850 3290
rect 3902 3238 3914 3290
rect 3966 3238 3978 3290
rect 4030 3238 11658 3290
rect 11710 3238 11722 3290
rect 11774 3238 11786 3290
rect 11838 3238 11850 3290
rect 11902 3238 11914 3290
rect 11966 3238 11978 3290
rect 12030 3238 19658 3290
rect 19710 3238 19722 3290
rect 19774 3238 19786 3290
rect 19838 3238 19850 3290
rect 19902 3238 19914 3290
rect 19966 3238 19978 3290
rect 20030 3238 27658 3290
rect 27710 3238 27722 3290
rect 27774 3238 27786 3290
rect 27838 3238 27850 3290
rect 27902 3238 27914 3290
rect 27966 3238 27978 3290
rect 28030 3238 28888 3290
rect 1104 3216 28888 3238
rect 10226 3136 10232 3188
rect 10284 3176 10290 3188
rect 10873 3179 10931 3185
rect 10873 3176 10885 3179
rect 10284 3148 10885 3176
rect 10284 3136 10290 3148
rect 10873 3145 10885 3148
rect 10919 3145 10931 3179
rect 10873 3139 10931 3145
rect 11054 3136 11060 3188
rect 11112 3176 11118 3188
rect 11514 3176 11520 3188
rect 11112 3148 11520 3176
rect 11112 3136 11118 3148
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 10594 3068 10600 3120
rect 10652 3108 10658 3120
rect 10652 3080 11560 3108
rect 10652 3068 10658 3080
rect 842 3000 848 3052
rect 900 3040 906 3052
rect 11532 3049 11560 3080
rect 12250 3068 12256 3120
rect 12308 3068 12314 3120
rect 1397 3043 1455 3049
rect 1397 3040 1409 3043
rect 900 3012 1409 3040
rect 900 3000 906 3012
rect 1397 3009 1409 3012
rect 1443 3009 1455 3043
rect 1397 3003 1455 3009
rect 10965 3043 11023 3049
rect 10965 3009 10977 3043
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 10686 2932 10692 2984
rect 10744 2932 10750 2984
rect 1581 2839 1639 2845
rect 1581 2805 1593 2839
rect 1627 2836 1639 2839
rect 10870 2836 10876 2848
rect 1627 2808 10876 2836
rect 1627 2805 1639 2808
rect 1581 2799 1639 2805
rect 10870 2796 10876 2808
rect 10928 2796 10934 2848
rect 10980 2836 11008 3003
rect 11793 2975 11851 2981
rect 11793 2972 11805 2975
rect 11348 2944 11805 2972
rect 11348 2913 11376 2944
rect 11793 2941 11805 2944
rect 11839 2941 11851 2975
rect 11793 2935 11851 2941
rect 11333 2907 11391 2913
rect 11333 2873 11345 2907
rect 11379 2873 11391 2907
rect 11333 2867 11391 2873
rect 13265 2839 13323 2845
rect 13265 2836 13277 2839
rect 10980 2808 13277 2836
rect 13265 2805 13277 2808
rect 13311 2836 13323 2839
rect 20622 2836 20628 2848
rect 13311 2808 20628 2836
rect 13311 2805 13323 2808
rect 13265 2799 13323 2805
rect 20622 2796 20628 2808
rect 20680 2796 20686 2848
rect 1104 2746 28888 2768
rect 1104 2694 2918 2746
rect 2970 2694 2982 2746
rect 3034 2694 3046 2746
rect 3098 2694 3110 2746
rect 3162 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 10918 2746
rect 10970 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 11238 2746
rect 11290 2694 18918 2746
rect 18970 2694 18982 2746
rect 19034 2694 19046 2746
rect 19098 2694 19110 2746
rect 19162 2694 19174 2746
rect 19226 2694 19238 2746
rect 19290 2694 26918 2746
rect 26970 2694 26982 2746
rect 27034 2694 27046 2746
rect 27098 2694 27110 2746
rect 27162 2694 27174 2746
rect 27226 2694 27238 2746
rect 27290 2694 28888 2746
rect 1104 2672 28888 2694
rect 11885 2635 11943 2641
rect 11885 2601 11897 2635
rect 11931 2632 11943 2635
rect 12250 2632 12256 2644
rect 11931 2604 12256 2632
rect 11931 2601 11943 2604
rect 11885 2595 11943 2601
rect 12250 2592 12256 2604
rect 12308 2592 12314 2644
rect 842 2388 848 2440
rect 900 2428 906 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 900 2400 1409 2428
rect 900 2388 906 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2428 12035 2431
rect 12342 2428 12348 2440
rect 12023 2400 12348 2428
rect 12023 2397 12035 2400
rect 11977 2391 12035 2397
rect 12342 2388 12348 2400
rect 12400 2388 12406 2440
rect 20622 2388 20628 2440
rect 20680 2428 20686 2440
rect 28077 2431 28135 2437
rect 28077 2428 28089 2431
rect 20680 2400 28089 2428
rect 20680 2388 20686 2400
rect 28077 2397 28089 2400
rect 28123 2397 28135 2431
rect 28077 2391 28135 2397
rect 28350 2320 28356 2372
rect 28408 2320 28414 2372
rect 1581 2295 1639 2301
rect 1581 2261 1593 2295
rect 1627 2292 1639 2295
rect 12158 2292 12164 2304
rect 1627 2264 12164 2292
rect 1627 2261 1639 2264
rect 1581 2255 1639 2261
rect 12158 2252 12164 2264
rect 12216 2252 12222 2304
rect 1104 2202 28888 2224
rect 1104 2150 3658 2202
rect 3710 2150 3722 2202
rect 3774 2150 3786 2202
rect 3838 2150 3850 2202
rect 3902 2150 3914 2202
rect 3966 2150 3978 2202
rect 4030 2150 11658 2202
rect 11710 2150 11722 2202
rect 11774 2150 11786 2202
rect 11838 2150 11850 2202
rect 11902 2150 11914 2202
rect 11966 2150 11978 2202
rect 12030 2150 19658 2202
rect 19710 2150 19722 2202
rect 19774 2150 19786 2202
rect 19838 2150 19850 2202
rect 19902 2150 19914 2202
rect 19966 2150 19978 2202
rect 20030 2150 27658 2202
rect 27710 2150 27722 2202
rect 27774 2150 27786 2202
rect 27838 2150 27850 2202
rect 27902 2150 27914 2202
rect 27966 2150 27978 2202
rect 28030 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 2918 27718 2970 27770
rect 2982 27718 3034 27770
rect 3046 27718 3098 27770
rect 3110 27718 3162 27770
rect 3174 27718 3226 27770
rect 3238 27718 3290 27770
rect 10918 27718 10970 27770
rect 10982 27718 11034 27770
rect 11046 27718 11098 27770
rect 11110 27718 11162 27770
rect 11174 27718 11226 27770
rect 11238 27718 11290 27770
rect 18918 27718 18970 27770
rect 18982 27718 19034 27770
rect 19046 27718 19098 27770
rect 19110 27718 19162 27770
rect 19174 27718 19226 27770
rect 19238 27718 19290 27770
rect 26918 27718 26970 27770
rect 26982 27718 27034 27770
rect 27046 27718 27098 27770
rect 27110 27718 27162 27770
rect 27174 27718 27226 27770
rect 27238 27718 27290 27770
rect 1032 27548 1084 27600
rect 940 27480 992 27532
rect 848 27412 900 27464
rect 10968 27548 11020 27600
rect 28356 27523 28408 27532
rect 28356 27489 28365 27523
rect 28365 27489 28399 27523
rect 28399 27489 28408 27523
rect 28356 27480 28408 27489
rect 12348 27412 12400 27464
rect 21272 27412 21324 27464
rect 1584 27319 1636 27328
rect 1584 27285 1593 27319
rect 1593 27285 1627 27319
rect 1627 27285 1636 27319
rect 1584 27276 1636 27285
rect 11428 27344 11480 27396
rect 12164 27276 12216 27328
rect 3658 27174 3710 27226
rect 3722 27174 3774 27226
rect 3786 27174 3838 27226
rect 3850 27174 3902 27226
rect 3914 27174 3966 27226
rect 3978 27174 4030 27226
rect 11658 27174 11710 27226
rect 11722 27174 11774 27226
rect 11786 27174 11838 27226
rect 11850 27174 11902 27226
rect 11914 27174 11966 27226
rect 11978 27174 12030 27226
rect 19658 27174 19710 27226
rect 19722 27174 19774 27226
rect 19786 27174 19838 27226
rect 19850 27174 19902 27226
rect 19914 27174 19966 27226
rect 19978 27174 20030 27226
rect 27658 27174 27710 27226
rect 27722 27174 27774 27226
rect 27786 27174 27838 27226
rect 27850 27174 27902 27226
rect 27914 27174 27966 27226
rect 27978 27174 28030 27226
rect 1584 27072 1636 27124
rect 10968 27072 11020 27124
rect 11428 27072 11480 27124
rect 13268 27004 13320 27056
rect 9220 26800 9272 26852
rect 12256 26936 12308 26988
rect 12440 26936 12492 26988
rect 21364 26936 21416 26988
rect 12164 26911 12216 26920
rect 12164 26877 12173 26911
rect 12173 26877 12207 26911
rect 12207 26877 12216 26911
rect 12164 26868 12216 26877
rect 28356 26911 28408 26920
rect 28356 26877 28365 26911
rect 28365 26877 28399 26911
rect 28399 26877 28408 26911
rect 28356 26868 28408 26877
rect 21272 26800 21324 26852
rect 10600 26775 10652 26784
rect 10600 26741 10609 26775
rect 10609 26741 10643 26775
rect 10643 26741 10652 26775
rect 10600 26732 10652 26741
rect 11428 26732 11480 26784
rect 12072 26732 12124 26784
rect 2918 26630 2970 26682
rect 2982 26630 3034 26682
rect 3046 26630 3098 26682
rect 3110 26630 3162 26682
rect 3174 26630 3226 26682
rect 3238 26630 3290 26682
rect 10918 26630 10970 26682
rect 10982 26630 11034 26682
rect 11046 26630 11098 26682
rect 11110 26630 11162 26682
rect 11174 26630 11226 26682
rect 11238 26630 11290 26682
rect 18918 26630 18970 26682
rect 18982 26630 19034 26682
rect 19046 26630 19098 26682
rect 19110 26630 19162 26682
rect 19174 26630 19226 26682
rect 19238 26630 19290 26682
rect 26918 26630 26970 26682
rect 26982 26630 27034 26682
rect 27046 26630 27098 26682
rect 27110 26630 27162 26682
rect 27174 26630 27226 26682
rect 27238 26630 27290 26682
rect 9220 26528 9272 26580
rect 10416 26392 10468 26444
rect 10600 26435 10652 26444
rect 10600 26401 10609 26435
rect 10609 26401 10643 26435
rect 10643 26401 10652 26435
rect 10600 26392 10652 26401
rect 11428 26435 11480 26444
rect 11428 26401 11437 26435
rect 11437 26401 11471 26435
rect 11471 26401 11480 26435
rect 11428 26392 11480 26401
rect 12164 26392 12216 26444
rect 848 26324 900 26376
rect 11336 26324 11388 26376
rect 12256 26324 12308 26376
rect 21364 26324 21416 26376
rect 13268 26256 13320 26308
rect 13544 26256 13596 26308
rect 28356 26299 28408 26308
rect 28356 26265 28365 26299
rect 28365 26265 28399 26299
rect 28399 26265 28408 26299
rect 28356 26256 28408 26265
rect 12072 26188 12124 26240
rect 12992 26231 13044 26240
rect 12992 26197 13001 26231
rect 13001 26197 13035 26231
rect 13035 26197 13044 26231
rect 12992 26188 13044 26197
rect 3658 26086 3710 26138
rect 3722 26086 3774 26138
rect 3786 26086 3838 26138
rect 3850 26086 3902 26138
rect 3914 26086 3966 26138
rect 3978 26086 4030 26138
rect 11658 26086 11710 26138
rect 11722 26086 11774 26138
rect 11786 26086 11838 26138
rect 11850 26086 11902 26138
rect 11914 26086 11966 26138
rect 11978 26086 12030 26138
rect 19658 26086 19710 26138
rect 19722 26086 19774 26138
rect 19786 26086 19838 26138
rect 19850 26086 19902 26138
rect 19914 26086 19966 26138
rect 19978 26086 20030 26138
rect 27658 26086 27710 26138
rect 27722 26086 27774 26138
rect 27786 26086 27838 26138
rect 27850 26086 27902 26138
rect 27914 26086 27966 26138
rect 27978 26086 28030 26138
rect 10416 25984 10468 26036
rect 12072 25984 12124 26036
rect 13544 25984 13596 26036
rect 848 25848 900 25900
rect 11612 25848 11664 25900
rect 11336 25780 11388 25832
rect 12992 25780 13044 25832
rect 10600 25644 10652 25696
rect 11428 25644 11480 25696
rect 12072 25644 12124 25696
rect 2918 25542 2970 25594
rect 2982 25542 3034 25594
rect 3046 25542 3098 25594
rect 3110 25542 3162 25594
rect 3174 25542 3226 25594
rect 3238 25542 3290 25594
rect 10918 25542 10970 25594
rect 10982 25542 11034 25594
rect 11046 25542 11098 25594
rect 11110 25542 11162 25594
rect 11174 25542 11226 25594
rect 11238 25542 11290 25594
rect 18918 25542 18970 25594
rect 18982 25542 19034 25594
rect 19046 25542 19098 25594
rect 19110 25542 19162 25594
rect 19174 25542 19226 25594
rect 19238 25542 19290 25594
rect 26918 25542 26970 25594
rect 26982 25542 27034 25594
rect 27046 25542 27098 25594
rect 27110 25542 27162 25594
rect 27174 25542 27226 25594
rect 27238 25542 27290 25594
rect 11428 25347 11480 25356
rect 11428 25313 11437 25347
rect 11437 25313 11471 25347
rect 11471 25313 11480 25347
rect 11428 25304 11480 25313
rect 11612 25304 11664 25356
rect 11336 25236 11388 25288
rect 28356 25211 28408 25220
rect 28356 25177 28365 25211
rect 28365 25177 28399 25211
rect 28399 25177 28408 25211
rect 28356 25168 28408 25177
rect 12808 25100 12860 25152
rect 3658 24998 3710 25050
rect 3722 24998 3774 25050
rect 3786 24998 3838 25050
rect 3850 24998 3902 25050
rect 3914 24998 3966 25050
rect 3978 24998 4030 25050
rect 11658 24998 11710 25050
rect 11722 24998 11774 25050
rect 11786 24998 11838 25050
rect 11850 24998 11902 25050
rect 11914 24998 11966 25050
rect 11978 24998 12030 25050
rect 19658 24998 19710 25050
rect 19722 24998 19774 25050
rect 19786 24998 19838 25050
rect 19850 24998 19902 25050
rect 19914 24998 19966 25050
rect 19978 24998 20030 25050
rect 27658 24998 27710 25050
rect 27722 24998 27774 25050
rect 27786 24998 27838 25050
rect 27850 24998 27902 25050
rect 27914 24998 27966 25050
rect 27978 24998 28030 25050
rect 12808 24828 12860 24880
rect 848 24760 900 24812
rect 13360 24760 13412 24812
rect 11336 24692 11388 24744
rect 12992 24692 13044 24744
rect 28356 24735 28408 24744
rect 28356 24701 28365 24735
rect 28365 24701 28399 24735
rect 28399 24701 28408 24735
rect 28356 24692 28408 24701
rect 11428 24556 11480 24608
rect 2918 24454 2970 24506
rect 2982 24454 3034 24506
rect 3046 24454 3098 24506
rect 3110 24454 3162 24506
rect 3174 24454 3226 24506
rect 3238 24454 3290 24506
rect 10918 24454 10970 24506
rect 10982 24454 11034 24506
rect 11046 24454 11098 24506
rect 11110 24454 11162 24506
rect 11174 24454 11226 24506
rect 11238 24454 11290 24506
rect 18918 24454 18970 24506
rect 18982 24454 19034 24506
rect 19046 24454 19098 24506
rect 19110 24454 19162 24506
rect 19174 24454 19226 24506
rect 19238 24454 19290 24506
rect 26918 24454 26970 24506
rect 26982 24454 27034 24506
rect 27046 24454 27098 24506
rect 27110 24454 27162 24506
rect 27174 24454 27226 24506
rect 27238 24454 27290 24506
rect 12992 24395 13044 24404
rect 12992 24361 13001 24395
rect 13001 24361 13035 24395
rect 13035 24361 13044 24395
rect 12992 24352 13044 24361
rect 12256 24284 12308 24336
rect 10600 24216 10652 24268
rect 848 24148 900 24200
rect 11336 24148 11388 24200
rect 11520 24148 11572 24200
rect 13360 24191 13412 24200
rect 13360 24157 13369 24191
rect 13369 24157 13403 24191
rect 13403 24157 13412 24191
rect 13360 24148 13412 24157
rect 1584 24055 1636 24064
rect 1584 24021 1593 24055
rect 1593 24021 1627 24055
rect 1627 24021 1636 24055
rect 1584 24012 1636 24021
rect 12624 24080 12676 24132
rect 28080 24080 28132 24132
rect 12716 24012 12768 24064
rect 3658 23910 3710 23962
rect 3722 23910 3774 23962
rect 3786 23910 3838 23962
rect 3850 23910 3902 23962
rect 3914 23910 3966 23962
rect 3978 23910 4030 23962
rect 11658 23910 11710 23962
rect 11722 23910 11774 23962
rect 11786 23910 11838 23962
rect 11850 23910 11902 23962
rect 11914 23910 11966 23962
rect 11978 23910 12030 23962
rect 19658 23910 19710 23962
rect 19722 23910 19774 23962
rect 19786 23910 19838 23962
rect 19850 23910 19902 23962
rect 19914 23910 19966 23962
rect 19978 23910 20030 23962
rect 27658 23910 27710 23962
rect 27722 23910 27774 23962
rect 27786 23910 27838 23962
rect 27850 23910 27902 23962
rect 27914 23910 27966 23962
rect 27978 23910 28030 23962
rect 1584 23808 1636 23860
rect 11520 23851 11572 23860
rect 11520 23817 11529 23851
rect 11529 23817 11563 23851
rect 11563 23817 11572 23851
rect 11520 23808 11572 23817
rect 12624 23808 12676 23860
rect 11428 23740 11480 23792
rect 14556 23672 14608 23724
rect 28080 23715 28132 23724
rect 28080 23681 28089 23715
rect 28089 23681 28123 23715
rect 28123 23681 28132 23715
rect 28080 23672 28132 23681
rect 12072 23647 12124 23656
rect 12072 23613 12081 23647
rect 12081 23613 12115 23647
rect 12115 23613 12124 23647
rect 12072 23604 12124 23613
rect 28356 23647 28408 23656
rect 28356 23613 28365 23647
rect 28365 23613 28399 23647
rect 28399 23613 28408 23647
rect 28356 23604 28408 23613
rect 2918 23366 2970 23418
rect 2982 23366 3034 23418
rect 3046 23366 3098 23418
rect 3110 23366 3162 23418
rect 3174 23366 3226 23418
rect 3238 23366 3290 23418
rect 10918 23366 10970 23418
rect 10982 23366 11034 23418
rect 11046 23366 11098 23418
rect 11110 23366 11162 23418
rect 11174 23366 11226 23418
rect 11238 23366 11290 23418
rect 18918 23366 18970 23418
rect 18982 23366 19034 23418
rect 19046 23366 19098 23418
rect 19110 23366 19162 23418
rect 19174 23366 19226 23418
rect 19238 23366 19290 23418
rect 26918 23366 26970 23418
rect 26982 23366 27034 23418
rect 27046 23366 27098 23418
rect 27110 23366 27162 23418
rect 27174 23366 27226 23418
rect 27238 23366 27290 23418
rect 12072 23196 12124 23248
rect 14556 23171 14608 23180
rect 14556 23137 14565 23171
rect 14565 23137 14599 23171
rect 14599 23137 14608 23171
rect 14556 23128 14608 23137
rect 14648 23171 14700 23180
rect 14648 23137 14657 23171
rect 14657 23137 14691 23171
rect 14691 23137 14700 23171
rect 14648 23128 14700 23137
rect 848 23060 900 23112
rect 12164 23060 12216 23112
rect 14924 23060 14976 23112
rect 11520 23035 11572 23044
rect 11520 23001 11529 23035
rect 11529 23001 11563 23035
rect 11563 23001 11572 23035
rect 11520 22992 11572 23001
rect 28356 23035 28408 23044
rect 28356 23001 28365 23035
rect 28365 23001 28399 23035
rect 28399 23001 28408 23035
rect 28356 22992 28408 23001
rect 11152 22924 11204 22976
rect 13084 22924 13136 22976
rect 13452 22924 13504 22976
rect 3658 22822 3710 22874
rect 3722 22822 3774 22874
rect 3786 22822 3838 22874
rect 3850 22822 3902 22874
rect 3914 22822 3966 22874
rect 3978 22822 4030 22874
rect 11658 22822 11710 22874
rect 11722 22822 11774 22874
rect 11786 22822 11838 22874
rect 11850 22822 11902 22874
rect 11914 22822 11966 22874
rect 11978 22822 12030 22874
rect 19658 22822 19710 22874
rect 19722 22822 19774 22874
rect 19786 22822 19838 22874
rect 19850 22822 19902 22874
rect 19914 22822 19966 22874
rect 19978 22822 20030 22874
rect 27658 22822 27710 22874
rect 27722 22822 27774 22874
rect 27786 22822 27838 22874
rect 27850 22822 27902 22874
rect 27914 22822 27966 22874
rect 27978 22822 28030 22874
rect 11152 22720 11204 22772
rect 14924 22720 14976 22772
rect 12624 22652 12676 22704
rect 13820 22652 13872 22704
rect 848 22584 900 22636
rect 12440 22627 12492 22636
rect 12440 22593 12449 22627
rect 12449 22593 12483 22627
rect 12483 22593 12492 22627
rect 12440 22584 12492 22593
rect 13452 22627 13504 22636
rect 13452 22593 13461 22627
rect 13461 22593 13495 22627
rect 13495 22593 13504 22627
rect 13452 22584 13504 22593
rect 12072 22559 12124 22568
rect 12072 22525 12081 22559
rect 12081 22525 12115 22559
rect 12115 22525 12124 22559
rect 12072 22516 12124 22525
rect 13084 22559 13136 22568
rect 13084 22525 13093 22559
rect 13093 22525 13127 22559
rect 13127 22525 13136 22559
rect 13084 22516 13136 22525
rect 12716 22448 12768 22500
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 11428 22380 11480 22432
rect 2918 22278 2970 22330
rect 2982 22278 3034 22330
rect 3046 22278 3098 22330
rect 3110 22278 3162 22330
rect 3174 22278 3226 22330
rect 3238 22278 3290 22330
rect 10918 22278 10970 22330
rect 10982 22278 11034 22330
rect 11046 22278 11098 22330
rect 11110 22278 11162 22330
rect 11174 22278 11226 22330
rect 11238 22278 11290 22330
rect 18918 22278 18970 22330
rect 18982 22278 19034 22330
rect 19046 22278 19098 22330
rect 19110 22278 19162 22330
rect 19174 22278 19226 22330
rect 19238 22278 19290 22330
rect 26918 22278 26970 22330
rect 26982 22278 27034 22330
rect 27046 22278 27098 22330
rect 27110 22278 27162 22330
rect 27174 22278 27226 22330
rect 27238 22278 27290 22330
rect 1584 22176 1636 22228
rect 11336 22040 11388 22092
rect 13084 22040 13136 22092
rect 14648 22108 14700 22160
rect 11428 22015 11480 22024
rect 11428 21981 11437 22015
rect 11437 21981 11471 22015
rect 11471 21981 11480 22015
rect 11428 21972 11480 21981
rect 12716 21972 12768 22024
rect 13728 21972 13780 22024
rect 12624 21904 12676 21956
rect 13452 21836 13504 21888
rect 14832 21904 14884 21956
rect 17868 21904 17920 21956
rect 28356 21947 28408 21956
rect 28356 21913 28365 21947
rect 28365 21913 28399 21947
rect 28399 21913 28408 21947
rect 28356 21904 28408 21913
rect 3658 21734 3710 21786
rect 3722 21734 3774 21786
rect 3786 21734 3838 21786
rect 3850 21734 3902 21786
rect 3914 21734 3966 21786
rect 3978 21734 4030 21786
rect 11658 21734 11710 21786
rect 11722 21734 11774 21786
rect 11786 21734 11838 21786
rect 11850 21734 11902 21786
rect 11914 21734 11966 21786
rect 11978 21734 12030 21786
rect 19658 21734 19710 21786
rect 19722 21734 19774 21786
rect 19786 21734 19838 21786
rect 19850 21734 19902 21786
rect 19914 21734 19966 21786
rect 19978 21734 20030 21786
rect 27658 21734 27710 21786
rect 27722 21734 27774 21786
rect 27786 21734 27838 21786
rect 27850 21734 27902 21786
rect 27914 21734 27966 21786
rect 27978 21734 28030 21786
rect 13728 21632 13780 21684
rect 14832 21632 14884 21684
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 13084 21539 13136 21548
rect 13084 21505 13093 21539
rect 13093 21505 13127 21539
rect 13127 21505 13136 21539
rect 13084 21496 13136 21505
rect 13452 21539 13504 21548
rect 13452 21505 13461 21539
rect 13461 21505 13495 21539
rect 13495 21505 13504 21539
rect 13452 21496 13504 21505
rect 17868 21496 17920 21548
rect 28356 21471 28408 21480
rect 28356 21437 28365 21471
rect 28365 21437 28399 21471
rect 28399 21437 28408 21471
rect 28356 21428 28408 21437
rect 14556 21292 14608 21344
rect 2918 21190 2970 21242
rect 2982 21190 3034 21242
rect 3046 21190 3098 21242
rect 3110 21190 3162 21242
rect 3174 21190 3226 21242
rect 3238 21190 3290 21242
rect 10918 21190 10970 21242
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 11238 21190 11290 21242
rect 18918 21190 18970 21242
rect 18982 21190 19034 21242
rect 19046 21190 19098 21242
rect 19110 21190 19162 21242
rect 19174 21190 19226 21242
rect 19238 21190 19290 21242
rect 26918 21190 26970 21242
rect 26982 21190 27034 21242
rect 27046 21190 27098 21242
rect 27110 21190 27162 21242
rect 27174 21190 27226 21242
rect 27238 21190 27290 21242
rect 12164 21020 12216 21072
rect 14556 20995 14608 21004
rect 14556 20961 14565 20995
rect 14565 20961 14599 20995
rect 14599 20961 14608 20995
rect 14556 20952 14608 20961
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 14648 20816 14700 20868
rect 11336 20748 11388 20800
rect 13912 20748 13964 20800
rect 3658 20646 3710 20698
rect 3722 20646 3774 20698
rect 3786 20646 3838 20698
rect 3850 20646 3902 20698
rect 3914 20646 3966 20698
rect 3978 20646 4030 20698
rect 11658 20646 11710 20698
rect 11722 20646 11774 20698
rect 11786 20646 11838 20698
rect 11850 20646 11902 20698
rect 11914 20646 11966 20698
rect 11978 20646 12030 20698
rect 19658 20646 19710 20698
rect 19722 20646 19774 20698
rect 19786 20646 19838 20698
rect 19850 20646 19902 20698
rect 19914 20646 19966 20698
rect 19978 20646 20030 20698
rect 27658 20646 27710 20698
rect 27722 20646 27774 20698
rect 27786 20646 27838 20698
rect 27850 20646 27902 20698
rect 27914 20646 27966 20698
rect 27978 20646 28030 20698
rect 12440 20544 12492 20596
rect 14648 20408 14700 20460
rect 12348 20340 12400 20392
rect 13912 20340 13964 20392
rect 28356 20383 28408 20392
rect 28356 20349 28365 20383
rect 28365 20349 28399 20383
rect 28399 20349 28408 20383
rect 28356 20340 28408 20349
rect 2918 20102 2970 20154
rect 2982 20102 3034 20154
rect 3046 20102 3098 20154
rect 3110 20102 3162 20154
rect 3174 20102 3226 20154
rect 3238 20102 3290 20154
rect 10918 20102 10970 20154
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 11238 20102 11290 20154
rect 18918 20102 18970 20154
rect 18982 20102 19034 20154
rect 19046 20102 19098 20154
rect 19110 20102 19162 20154
rect 19174 20102 19226 20154
rect 19238 20102 19290 20154
rect 26918 20102 26970 20154
rect 26982 20102 27034 20154
rect 27046 20102 27098 20154
rect 27110 20102 27162 20154
rect 27174 20102 27226 20154
rect 27238 20102 27290 20154
rect 12348 19864 12400 19916
rect 13820 19907 13872 19916
rect 13820 19873 13829 19907
rect 13829 19873 13863 19907
rect 13863 19873 13872 19907
rect 13820 19864 13872 19873
rect 1400 19839 1452 19848
rect 1400 19805 1409 19839
rect 1409 19805 1443 19839
rect 1443 19805 1452 19839
rect 1400 19796 1452 19805
rect 11428 19839 11480 19848
rect 11428 19805 11437 19839
rect 11437 19805 11471 19839
rect 11471 19805 11480 19839
rect 11428 19796 11480 19805
rect 12256 19796 12308 19848
rect 12440 19728 12492 19780
rect 28356 19771 28408 19780
rect 28356 19737 28365 19771
rect 28365 19737 28399 19771
rect 28399 19737 28408 19771
rect 28356 19728 28408 19737
rect 12992 19660 13044 19712
rect 13544 19703 13596 19712
rect 13544 19669 13553 19703
rect 13553 19669 13587 19703
rect 13587 19669 13596 19703
rect 13544 19660 13596 19669
rect 3658 19558 3710 19610
rect 3722 19558 3774 19610
rect 3786 19558 3838 19610
rect 3850 19558 3902 19610
rect 3914 19558 3966 19610
rect 3978 19558 4030 19610
rect 11658 19558 11710 19610
rect 11722 19558 11774 19610
rect 11786 19558 11838 19610
rect 11850 19558 11902 19610
rect 11914 19558 11966 19610
rect 11978 19558 12030 19610
rect 19658 19558 19710 19610
rect 19722 19558 19774 19610
rect 19786 19558 19838 19610
rect 19850 19558 19902 19610
rect 19914 19558 19966 19610
rect 19978 19558 20030 19610
rect 27658 19558 27710 19610
rect 27722 19558 27774 19610
rect 27786 19558 27838 19610
rect 27850 19558 27902 19610
rect 27914 19558 27966 19610
rect 27978 19558 28030 19610
rect 848 19320 900 19372
rect 11428 19456 11480 19508
rect 12256 19456 12308 19508
rect 13544 19456 13596 19508
rect 11336 19388 11388 19440
rect 12348 19320 12400 19372
rect 13728 19388 13780 19440
rect 11428 19252 11480 19304
rect 12164 19252 12216 19304
rect 12992 19363 13044 19372
rect 12992 19329 13001 19363
rect 13001 19329 13035 19363
rect 13035 19329 13044 19363
rect 12992 19320 13044 19329
rect 23480 19320 23532 19372
rect 14556 19252 14608 19304
rect 2918 19014 2970 19066
rect 2982 19014 3034 19066
rect 3046 19014 3098 19066
rect 3110 19014 3162 19066
rect 3174 19014 3226 19066
rect 3238 19014 3290 19066
rect 10918 19014 10970 19066
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 11238 19014 11290 19066
rect 18918 19014 18970 19066
rect 18982 19014 19034 19066
rect 19046 19014 19098 19066
rect 19110 19014 19162 19066
rect 19174 19014 19226 19066
rect 19238 19014 19290 19066
rect 26918 19014 26970 19066
rect 26982 19014 27034 19066
rect 27046 19014 27098 19066
rect 27110 19014 27162 19066
rect 27174 19014 27226 19066
rect 27238 19014 27290 19066
rect 13820 18776 13872 18828
rect 14648 18819 14700 18828
rect 14648 18785 14657 18819
rect 14657 18785 14691 18819
rect 14691 18785 14700 18819
rect 14648 18776 14700 18785
rect 14556 18751 14608 18760
rect 14556 18717 14565 18751
rect 14565 18717 14599 18751
rect 14599 18717 14608 18751
rect 14556 18708 14608 18717
rect 23480 18708 23532 18760
rect 12348 18640 12400 18692
rect 28356 18683 28408 18692
rect 28356 18649 28365 18683
rect 28365 18649 28399 18683
rect 28399 18649 28408 18683
rect 28356 18640 28408 18649
rect 12716 18572 12768 18624
rect 14464 18615 14516 18624
rect 14464 18581 14473 18615
rect 14473 18581 14507 18615
rect 14507 18581 14516 18615
rect 14464 18572 14516 18581
rect 3658 18470 3710 18522
rect 3722 18470 3774 18522
rect 3786 18470 3838 18522
rect 3850 18470 3902 18522
rect 3914 18470 3966 18522
rect 3978 18470 4030 18522
rect 11658 18470 11710 18522
rect 11722 18470 11774 18522
rect 11786 18470 11838 18522
rect 11850 18470 11902 18522
rect 11914 18470 11966 18522
rect 11978 18470 12030 18522
rect 19658 18470 19710 18522
rect 19722 18470 19774 18522
rect 19786 18470 19838 18522
rect 19850 18470 19902 18522
rect 19914 18470 19966 18522
rect 19978 18470 20030 18522
rect 27658 18470 27710 18522
rect 27722 18470 27774 18522
rect 27786 18470 27838 18522
rect 27850 18470 27902 18522
rect 27914 18470 27966 18522
rect 27978 18470 28030 18522
rect 14556 18368 14608 18420
rect 13728 18300 13780 18352
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 12716 18275 12768 18284
rect 12716 18241 12725 18275
rect 12725 18241 12759 18275
rect 12759 18241 12768 18275
rect 12716 18232 12768 18241
rect 14464 18232 14516 18284
rect 12348 18207 12400 18216
rect 12348 18173 12357 18207
rect 12357 18173 12391 18207
rect 12391 18173 12400 18207
rect 12348 18164 12400 18173
rect 28356 18207 28408 18216
rect 28356 18173 28365 18207
rect 28365 18173 28399 18207
rect 28399 18173 28408 18207
rect 28356 18164 28408 18173
rect 2918 17926 2970 17978
rect 2982 17926 3034 17978
rect 3046 17926 3098 17978
rect 3110 17926 3162 17978
rect 3174 17926 3226 17978
rect 3238 17926 3290 17978
rect 10918 17926 10970 17978
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 11238 17926 11290 17978
rect 18918 17926 18970 17978
rect 18982 17926 19034 17978
rect 19046 17926 19098 17978
rect 19110 17926 19162 17978
rect 19174 17926 19226 17978
rect 19238 17926 19290 17978
rect 26918 17926 26970 17978
rect 26982 17926 27034 17978
rect 27046 17926 27098 17978
rect 27110 17926 27162 17978
rect 27174 17926 27226 17978
rect 27238 17926 27290 17978
rect 12348 17824 12400 17876
rect 14556 17731 14608 17740
rect 14556 17697 14565 17731
rect 14565 17697 14599 17731
rect 14599 17697 14608 17731
rect 14556 17688 14608 17697
rect 14648 17731 14700 17740
rect 14648 17697 14657 17731
rect 14657 17697 14691 17731
rect 14691 17697 14700 17731
rect 14648 17688 14700 17697
rect 1400 17663 1452 17672
rect 1400 17629 1409 17663
rect 1409 17629 1443 17663
rect 1443 17629 1452 17663
rect 1400 17620 1452 17629
rect 11520 17620 11572 17672
rect 12164 17663 12216 17672
rect 12164 17629 12173 17663
rect 12173 17629 12207 17663
rect 12207 17629 12216 17663
rect 12164 17620 12216 17629
rect 11336 17484 11388 17536
rect 12440 17484 12492 17536
rect 14464 17527 14516 17536
rect 14464 17493 14473 17527
rect 14473 17493 14507 17527
rect 14507 17493 14516 17527
rect 14464 17484 14516 17493
rect 3658 17382 3710 17434
rect 3722 17382 3774 17434
rect 3786 17382 3838 17434
rect 3850 17382 3902 17434
rect 3914 17382 3966 17434
rect 3978 17382 4030 17434
rect 11658 17382 11710 17434
rect 11722 17382 11774 17434
rect 11786 17382 11838 17434
rect 11850 17382 11902 17434
rect 11914 17382 11966 17434
rect 11978 17382 12030 17434
rect 19658 17382 19710 17434
rect 19722 17382 19774 17434
rect 19786 17382 19838 17434
rect 19850 17382 19902 17434
rect 19914 17382 19966 17434
rect 19978 17382 20030 17434
rect 27658 17382 27710 17434
rect 27722 17382 27774 17434
rect 27786 17382 27838 17434
rect 27850 17382 27902 17434
rect 27914 17382 27966 17434
rect 27978 17382 28030 17434
rect 12440 17187 12492 17196
rect 12440 17153 12449 17187
rect 12449 17153 12483 17187
rect 12483 17153 12492 17187
rect 12440 17144 12492 17153
rect 11520 17076 11572 17128
rect 12348 17076 12400 17128
rect 12992 17076 13044 17128
rect 13728 17212 13780 17264
rect 14464 17144 14516 17196
rect 28356 17119 28408 17128
rect 28356 17085 28365 17119
rect 28365 17085 28399 17119
rect 28399 17085 28408 17119
rect 28356 17076 28408 17085
rect 2918 16838 2970 16890
rect 2982 16838 3034 16890
rect 3046 16838 3098 16890
rect 3110 16838 3162 16890
rect 3174 16838 3226 16890
rect 3238 16838 3290 16890
rect 10918 16838 10970 16890
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 11238 16838 11290 16890
rect 18918 16838 18970 16890
rect 18982 16838 19034 16890
rect 19046 16838 19098 16890
rect 19110 16838 19162 16890
rect 19174 16838 19226 16890
rect 19238 16838 19290 16890
rect 26918 16838 26970 16890
rect 26982 16838 27034 16890
rect 27046 16838 27098 16890
rect 27110 16838 27162 16890
rect 27174 16838 27226 16890
rect 27238 16838 27290 16890
rect 1400 16575 1452 16584
rect 1400 16541 1409 16575
rect 1409 16541 1443 16575
rect 1443 16541 1452 16575
rect 1400 16532 1452 16541
rect 11520 16532 11572 16584
rect 12072 16532 12124 16584
rect 21364 16532 21416 16584
rect 10876 16396 10928 16448
rect 28356 16507 28408 16516
rect 28356 16473 28365 16507
rect 28365 16473 28399 16507
rect 28399 16473 28408 16507
rect 28356 16464 28408 16473
rect 12440 16396 12492 16448
rect 12900 16396 12952 16448
rect 13452 16396 13504 16448
rect 3658 16294 3710 16346
rect 3722 16294 3774 16346
rect 3786 16294 3838 16346
rect 3850 16294 3902 16346
rect 3914 16294 3966 16346
rect 3978 16294 4030 16346
rect 11658 16294 11710 16346
rect 11722 16294 11774 16346
rect 11786 16294 11838 16346
rect 11850 16294 11902 16346
rect 11914 16294 11966 16346
rect 11978 16294 12030 16346
rect 19658 16294 19710 16346
rect 19722 16294 19774 16346
rect 19786 16294 19838 16346
rect 19850 16294 19902 16346
rect 19914 16294 19966 16346
rect 19978 16294 20030 16346
rect 27658 16294 27710 16346
rect 27722 16294 27774 16346
rect 27786 16294 27838 16346
rect 27850 16294 27902 16346
rect 27914 16294 27966 16346
rect 27978 16294 28030 16346
rect 10876 16235 10928 16244
rect 10876 16201 10885 16235
rect 10885 16201 10919 16235
rect 10919 16201 10928 16235
rect 10876 16192 10928 16201
rect 12440 16124 12492 16176
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 10692 16031 10744 16040
rect 10692 15997 10701 16031
rect 10701 15997 10735 16031
rect 10735 15997 10744 16031
rect 10692 15988 10744 15997
rect 10784 15852 10836 15904
rect 11520 16099 11572 16108
rect 11520 16065 11529 16099
rect 11529 16065 11563 16099
rect 11563 16065 11572 16099
rect 11520 16056 11572 16065
rect 28080 15852 28132 15904
rect 2918 15750 2970 15802
rect 2982 15750 3034 15802
rect 3046 15750 3098 15802
rect 3110 15750 3162 15802
rect 3174 15750 3226 15802
rect 3238 15750 3290 15802
rect 10918 15750 10970 15802
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 11238 15750 11290 15802
rect 18918 15750 18970 15802
rect 18982 15750 19034 15802
rect 19046 15750 19098 15802
rect 19110 15750 19162 15802
rect 19174 15750 19226 15802
rect 19238 15750 19290 15802
rect 26918 15750 26970 15802
rect 26982 15750 27034 15802
rect 27046 15750 27098 15802
rect 27110 15750 27162 15802
rect 27174 15750 27226 15802
rect 27238 15750 27290 15802
rect 11428 15648 11480 15700
rect 12072 15691 12124 15700
rect 12072 15657 12081 15691
rect 12081 15657 12115 15691
rect 12115 15657 12124 15691
rect 12072 15648 12124 15657
rect 10692 15580 10744 15632
rect 11336 15512 11388 15564
rect 14648 15512 14700 15564
rect 11428 15444 11480 15496
rect 12256 15444 12308 15496
rect 28080 15487 28132 15496
rect 28080 15453 28089 15487
rect 28089 15453 28123 15487
rect 28123 15453 28132 15487
rect 28080 15444 28132 15453
rect 11612 15419 11664 15428
rect 11612 15385 11621 15419
rect 11621 15385 11655 15419
rect 11655 15385 11664 15419
rect 11612 15376 11664 15385
rect 13452 15376 13504 15428
rect 21364 15376 21416 15428
rect 28356 15419 28408 15428
rect 28356 15385 28365 15419
rect 28365 15385 28399 15419
rect 28399 15385 28408 15419
rect 28356 15376 28408 15385
rect 12624 15308 12676 15360
rect 3658 15206 3710 15258
rect 3722 15206 3774 15258
rect 3786 15206 3838 15258
rect 3850 15206 3902 15258
rect 3914 15206 3966 15258
rect 3978 15206 4030 15258
rect 11658 15206 11710 15258
rect 11722 15206 11774 15258
rect 11786 15206 11838 15258
rect 11850 15206 11902 15258
rect 11914 15206 11966 15258
rect 11978 15206 12030 15258
rect 19658 15206 19710 15258
rect 19722 15206 19774 15258
rect 19786 15206 19838 15258
rect 19850 15206 19902 15258
rect 19914 15206 19966 15258
rect 19978 15206 20030 15258
rect 27658 15206 27710 15258
rect 27722 15206 27774 15258
rect 27786 15206 27838 15258
rect 27850 15206 27902 15258
rect 27914 15206 27966 15258
rect 27978 15206 28030 15258
rect 10784 15104 10836 15156
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 112 14900 164 14952
rect 11796 14968 11848 15020
rect 28080 15011 28132 15020
rect 28080 14977 28089 15011
rect 28089 14977 28123 15011
rect 28123 14977 28132 15011
rect 28080 14968 28132 14977
rect 10692 14900 10744 14952
rect 28356 14943 28408 14952
rect 28356 14909 28365 14943
rect 28365 14909 28399 14943
rect 28399 14909 28408 14943
rect 28356 14900 28408 14909
rect 11520 14832 11572 14884
rect 10784 14764 10836 14816
rect 12164 14764 12216 14816
rect 12808 14807 12860 14816
rect 12808 14773 12817 14807
rect 12817 14773 12851 14807
rect 12851 14773 12860 14807
rect 12808 14764 12860 14773
rect 2918 14662 2970 14714
rect 2982 14662 3034 14714
rect 3046 14662 3098 14714
rect 3110 14662 3162 14714
rect 3174 14662 3226 14714
rect 3238 14662 3290 14714
rect 10918 14662 10970 14714
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 11238 14662 11290 14714
rect 18918 14662 18970 14714
rect 18982 14662 19034 14714
rect 19046 14662 19098 14714
rect 19110 14662 19162 14714
rect 19174 14662 19226 14714
rect 19238 14662 19290 14714
rect 26918 14662 26970 14714
rect 26982 14662 27034 14714
rect 27046 14662 27098 14714
rect 27110 14662 27162 14714
rect 27174 14662 27226 14714
rect 27238 14662 27290 14714
rect 10784 14424 10836 14476
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 10692 14356 10744 14408
rect 11796 14356 11848 14408
rect 12716 14331 12768 14340
rect 12716 14297 12725 14331
rect 12725 14297 12759 14331
rect 12759 14297 12768 14331
rect 12716 14288 12768 14297
rect 12164 14220 12216 14272
rect 12440 14220 12492 14272
rect 28080 14220 28132 14272
rect 3658 14118 3710 14170
rect 3722 14118 3774 14170
rect 3786 14118 3838 14170
rect 3850 14118 3902 14170
rect 3914 14118 3966 14170
rect 3978 14118 4030 14170
rect 11658 14118 11710 14170
rect 11722 14118 11774 14170
rect 11786 14118 11838 14170
rect 11850 14118 11902 14170
rect 11914 14118 11966 14170
rect 11978 14118 12030 14170
rect 19658 14118 19710 14170
rect 19722 14118 19774 14170
rect 19786 14118 19838 14170
rect 19850 14118 19902 14170
rect 19914 14118 19966 14170
rect 19978 14118 20030 14170
rect 27658 14118 27710 14170
rect 27722 14118 27774 14170
rect 27786 14118 27838 14170
rect 27850 14118 27902 14170
rect 27914 14118 27966 14170
rect 27978 14118 28030 14170
rect 11520 14016 11572 14068
rect 12348 13880 12400 13932
rect 10324 13812 10376 13864
rect 28356 13855 28408 13864
rect 28356 13821 28365 13855
rect 28365 13821 28399 13855
rect 28399 13821 28408 13855
rect 28356 13812 28408 13821
rect 11520 13719 11572 13728
rect 11520 13685 11529 13719
rect 11529 13685 11563 13719
rect 11563 13685 11572 13719
rect 11520 13676 11572 13685
rect 2918 13574 2970 13626
rect 2982 13574 3034 13626
rect 3046 13574 3098 13626
rect 3110 13574 3162 13626
rect 3174 13574 3226 13626
rect 3238 13574 3290 13626
rect 10918 13574 10970 13626
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 11238 13574 11290 13626
rect 18918 13574 18970 13626
rect 18982 13574 19034 13626
rect 19046 13574 19098 13626
rect 19110 13574 19162 13626
rect 19174 13574 19226 13626
rect 19238 13574 19290 13626
rect 26918 13574 26970 13626
rect 26982 13574 27034 13626
rect 27046 13574 27098 13626
rect 27110 13574 27162 13626
rect 27174 13574 27226 13626
rect 27238 13574 27290 13626
rect 10784 13472 10836 13524
rect 12348 13472 12400 13524
rect 11520 13336 11572 13388
rect 12164 13336 12216 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 10692 13268 10744 13320
rect 13360 13268 13412 13320
rect 12348 13200 12400 13252
rect 28356 13243 28408 13252
rect 28356 13209 28365 13243
rect 28365 13209 28399 13243
rect 28399 13209 28408 13243
rect 28356 13200 28408 13209
rect 10876 13132 10928 13184
rect 12624 13132 12676 13184
rect 3658 13030 3710 13082
rect 3722 13030 3774 13082
rect 3786 13030 3838 13082
rect 3850 13030 3902 13082
rect 3914 13030 3966 13082
rect 3978 13030 4030 13082
rect 11658 13030 11710 13082
rect 11722 13030 11774 13082
rect 11786 13030 11838 13082
rect 11850 13030 11902 13082
rect 11914 13030 11966 13082
rect 11978 13030 12030 13082
rect 19658 13030 19710 13082
rect 19722 13030 19774 13082
rect 19786 13030 19838 13082
rect 19850 13030 19902 13082
rect 19914 13030 19966 13082
rect 19978 13030 20030 13082
rect 27658 13030 27710 13082
rect 27722 13030 27774 13082
rect 27786 13030 27838 13082
rect 27850 13030 27902 13082
rect 27914 13030 27966 13082
rect 27978 13030 28030 13082
rect 10876 12971 10928 12980
rect 10876 12937 10885 12971
rect 10885 12937 10919 12971
rect 10919 12937 10928 12971
rect 10876 12928 10928 12937
rect 13360 12928 13412 12980
rect 12440 12860 12492 12912
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 11980 12792 12032 12844
rect 10784 12767 10836 12776
rect 10784 12733 10793 12767
rect 10793 12733 10827 12767
rect 10827 12733 10836 12767
rect 10784 12724 10836 12733
rect 12624 12724 12676 12776
rect 10600 12588 10652 12640
rect 10692 12588 10744 12640
rect 11336 12631 11388 12640
rect 11336 12597 11345 12631
rect 11345 12597 11379 12631
rect 11379 12597 11388 12631
rect 11336 12588 11388 12597
rect 2918 12486 2970 12538
rect 2982 12486 3034 12538
rect 3046 12486 3098 12538
rect 3110 12486 3162 12538
rect 3174 12486 3226 12538
rect 3238 12486 3290 12538
rect 10918 12486 10970 12538
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 11238 12486 11290 12538
rect 18918 12486 18970 12538
rect 18982 12486 19034 12538
rect 19046 12486 19098 12538
rect 19110 12486 19162 12538
rect 19174 12486 19226 12538
rect 19238 12486 19290 12538
rect 26918 12486 26970 12538
rect 26982 12486 27034 12538
rect 27046 12486 27098 12538
rect 27110 12486 27162 12538
rect 27174 12486 27226 12538
rect 27238 12486 27290 12538
rect 11336 12248 11388 12300
rect 10692 12223 10744 12232
rect 10692 12189 10701 12223
rect 10701 12189 10735 12223
rect 10735 12189 10744 12223
rect 10692 12180 10744 12189
rect 11980 12180 12032 12232
rect 12348 12112 12400 12164
rect 28356 12155 28408 12164
rect 28356 12121 28365 12155
rect 28365 12121 28399 12155
rect 28399 12121 28408 12155
rect 28356 12112 28408 12121
rect 3658 11942 3710 11994
rect 3722 11942 3774 11994
rect 3786 11942 3838 11994
rect 3850 11942 3902 11994
rect 3914 11942 3966 11994
rect 3978 11942 4030 11994
rect 11658 11942 11710 11994
rect 11722 11942 11774 11994
rect 11786 11942 11838 11994
rect 11850 11942 11902 11994
rect 11914 11942 11966 11994
rect 11978 11942 12030 11994
rect 19658 11942 19710 11994
rect 19722 11942 19774 11994
rect 19786 11942 19838 11994
rect 19850 11942 19902 11994
rect 19914 11942 19966 11994
rect 19978 11942 20030 11994
rect 27658 11942 27710 11994
rect 27722 11942 27774 11994
rect 27786 11942 27838 11994
rect 27850 11942 27902 11994
rect 27914 11942 27966 11994
rect 27978 11942 28030 11994
rect 12440 11772 12492 11824
rect 1400 11747 1452 11756
rect 1400 11713 1409 11747
rect 1409 11713 1443 11747
rect 1443 11713 1452 11747
rect 1400 11704 1452 11713
rect 10692 11636 10744 11688
rect 11704 11636 11756 11688
rect 12808 11636 12860 11688
rect 11428 11568 11480 11620
rect 11336 11500 11388 11552
rect 28356 11679 28408 11688
rect 28356 11645 28365 11679
rect 28365 11645 28399 11679
rect 28399 11645 28408 11679
rect 28356 11636 28408 11645
rect 2918 11398 2970 11450
rect 2982 11398 3034 11450
rect 3046 11398 3098 11450
rect 3110 11398 3162 11450
rect 3174 11398 3226 11450
rect 3238 11398 3290 11450
rect 10918 11398 10970 11450
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 11238 11398 11290 11450
rect 18918 11398 18970 11450
rect 18982 11398 19034 11450
rect 19046 11398 19098 11450
rect 19110 11398 19162 11450
rect 19174 11398 19226 11450
rect 19238 11398 19290 11450
rect 26918 11398 26970 11450
rect 26982 11398 27034 11450
rect 27046 11398 27098 11450
rect 27110 11398 27162 11450
rect 27174 11398 27226 11450
rect 27238 11398 27290 11450
rect 11244 11160 11296 11212
rect 11428 11160 11480 11212
rect 12072 11160 12124 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 10692 11135 10744 11144
rect 10692 11101 10701 11135
rect 10701 11101 10735 11135
rect 10735 11101 10744 11135
rect 10692 11092 10744 11101
rect 11060 11135 11112 11144
rect 11060 11101 11069 11135
rect 11069 11101 11103 11135
rect 11103 11101 11112 11135
rect 11060 11092 11112 11101
rect 12348 11024 12400 11076
rect 12440 11024 12492 11076
rect 3658 10854 3710 10906
rect 3722 10854 3774 10906
rect 3786 10854 3838 10906
rect 3850 10854 3902 10906
rect 3914 10854 3966 10906
rect 3978 10854 4030 10906
rect 11658 10854 11710 10906
rect 11722 10854 11774 10906
rect 11786 10854 11838 10906
rect 11850 10854 11902 10906
rect 11914 10854 11966 10906
rect 11978 10854 12030 10906
rect 19658 10854 19710 10906
rect 19722 10854 19774 10906
rect 19786 10854 19838 10906
rect 19850 10854 19902 10906
rect 19914 10854 19966 10906
rect 19978 10854 20030 10906
rect 27658 10854 27710 10906
rect 27722 10854 27774 10906
rect 27786 10854 27838 10906
rect 27850 10854 27902 10906
rect 27914 10854 27966 10906
rect 27978 10854 28030 10906
rect 10600 10752 10652 10804
rect 11060 10752 11112 10804
rect 12072 10752 12124 10804
rect 10324 10727 10376 10736
rect 10324 10693 10333 10727
rect 10333 10693 10367 10727
rect 10367 10693 10376 10727
rect 10324 10684 10376 10693
rect 11336 10684 11388 10736
rect 11428 10616 11480 10668
rect 12440 10616 12492 10668
rect 10784 10591 10836 10600
rect 10784 10557 10793 10591
rect 10793 10557 10827 10591
rect 10827 10557 10836 10591
rect 10784 10548 10836 10557
rect 13176 10548 13228 10600
rect 28356 10591 28408 10600
rect 28356 10557 28365 10591
rect 28365 10557 28399 10591
rect 28399 10557 28408 10591
rect 28356 10548 28408 10557
rect 11520 10480 11572 10532
rect 12072 10412 12124 10464
rect 12256 10412 12308 10464
rect 2918 10310 2970 10362
rect 2982 10310 3034 10362
rect 3046 10310 3098 10362
rect 3110 10310 3162 10362
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 10918 10310 10970 10362
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 11238 10310 11290 10362
rect 18918 10310 18970 10362
rect 18982 10310 19034 10362
rect 19046 10310 19098 10362
rect 19110 10310 19162 10362
rect 19174 10310 19226 10362
rect 19238 10310 19290 10362
rect 26918 10310 26970 10362
rect 26982 10310 27034 10362
rect 27046 10310 27098 10362
rect 27110 10310 27162 10362
rect 27174 10310 27226 10362
rect 27238 10310 27290 10362
rect 13176 10115 13228 10124
rect 13176 10081 13185 10115
rect 13185 10081 13219 10115
rect 13219 10081 13228 10115
rect 13176 10072 13228 10081
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 12348 9936 12400 9988
rect 28356 9979 28408 9988
rect 28356 9945 28365 9979
rect 28365 9945 28399 9979
rect 28399 9945 28408 9979
rect 28356 9936 28408 9945
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 11336 9868 11388 9920
rect 3658 9766 3710 9818
rect 3722 9766 3774 9818
rect 3786 9766 3838 9818
rect 3850 9766 3902 9818
rect 3914 9766 3966 9818
rect 3978 9766 4030 9818
rect 11658 9766 11710 9818
rect 11722 9766 11774 9818
rect 11786 9766 11838 9818
rect 11850 9766 11902 9818
rect 11914 9766 11966 9818
rect 11978 9766 12030 9818
rect 19658 9766 19710 9818
rect 19722 9766 19774 9818
rect 19786 9766 19838 9818
rect 19850 9766 19902 9818
rect 19914 9766 19966 9818
rect 19978 9766 20030 9818
rect 27658 9766 27710 9818
rect 27722 9766 27774 9818
rect 27786 9766 27838 9818
rect 27850 9766 27902 9818
rect 27914 9766 27966 9818
rect 27978 9766 28030 9818
rect 1584 9664 1636 9716
rect 10692 9596 10744 9648
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 12256 9596 12308 9648
rect 10784 9503 10836 9512
rect 10784 9469 10793 9503
rect 10793 9469 10827 9503
rect 10827 9469 10836 9503
rect 10784 9460 10836 9469
rect 10784 9324 10836 9376
rect 28080 9324 28132 9376
rect 2918 9222 2970 9274
rect 2982 9222 3034 9274
rect 3046 9222 3098 9274
rect 3110 9222 3162 9274
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 10918 9222 10970 9274
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 11238 9222 11290 9274
rect 18918 9222 18970 9274
rect 18982 9222 19034 9274
rect 19046 9222 19098 9274
rect 19110 9222 19162 9274
rect 19174 9222 19226 9274
rect 19238 9222 19290 9274
rect 26918 9222 26970 9274
rect 26982 9222 27034 9274
rect 27046 9222 27098 9274
rect 27110 9222 27162 9274
rect 27174 9222 27226 9274
rect 27238 9222 27290 9274
rect 12256 9120 12308 9172
rect 12072 8916 12124 8968
rect 28080 8959 28132 8968
rect 28080 8925 28089 8959
rect 28089 8925 28123 8959
rect 28123 8925 28132 8959
rect 28080 8916 28132 8925
rect 28356 8891 28408 8900
rect 28356 8857 28365 8891
rect 28365 8857 28399 8891
rect 28399 8857 28408 8891
rect 28356 8848 28408 8857
rect 3658 8678 3710 8730
rect 3722 8678 3774 8730
rect 3786 8678 3838 8730
rect 3850 8678 3902 8730
rect 3914 8678 3966 8730
rect 3978 8678 4030 8730
rect 11658 8678 11710 8730
rect 11722 8678 11774 8730
rect 11786 8678 11838 8730
rect 11850 8678 11902 8730
rect 11914 8678 11966 8730
rect 11978 8678 12030 8730
rect 19658 8678 19710 8730
rect 19722 8678 19774 8730
rect 19786 8678 19838 8730
rect 19850 8678 19902 8730
rect 19914 8678 19966 8730
rect 19978 8678 20030 8730
rect 27658 8678 27710 8730
rect 27722 8678 27774 8730
rect 27786 8678 27838 8730
rect 27850 8678 27902 8730
rect 27914 8678 27966 8730
rect 27978 8678 28030 8730
rect 10784 8576 10836 8628
rect 12072 8508 12124 8560
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 11336 8440 11388 8492
rect 11428 8372 11480 8424
rect 10692 8236 10744 8288
rect 28356 8415 28408 8424
rect 28356 8381 28365 8415
rect 28365 8381 28399 8415
rect 28399 8381 28408 8415
rect 28356 8372 28408 8381
rect 2918 8134 2970 8186
rect 2982 8134 3034 8186
rect 3046 8134 3098 8186
rect 3110 8134 3162 8186
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 10918 8134 10970 8186
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 11238 8134 11290 8186
rect 18918 8134 18970 8186
rect 18982 8134 19034 8186
rect 19046 8134 19098 8186
rect 19110 8134 19162 8186
rect 19174 8134 19226 8186
rect 19238 8134 19290 8186
rect 26918 8134 26970 8186
rect 26982 8134 27034 8186
rect 27046 8134 27098 8186
rect 27110 8134 27162 8186
rect 27174 8134 27226 8186
rect 27238 8134 27290 8186
rect 10692 7939 10744 7948
rect 10692 7905 10701 7939
rect 10701 7905 10735 7939
rect 10735 7905 10744 7939
rect 10692 7896 10744 7905
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 12072 7828 12124 7880
rect 12348 7828 12400 7880
rect 10968 7803 11020 7812
rect 10968 7769 10977 7803
rect 10977 7769 11011 7803
rect 11011 7769 11020 7803
rect 10968 7760 11020 7769
rect 10140 7692 10192 7744
rect 12440 7735 12492 7744
rect 12440 7701 12449 7735
rect 12449 7701 12483 7735
rect 12483 7701 12492 7735
rect 12440 7692 12492 7701
rect 28080 7692 28132 7744
rect 3658 7590 3710 7642
rect 3722 7590 3774 7642
rect 3786 7590 3838 7642
rect 3850 7590 3902 7642
rect 3914 7590 3966 7642
rect 3978 7590 4030 7642
rect 11658 7590 11710 7642
rect 11722 7590 11774 7642
rect 11786 7590 11838 7642
rect 11850 7590 11902 7642
rect 11914 7590 11966 7642
rect 11978 7590 12030 7642
rect 19658 7590 19710 7642
rect 19722 7590 19774 7642
rect 19786 7590 19838 7642
rect 19850 7590 19902 7642
rect 19914 7590 19966 7642
rect 19978 7590 20030 7642
rect 27658 7590 27710 7642
rect 27722 7590 27774 7642
rect 27786 7590 27838 7642
rect 27850 7590 27902 7642
rect 27914 7590 27966 7642
rect 27978 7590 28030 7642
rect 10968 7488 11020 7540
rect 12440 7488 12492 7540
rect 11336 7420 11388 7472
rect 28080 7395 28132 7404
rect 28080 7361 28089 7395
rect 28089 7361 28123 7395
rect 28123 7361 28132 7395
rect 28080 7352 28132 7361
rect 11428 7284 11480 7336
rect 28356 7327 28408 7336
rect 28356 7293 28365 7327
rect 28365 7293 28399 7327
rect 28399 7293 28408 7327
rect 28356 7284 28408 7293
rect 2918 7046 2970 7098
rect 2982 7046 3034 7098
rect 3046 7046 3098 7098
rect 3110 7046 3162 7098
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 10918 7046 10970 7098
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 11238 7046 11290 7098
rect 18918 7046 18970 7098
rect 18982 7046 19034 7098
rect 19046 7046 19098 7098
rect 19110 7046 19162 7098
rect 19174 7046 19226 7098
rect 19238 7046 19290 7098
rect 26918 7046 26970 7098
rect 26982 7046 27034 7098
rect 27046 7046 27098 7098
rect 27110 7046 27162 7098
rect 27174 7046 27226 7098
rect 27238 7046 27290 7098
rect 10692 6808 10744 6860
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 12808 6783 12860 6792
rect 12808 6749 12817 6783
rect 12817 6749 12851 6783
rect 12851 6749 12860 6783
rect 12808 6740 12860 6749
rect 28080 6783 28132 6792
rect 28080 6749 28089 6783
rect 28089 6749 28123 6783
rect 28123 6749 28132 6783
rect 28080 6740 28132 6749
rect 28356 6715 28408 6724
rect 28356 6681 28365 6715
rect 28365 6681 28399 6715
rect 28399 6681 28408 6715
rect 28356 6672 28408 6681
rect 10048 6604 10100 6656
rect 3658 6502 3710 6554
rect 3722 6502 3774 6554
rect 3786 6502 3838 6554
rect 3850 6502 3902 6554
rect 3914 6502 3966 6554
rect 3978 6502 4030 6554
rect 11658 6502 11710 6554
rect 11722 6502 11774 6554
rect 11786 6502 11838 6554
rect 11850 6502 11902 6554
rect 11914 6502 11966 6554
rect 11978 6502 12030 6554
rect 19658 6502 19710 6554
rect 19722 6502 19774 6554
rect 19786 6502 19838 6554
rect 19850 6502 19902 6554
rect 19914 6502 19966 6554
rect 19978 6502 20030 6554
rect 27658 6502 27710 6554
rect 27722 6502 27774 6554
rect 27786 6502 27838 6554
rect 27850 6502 27902 6554
rect 27914 6502 27966 6554
rect 27978 6502 28030 6554
rect 10048 6443 10100 6452
rect 10048 6409 10057 6443
rect 10057 6409 10091 6443
rect 10091 6409 10100 6443
rect 10048 6400 10100 6409
rect 10140 6400 10192 6452
rect 10692 6332 10744 6384
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 10140 6307 10192 6316
rect 10140 6273 10149 6307
rect 10149 6273 10183 6307
rect 10183 6273 10192 6307
rect 10140 6264 10192 6273
rect 12256 6332 12308 6384
rect 10784 6196 10836 6248
rect 10416 6128 10468 6180
rect 10508 6103 10560 6112
rect 10508 6069 10517 6103
rect 10517 6069 10551 6103
rect 10551 6069 10560 6103
rect 10508 6060 10560 6069
rect 28080 6060 28132 6112
rect 2918 5958 2970 6010
rect 2982 5958 3034 6010
rect 3046 5958 3098 6010
rect 3110 5958 3162 6010
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 10918 5958 10970 6010
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 11238 5958 11290 6010
rect 18918 5958 18970 6010
rect 18982 5958 19034 6010
rect 19046 5958 19098 6010
rect 19110 5958 19162 6010
rect 19174 5958 19226 6010
rect 19238 5958 19290 6010
rect 26918 5958 26970 6010
rect 26982 5958 27034 6010
rect 27046 5958 27098 6010
rect 27110 5958 27162 6010
rect 27174 5958 27226 6010
rect 27238 5958 27290 6010
rect 10140 5856 10192 5908
rect 10508 5788 10560 5840
rect 10692 5763 10744 5772
rect 10692 5729 10701 5763
rect 10701 5729 10735 5763
rect 10735 5729 10744 5763
rect 10692 5720 10744 5729
rect 12256 5584 12308 5636
rect 28356 5627 28408 5636
rect 28356 5593 28365 5627
rect 28365 5593 28399 5627
rect 28399 5593 28408 5627
rect 28356 5584 28408 5593
rect 3658 5414 3710 5466
rect 3722 5414 3774 5466
rect 3786 5414 3838 5466
rect 3850 5414 3902 5466
rect 3914 5414 3966 5466
rect 3978 5414 4030 5466
rect 11658 5414 11710 5466
rect 11722 5414 11774 5466
rect 11786 5414 11838 5466
rect 11850 5414 11902 5466
rect 11914 5414 11966 5466
rect 11978 5414 12030 5466
rect 19658 5414 19710 5466
rect 19722 5414 19774 5466
rect 19786 5414 19838 5466
rect 19850 5414 19902 5466
rect 19914 5414 19966 5466
rect 19978 5414 20030 5466
rect 27658 5414 27710 5466
rect 27722 5414 27774 5466
rect 27786 5414 27838 5466
rect 27850 5414 27902 5466
rect 27914 5414 27966 5466
rect 27978 5414 28030 5466
rect 10416 5312 10468 5364
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 12532 5176 12584 5228
rect 28080 5219 28132 5228
rect 28080 5185 28089 5219
rect 28089 5185 28123 5219
rect 28123 5185 28132 5219
rect 28080 5176 28132 5185
rect 10784 5108 10836 5160
rect 12992 5108 13044 5160
rect 28356 5151 28408 5160
rect 28356 5117 28365 5151
rect 28365 5117 28399 5151
rect 28399 5117 28408 5151
rect 28356 5108 28408 5117
rect 7564 4972 7616 5024
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 2918 4870 2970 4922
rect 2982 4870 3034 4922
rect 3046 4870 3098 4922
rect 3110 4870 3162 4922
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 10918 4870 10970 4922
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 11238 4870 11290 4922
rect 18918 4870 18970 4922
rect 18982 4870 19034 4922
rect 19046 4870 19098 4922
rect 19110 4870 19162 4922
rect 19174 4870 19226 4922
rect 19238 4870 19290 4922
rect 26918 4870 26970 4922
rect 26982 4870 27034 4922
rect 27046 4870 27098 4922
rect 27110 4870 27162 4922
rect 27174 4870 27226 4922
rect 27238 4870 27290 4922
rect 7564 4768 7616 4820
rect 10600 4675 10652 4684
rect 10600 4641 10609 4675
rect 10609 4641 10643 4675
rect 10643 4641 10652 4675
rect 10600 4632 10652 4641
rect 11520 4632 11572 4684
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 12256 4632 12308 4684
rect 12992 4675 13044 4684
rect 12992 4641 13001 4675
rect 13001 4641 13035 4675
rect 13035 4641 13044 4675
rect 12992 4632 13044 4641
rect 12716 4564 12768 4616
rect 12532 4496 12584 4548
rect 12440 4471 12492 4480
rect 12440 4437 12449 4471
rect 12449 4437 12483 4471
rect 12483 4437 12492 4471
rect 12440 4428 12492 4437
rect 12808 4471 12860 4480
rect 12808 4437 12817 4471
rect 12817 4437 12851 4471
rect 12851 4437 12860 4471
rect 12808 4428 12860 4437
rect 3658 4326 3710 4378
rect 3722 4326 3774 4378
rect 3786 4326 3838 4378
rect 3850 4326 3902 4378
rect 3914 4326 3966 4378
rect 3978 4326 4030 4378
rect 11658 4326 11710 4378
rect 11722 4326 11774 4378
rect 11786 4326 11838 4378
rect 11850 4326 11902 4378
rect 11914 4326 11966 4378
rect 11978 4326 12030 4378
rect 19658 4326 19710 4378
rect 19722 4326 19774 4378
rect 19786 4326 19838 4378
rect 19850 4326 19902 4378
rect 19914 4326 19966 4378
rect 19978 4326 20030 4378
rect 27658 4326 27710 4378
rect 27722 4326 27774 4378
rect 27786 4326 27838 4378
rect 27850 4326 27902 4378
rect 27914 4326 27966 4378
rect 27978 4326 28030 4378
rect 12532 4224 12584 4276
rect 28080 4224 28132 4276
rect 11520 4156 11572 4208
rect 12256 4156 12308 4208
rect 11428 4088 11480 4140
rect 10600 4020 10652 4072
rect 12440 4020 12492 4072
rect 12808 4020 12860 4072
rect 28356 4063 28408 4072
rect 28356 4029 28365 4063
rect 28365 4029 28399 4063
rect 28399 4029 28408 4063
rect 28356 4020 28408 4029
rect 2918 3782 2970 3834
rect 2982 3782 3034 3834
rect 3046 3782 3098 3834
rect 3110 3782 3162 3834
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 10918 3782 10970 3834
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 11238 3782 11290 3834
rect 18918 3782 18970 3834
rect 18982 3782 19034 3834
rect 19046 3782 19098 3834
rect 19110 3782 19162 3834
rect 19174 3782 19226 3834
rect 19238 3782 19290 3834
rect 26918 3782 26970 3834
rect 26982 3782 27034 3834
rect 27046 3782 27098 3834
rect 27110 3782 27162 3834
rect 27174 3782 27226 3834
rect 27238 3782 27290 3834
rect 10692 3680 10744 3732
rect 10600 3587 10652 3596
rect 10600 3553 10609 3587
rect 10609 3553 10643 3587
rect 10643 3553 10652 3587
rect 10600 3544 10652 3553
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 12716 3544 12768 3596
rect 12992 3587 13044 3596
rect 12992 3553 13001 3587
rect 13001 3553 13035 3587
rect 13035 3553 13044 3587
rect 12992 3544 13044 3553
rect 11152 3408 11204 3460
rect 12256 3408 12308 3460
rect 12348 3408 12400 3460
rect 10232 3340 10284 3392
rect 12164 3340 12216 3392
rect 28356 3451 28408 3460
rect 28356 3417 28365 3451
rect 28365 3417 28399 3451
rect 28399 3417 28408 3451
rect 28356 3408 28408 3417
rect 3658 3238 3710 3290
rect 3722 3238 3774 3290
rect 3786 3238 3838 3290
rect 3850 3238 3902 3290
rect 3914 3238 3966 3290
rect 3978 3238 4030 3290
rect 11658 3238 11710 3290
rect 11722 3238 11774 3290
rect 11786 3238 11838 3290
rect 11850 3238 11902 3290
rect 11914 3238 11966 3290
rect 11978 3238 12030 3290
rect 19658 3238 19710 3290
rect 19722 3238 19774 3290
rect 19786 3238 19838 3290
rect 19850 3238 19902 3290
rect 19914 3238 19966 3290
rect 19978 3238 20030 3290
rect 27658 3238 27710 3290
rect 27722 3238 27774 3290
rect 27786 3238 27838 3290
rect 27850 3238 27902 3290
rect 27914 3238 27966 3290
rect 27978 3238 28030 3290
rect 10232 3136 10284 3188
rect 11060 3136 11112 3188
rect 11520 3136 11572 3188
rect 10600 3068 10652 3120
rect 848 3000 900 3052
rect 12256 3068 12308 3120
rect 10692 2975 10744 2984
rect 10692 2941 10701 2975
rect 10701 2941 10735 2975
rect 10735 2941 10744 2975
rect 10692 2932 10744 2941
rect 10876 2796 10928 2848
rect 20628 2796 20680 2848
rect 2918 2694 2970 2746
rect 2982 2694 3034 2746
rect 3046 2694 3098 2746
rect 3110 2694 3162 2746
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 10918 2694 10970 2746
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 11238 2694 11290 2746
rect 18918 2694 18970 2746
rect 18982 2694 19034 2746
rect 19046 2694 19098 2746
rect 19110 2694 19162 2746
rect 19174 2694 19226 2746
rect 19238 2694 19290 2746
rect 26918 2694 26970 2746
rect 26982 2694 27034 2746
rect 27046 2694 27098 2746
rect 27110 2694 27162 2746
rect 27174 2694 27226 2746
rect 27238 2694 27290 2746
rect 12256 2592 12308 2644
rect 848 2388 900 2440
rect 12348 2388 12400 2440
rect 20628 2388 20680 2440
rect 28356 2363 28408 2372
rect 28356 2329 28365 2363
rect 28365 2329 28399 2363
rect 28399 2329 28408 2363
rect 28356 2320 28408 2329
rect 12164 2252 12216 2304
rect 3658 2150 3710 2202
rect 3722 2150 3774 2202
rect 3786 2150 3838 2202
rect 3850 2150 3902 2202
rect 3914 2150 3966 2202
rect 3978 2150 4030 2202
rect 11658 2150 11710 2202
rect 11722 2150 11774 2202
rect 11786 2150 11838 2202
rect 11850 2150 11902 2202
rect 11914 2150 11966 2202
rect 11978 2150 12030 2202
rect 19658 2150 19710 2202
rect 19722 2150 19774 2202
rect 19786 2150 19838 2202
rect 19850 2150 19902 2202
rect 19914 2150 19966 2202
rect 19978 2150 20030 2202
rect 27658 2150 27710 2202
rect 27722 2150 27774 2202
rect 27786 2150 27838 2202
rect 27850 2150 27902 2202
rect 27914 2150 27966 2202
rect 27978 2150 28030 2202
<< metal2 >>
rect 1030 28656 1086 28665
rect 1030 28591 1086 28600
rect 938 27840 994 27849
rect 938 27775 994 27784
rect 952 27538 980 27775
rect 1044 27606 1072 28591
rect 2916 27772 3292 27781
rect 2972 27770 2996 27772
rect 3052 27770 3076 27772
rect 3132 27770 3156 27772
rect 3212 27770 3236 27772
rect 2972 27718 2982 27770
rect 3226 27718 3236 27770
rect 2972 27716 2996 27718
rect 3052 27716 3076 27718
rect 3132 27716 3156 27718
rect 3212 27716 3236 27718
rect 2916 27707 3292 27716
rect 10916 27772 11292 27781
rect 10972 27770 10996 27772
rect 11052 27770 11076 27772
rect 11132 27770 11156 27772
rect 11212 27770 11236 27772
rect 10972 27718 10982 27770
rect 11226 27718 11236 27770
rect 10972 27716 10996 27718
rect 11052 27716 11076 27718
rect 11132 27716 11156 27718
rect 11212 27716 11236 27718
rect 10916 27707 11292 27716
rect 18916 27772 19292 27781
rect 18972 27770 18996 27772
rect 19052 27770 19076 27772
rect 19132 27770 19156 27772
rect 19212 27770 19236 27772
rect 18972 27718 18982 27770
rect 19226 27718 19236 27770
rect 18972 27716 18996 27718
rect 19052 27716 19076 27718
rect 19132 27716 19156 27718
rect 19212 27716 19236 27718
rect 18916 27707 19292 27716
rect 26916 27772 27292 27781
rect 26972 27770 26996 27772
rect 27052 27770 27076 27772
rect 27132 27770 27156 27772
rect 27212 27770 27236 27772
rect 26972 27718 26982 27770
rect 27226 27718 27236 27770
rect 26972 27716 26996 27718
rect 27052 27716 27076 27718
rect 27132 27716 27156 27718
rect 27212 27716 27236 27718
rect 26916 27707 27292 27716
rect 1032 27600 1084 27606
rect 1032 27542 1084 27548
rect 10968 27600 11020 27606
rect 10968 27542 11020 27548
rect 28354 27568 28410 27577
rect 940 27532 992 27538
rect 940 27474 992 27480
rect 848 27464 900 27470
rect 848 27406 900 27412
rect 860 27169 888 27406
rect 1584 27328 1636 27334
rect 1584 27270 1636 27276
rect 846 27160 902 27169
rect 1596 27130 1624 27270
rect 3656 27228 4032 27237
rect 3712 27226 3736 27228
rect 3792 27226 3816 27228
rect 3872 27226 3896 27228
rect 3952 27226 3976 27228
rect 3712 27174 3722 27226
rect 3966 27174 3976 27226
rect 3712 27172 3736 27174
rect 3792 27172 3816 27174
rect 3872 27172 3896 27174
rect 3952 27172 3976 27174
rect 3656 27163 4032 27172
rect 10980 27130 11008 27542
rect 28354 27503 28356 27512
rect 28408 27503 28410 27512
rect 28356 27474 28408 27480
rect 12348 27464 12400 27470
rect 12348 27406 12400 27412
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 11428 27396 11480 27402
rect 11428 27338 11480 27344
rect 11440 27130 11468 27338
rect 12164 27328 12216 27334
rect 12164 27270 12216 27276
rect 11656 27228 12032 27237
rect 11712 27226 11736 27228
rect 11792 27226 11816 27228
rect 11872 27226 11896 27228
rect 11952 27226 11976 27228
rect 11712 27174 11722 27226
rect 11966 27174 11976 27226
rect 11712 27172 11736 27174
rect 11792 27172 11816 27174
rect 11872 27172 11896 27174
rect 11952 27172 11976 27174
rect 11656 27163 12032 27172
rect 846 27095 902 27104
rect 1584 27124 1636 27130
rect 1584 27066 1636 27072
rect 10968 27124 11020 27130
rect 10968 27066 11020 27072
rect 11428 27124 11480 27130
rect 11428 27066 11480 27072
rect 12176 26926 12204 27270
rect 12256 26988 12308 26994
rect 12256 26930 12308 26936
rect 12164 26920 12216 26926
rect 12164 26862 12216 26868
rect 9220 26852 9272 26858
rect 9220 26794 9272 26800
rect 2916 26684 3292 26693
rect 2972 26682 2996 26684
rect 3052 26682 3076 26684
rect 3132 26682 3156 26684
rect 3212 26682 3236 26684
rect 2972 26630 2982 26682
rect 3226 26630 3236 26682
rect 2972 26628 2996 26630
rect 3052 26628 3076 26630
rect 3132 26628 3156 26630
rect 3212 26628 3236 26630
rect 2916 26619 3292 26628
rect 9232 26586 9260 26794
rect 10600 26784 10652 26790
rect 10600 26726 10652 26732
rect 11428 26784 11480 26790
rect 11428 26726 11480 26732
rect 12072 26784 12124 26790
rect 12072 26726 12124 26732
rect 9220 26580 9272 26586
rect 9220 26522 9272 26528
rect 10612 26450 10640 26726
rect 10916 26684 11292 26693
rect 10972 26682 10996 26684
rect 11052 26682 11076 26684
rect 11132 26682 11156 26684
rect 11212 26682 11236 26684
rect 10972 26630 10982 26682
rect 11226 26630 11236 26682
rect 10972 26628 10996 26630
rect 11052 26628 11076 26630
rect 11132 26628 11156 26630
rect 11212 26628 11236 26630
rect 10916 26619 11292 26628
rect 11440 26450 11468 26726
rect 10416 26444 10468 26450
rect 10416 26386 10468 26392
rect 10600 26444 10652 26450
rect 10600 26386 10652 26392
rect 11428 26444 11480 26450
rect 11428 26386 11480 26392
rect 848 26376 900 26382
rect 848 26318 900 26324
rect 860 26081 888 26318
rect 3656 26140 4032 26149
rect 3712 26138 3736 26140
rect 3792 26138 3816 26140
rect 3872 26138 3896 26140
rect 3952 26138 3976 26140
rect 3712 26086 3722 26138
rect 3966 26086 3976 26138
rect 3712 26084 3736 26086
rect 3792 26084 3816 26086
rect 3872 26084 3896 26086
rect 3952 26084 3976 26086
rect 846 26072 902 26081
rect 3656 26075 4032 26084
rect 10428 26042 10456 26386
rect 11336 26376 11388 26382
rect 11336 26318 11388 26324
rect 846 26007 902 26016
rect 10416 26036 10468 26042
rect 10416 25978 10468 25984
rect 848 25900 900 25906
rect 848 25842 900 25848
rect 860 25537 888 25842
rect 11348 25838 11376 26318
rect 12084 26246 12112 26726
rect 12176 26450 12204 26862
rect 12164 26444 12216 26450
rect 12164 26386 12216 26392
rect 12268 26382 12296 26930
rect 12256 26376 12308 26382
rect 12256 26318 12308 26324
rect 12072 26240 12124 26246
rect 12072 26182 12124 26188
rect 11656 26140 12032 26149
rect 11712 26138 11736 26140
rect 11792 26138 11816 26140
rect 11872 26138 11896 26140
rect 11952 26138 11976 26140
rect 11712 26086 11722 26138
rect 11966 26086 11976 26138
rect 11712 26084 11736 26086
rect 11792 26084 11816 26086
rect 11872 26084 11896 26086
rect 11952 26084 11976 26086
rect 11656 26075 12032 26084
rect 12084 26042 12112 26182
rect 12072 26036 12124 26042
rect 12072 25978 12124 25984
rect 11612 25900 11664 25906
rect 11612 25842 11664 25848
rect 11336 25832 11388 25838
rect 11336 25774 11388 25780
rect 10600 25696 10652 25702
rect 10600 25638 10652 25644
rect 2916 25596 3292 25605
rect 2972 25594 2996 25596
rect 3052 25594 3076 25596
rect 3132 25594 3156 25596
rect 3212 25594 3236 25596
rect 2972 25542 2982 25594
rect 3226 25542 3236 25594
rect 2972 25540 2996 25542
rect 3052 25540 3076 25542
rect 3132 25540 3156 25542
rect 3212 25540 3236 25542
rect 846 25528 902 25537
rect 2916 25531 3292 25540
rect 846 25463 902 25472
rect 3656 25052 4032 25061
rect 3712 25050 3736 25052
rect 3792 25050 3816 25052
rect 3872 25050 3896 25052
rect 3952 25050 3976 25052
rect 3712 24998 3722 25050
rect 3966 24998 3976 25050
rect 3712 24996 3736 24998
rect 3792 24996 3816 24998
rect 3872 24996 3896 24998
rect 3952 24996 3976 24998
rect 3656 24987 4032 24996
rect 848 24812 900 24818
rect 848 24754 900 24760
rect 860 24721 888 24754
rect 846 24712 902 24721
rect 846 24647 902 24656
rect 2916 24508 3292 24517
rect 2972 24506 2996 24508
rect 3052 24506 3076 24508
rect 3132 24506 3156 24508
rect 3212 24506 3236 24508
rect 2972 24454 2982 24506
rect 3226 24454 3236 24506
rect 2972 24452 2996 24454
rect 3052 24452 3076 24454
rect 3132 24452 3156 24454
rect 3212 24452 3236 24454
rect 2916 24443 3292 24452
rect 10612 24274 10640 25638
rect 10916 25596 11292 25605
rect 10972 25594 10996 25596
rect 11052 25594 11076 25596
rect 11132 25594 11156 25596
rect 11212 25594 11236 25596
rect 10972 25542 10982 25594
rect 11226 25542 11236 25594
rect 10972 25540 10996 25542
rect 11052 25540 11076 25542
rect 11132 25540 11156 25542
rect 11212 25540 11236 25542
rect 10916 25531 11292 25540
rect 11348 25294 11376 25774
rect 11428 25696 11480 25702
rect 11428 25638 11480 25644
rect 11440 25362 11468 25638
rect 11624 25362 11652 25842
rect 12072 25696 12124 25702
rect 12072 25638 12124 25644
rect 11428 25356 11480 25362
rect 11428 25298 11480 25304
rect 11612 25356 11664 25362
rect 11612 25298 11664 25304
rect 11336 25288 11388 25294
rect 11336 25230 11388 25236
rect 11348 24750 11376 25230
rect 11656 25052 12032 25061
rect 11712 25050 11736 25052
rect 11792 25050 11816 25052
rect 11872 25050 11896 25052
rect 11952 25050 11976 25052
rect 11712 24998 11722 25050
rect 11966 24998 11976 25050
rect 11712 24996 11736 24998
rect 11792 24996 11816 24998
rect 11872 24996 11896 24998
rect 11952 24996 11976 24998
rect 11656 24987 12032 24996
rect 11336 24744 11388 24750
rect 11336 24686 11388 24692
rect 10916 24508 11292 24517
rect 10972 24506 10996 24508
rect 11052 24506 11076 24508
rect 11132 24506 11156 24508
rect 11212 24506 11236 24508
rect 10972 24454 10982 24506
rect 11226 24454 11236 24506
rect 10972 24452 10996 24454
rect 11052 24452 11076 24454
rect 11132 24452 11156 24454
rect 11212 24452 11236 24454
rect 10916 24443 11292 24452
rect 10600 24268 10652 24274
rect 10600 24210 10652 24216
rect 11348 24206 11376 24686
rect 11428 24608 11480 24614
rect 11428 24550 11480 24556
rect 848 24200 900 24206
rect 848 24142 900 24148
rect 11336 24200 11388 24206
rect 11336 24142 11388 24148
rect 860 23905 888 24142
rect 1584 24064 1636 24070
rect 1584 24006 1636 24012
rect 846 23896 902 23905
rect 1596 23866 1624 24006
rect 3656 23964 4032 23973
rect 3712 23962 3736 23964
rect 3792 23962 3816 23964
rect 3872 23962 3896 23964
rect 3952 23962 3976 23964
rect 3712 23910 3722 23962
rect 3966 23910 3976 23962
rect 3712 23908 3736 23910
rect 3792 23908 3816 23910
rect 3872 23908 3896 23910
rect 3952 23908 3976 23910
rect 3656 23899 4032 23908
rect 846 23831 902 23840
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 2916 23420 3292 23429
rect 2972 23418 2996 23420
rect 3052 23418 3076 23420
rect 3132 23418 3156 23420
rect 3212 23418 3236 23420
rect 2972 23366 2982 23418
rect 3226 23366 3236 23418
rect 2972 23364 2996 23366
rect 3052 23364 3076 23366
rect 3132 23364 3156 23366
rect 3212 23364 3236 23366
rect 2916 23355 3292 23364
rect 10916 23420 11292 23429
rect 10972 23418 10996 23420
rect 11052 23418 11076 23420
rect 11132 23418 11156 23420
rect 11212 23418 11236 23420
rect 10972 23366 10982 23418
rect 11226 23366 11236 23418
rect 10972 23364 10996 23366
rect 11052 23364 11076 23366
rect 11132 23364 11156 23366
rect 11212 23364 11236 23366
rect 10916 23355 11292 23364
rect 848 23112 900 23118
rect 846 23080 848 23089
rect 900 23080 902 23089
rect 846 23015 902 23024
rect 11152 22976 11204 22982
rect 11152 22918 11204 22924
rect 3656 22876 4032 22885
rect 3712 22874 3736 22876
rect 3792 22874 3816 22876
rect 3872 22874 3896 22876
rect 3952 22874 3976 22876
rect 3712 22822 3722 22874
rect 3966 22822 3976 22874
rect 3712 22820 3736 22822
rect 3792 22820 3816 22822
rect 3872 22820 3896 22822
rect 3952 22820 3976 22822
rect 3656 22811 4032 22820
rect 11164 22778 11192 22918
rect 11152 22772 11204 22778
rect 11152 22714 11204 22720
rect 848 22636 900 22642
rect 848 22578 900 22584
rect 860 22273 888 22578
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 846 22264 902 22273
rect 1596 22234 1624 22374
rect 2916 22332 3292 22341
rect 2972 22330 2996 22332
rect 3052 22330 3076 22332
rect 3132 22330 3156 22332
rect 3212 22330 3236 22332
rect 2972 22278 2982 22330
rect 3226 22278 3236 22330
rect 2972 22276 2996 22278
rect 3052 22276 3076 22278
rect 3132 22276 3156 22278
rect 3212 22276 3236 22278
rect 2916 22267 3292 22276
rect 10916 22332 11292 22341
rect 10972 22330 10996 22332
rect 11052 22330 11076 22332
rect 11132 22330 11156 22332
rect 11212 22330 11236 22332
rect 10972 22278 10982 22330
rect 11226 22278 11236 22330
rect 10972 22276 10996 22278
rect 11052 22276 11076 22278
rect 11132 22276 11156 22278
rect 11212 22276 11236 22278
rect 10916 22267 11292 22276
rect 846 22199 902 22208
rect 1584 22228 1636 22234
rect 1584 22170 1636 22176
rect 11348 22098 11376 24142
rect 11440 23798 11468 24550
rect 12084 24290 12112 25638
rect 12256 24336 12308 24342
rect 12084 24284 12256 24290
rect 12084 24278 12308 24284
rect 12084 24262 12296 24278
rect 11520 24200 11572 24206
rect 11520 24142 11572 24148
rect 11532 23866 11560 24142
rect 11656 23964 12032 23973
rect 11712 23962 11736 23964
rect 11792 23962 11816 23964
rect 11872 23962 11896 23964
rect 11952 23962 11976 23964
rect 11712 23910 11722 23962
rect 11966 23910 11976 23962
rect 11712 23908 11736 23910
rect 11792 23908 11816 23910
rect 11872 23908 11896 23910
rect 11952 23908 11976 23910
rect 11656 23899 12032 23908
rect 11520 23860 11572 23866
rect 11520 23802 11572 23808
rect 11428 23792 11480 23798
rect 11428 23734 11480 23740
rect 12084 23662 12112 24262
rect 12072 23656 12124 23662
rect 12072 23598 12124 23604
rect 12084 23254 12112 23598
rect 12072 23248 12124 23254
rect 12360 23202 12388 27406
rect 19656 27228 20032 27237
rect 19712 27226 19736 27228
rect 19792 27226 19816 27228
rect 19872 27226 19896 27228
rect 19952 27226 19976 27228
rect 19712 27174 19722 27226
rect 19966 27174 19976 27226
rect 19712 27172 19736 27174
rect 19792 27172 19816 27174
rect 19872 27172 19896 27174
rect 19952 27172 19976 27174
rect 19656 27163 20032 27172
rect 13268 27056 13320 27062
rect 13268 26998 13320 27004
rect 12440 26988 12492 26994
rect 12440 26930 12492 26936
rect 12072 23190 12124 23196
rect 11520 23044 11572 23050
rect 11520 22986 11572 22992
rect 11428 22432 11480 22438
rect 11428 22374 11480 22380
rect 11336 22092 11388 22098
rect 11336 22034 11388 22040
rect 11440 22030 11468 22374
rect 11428 22024 11480 22030
rect 11428 21966 11480 21972
rect 3656 21788 4032 21797
rect 3712 21786 3736 21788
rect 3792 21786 3816 21788
rect 3872 21786 3896 21788
rect 3952 21786 3976 21788
rect 3712 21734 3722 21786
rect 3966 21734 3976 21786
rect 3712 21732 3736 21734
rect 3792 21732 3816 21734
rect 3872 21732 3896 21734
rect 3952 21732 3976 21734
rect 3656 21723 4032 21732
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1412 21457 1440 21490
rect 1398 21448 1454 21457
rect 1398 21383 1454 21392
rect 2916 21244 3292 21253
rect 2972 21242 2996 21244
rect 3052 21242 3076 21244
rect 3132 21242 3156 21244
rect 3212 21242 3236 21244
rect 2972 21190 2982 21242
rect 3226 21190 3236 21242
rect 2972 21188 2996 21190
rect 3052 21188 3076 21190
rect 3132 21188 3156 21190
rect 3212 21188 3236 21190
rect 2916 21179 3292 21188
rect 10916 21244 11292 21253
rect 10972 21242 10996 21244
rect 11052 21242 11076 21244
rect 11132 21242 11156 21244
rect 11212 21242 11236 21244
rect 10972 21190 10982 21242
rect 11226 21190 11236 21242
rect 10972 21188 10996 21190
rect 11052 21188 11076 21190
rect 11132 21188 11156 21190
rect 11212 21188 11236 21190
rect 10916 21179 11292 21188
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1412 20641 1440 20878
rect 11336 20800 11388 20806
rect 11336 20742 11388 20748
rect 3656 20700 4032 20709
rect 3712 20698 3736 20700
rect 3792 20698 3816 20700
rect 3872 20698 3896 20700
rect 3952 20698 3976 20700
rect 3712 20646 3722 20698
rect 3966 20646 3976 20698
rect 3712 20644 3736 20646
rect 3792 20644 3816 20646
rect 3872 20644 3896 20646
rect 3952 20644 3976 20646
rect 1398 20632 1454 20641
rect 3656 20635 4032 20644
rect 1398 20567 1454 20576
rect 2916 20156 3292 20165
rect 2972 20154 2996 20156
rect 3052 20154 3076 20156
rect 3132 20154 3156 20156
rect 3212 20154 3236 20156
rect 2972 20102 2982 20154
rect 3226 20102 3236 20154
rect 2972 20100 2996 20102
rect 3052 20100 3076 20102
rect 3132 20100 3156 20102
rect 3212 20100 3236 20102
rect 2916 20091 3292 20100
rect 10916 20156 11292 20165
rect 10972 20154 10996 20156
rect 11052 20154 11076 20156
rect 11132 20154 11156 20156
rect 11212 20154 11236 20156
rect 10972 20102 10982 20154
rect 11226 20102 11236 20154
rect 10972 20100 10996 20102
rect 11052 20100 11076 20102
rect 11132 20100 11156 20102
rect 11212 20100 11236 20102
rect 10916 20091 11292 20100
rect 1400 19848 1452 19854
rect 1398 19816 1400 19825
rect 1452 19816 1454 19825
rect 1398 19751 1454 19760
rect 3656 19612 4032 19621
rect 3712 19610 3736 19612
rect 3792 19610 3816 19612
rect 3872 19610 3896 19612
rect 3952 19610 3976 19612
rect 3712 19558 3722 19610
rect 3966 19558 3976 19610
rect 3712 19556 3736 19558
rect 3792 19556 3816 19558
rect 3872 19556 3896 19558
rect 3952 19556 3976 19558
rect 3656 19547 4032 19556
rect 11348 19446 11376 20742
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 11440 19514 11468 19790
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 11336 19440 11388 19446
rect 11336 19382 11388 19388
rect 848 19372 900 19378
rect 848 19314 900 19320
rect 860 19009 888 19314
rect 11428 19304 11480 19310
rect 11428 19246 11480 19252
rect 2916 19068 3292 19077
rect 2972 19066 2996 19068
rect 3052 19066 3076 19068
rect 3132 19066 3156 19068
rect 3212 19066 3236 19068
rect 2972 19014 2982 19066
rect 3226 19014 3236 19066
rect 2972 19012 2996 19014
rect 3052 19012 3076 19014
rect 3132 19012 3156 19014
rect 3212 19012 3236 19014
rect 846 19000 902 19009
rect 2916 19003 3292 19012
rect 10916 19068 11292 19077
rect 10972 19066 10996 19068
rect 11052 19066 11076 19068
rect 11132 19066 11156 19068
rect 11212 19066 11236 19068
rect 10972 19014 10982 19066
rect 11226 19014 11236 19066
rect 10972 19012 10996 19014
rect 11052 19012 11076 19014
rect 11132 19012 11156 19014
rect 11212 19012 11236 19014
rect 10916 19003 11292 19012
rect 846 18935 902 18944
rect 3656 18524 4032 18533
rect 3712 18522 3736 18524
rect 3792 18522 3816 18524
rect 3872 18522 3896 18524
rect 3952 18522 3976 18524
rect 3712 18470 3722 18522
rect 3966 18470 3976 18522
rect 3712 18468 3736 18470
rect 3792 18468 3816 18470
rect 3872 18468 3896 18470
rect 3952 18468 3976 18470
rect 3656 18459 4032 18468
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1412 18057 1440 18226
rect 1398 18048 1454 18057
rect 1398 17983 1454 17992
rect 2916 17980 3292 17989
rect 2972 17978 2996 17980
rect 3052 17978 3076 17980
rect 3132 17978 3156 17980
rect 3212 17978 3236 17980
rect 2972 17926 2982 17978
rect 3226 17926 3236 17978
rect 2972 17924 2996 17926
rect 3052 17924 3076 17926
rect 3132 17924 3156 17926
rect 3212 17924 3236 17926
rect 2916 17915 3292 17924
rect 10916 17980 11292 17989
rect 10972 17978 10996 17980
rect 11052 17978 11076 17980
rect 11132 17978 11156 17980
rect 11212 17978 11236 17980
rect 10972 17926 10982 17978
rect 11226 17926 11236 17978
rect 10972 17924 10996 17926
rect 11052 17924 11076 17926
rect 11132 17924 11156 17926
rect 11212 17924 11236 17926
rect 10916 17915 11292 17924
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1412 17377 1440 17614
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 3656 17436 4032 17445
rect 3712 17434 3736 17436
rect 3792 17434 3816 17436
rect 3872 17434 3896 17436
rect 3952 17434 3976 17436
rect 3712 17382 3722 17434
rect 3966 17382 3976 17434
rect 3712 17380 3736 17382
rect 3792 17380 3816 17382
rect 3872 17380 3896 17382
rect 3952 17380 3976 17382
rect 1398 17368 1454 17377
rect 3656 17371 4032 17380
rect 1398 17303 1454 17312
rect 2916 16892 3292 16901
rect 2972 16890 2996 16892
rect 3052 16890 3076 16892
rect 3132 16890 3156 16892
rect 3212 16890 3236 16892
rect 2972 16838 2982 16890
rect 3226 16838 3236 16890
rect 2972 16836 2996 16838
rect 3052 16836 3076 16838
rect 3132 16836 3156 16838
rect 3212 16836 3236 16838
rect 2916 16827 3292 16836
rect 10916 16892 11292 16901
rect 10972 16890 10996 16892
rect 11052 16890 11076 16892
rect 11132 16890 11156 16892
rect 11212 16890 11236 16892
rect 10972 16838 10982 16890
rect 11226 16838 11236 16890
rect 10972 16836 10996 16838
rect 11052 16836 11076 16838
rect 11132 16836 11156 16838
rect 11212 16836 11236 16838
rect 10916 16827 11292 16836
rect 1400 16584 1452 16590
rect 1398 16552 1400 16561
rect 1452 16552 1454 16561
rect 1398 16487 1454 16496
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 3656 16348 4032 16357
rect 3712 16346 3736 16348
rect 3792 16346 3816 16348
rect 3872 16346 3896 16348
rect 3952 16346 3976 16348
rect 3712 16294 3722 16346
rect 3966 16294 3976 16346
rect 3712 16292 3736 16294
rect 3792 16292 3816 16294
rect 3872 16292 3896 16294
rect 3952 16292 3976 16294
rect 3656 16283 4032 16292
rect 10888 16250 10916 16390
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1412 15745 1440 16050
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 2916 15804 3292 15813
rect 2972 15802 2996 15804
rect 3052 15802 3076 15804
rect 3132 15802 3156 15804
rect 3212 15802 3236 15804
rect 2972 15750 2982 15802
rect 3226 15750 3236 15802
rect 2972 15748 2996 15750
rect 3052 15748 3076 15750
rect 3132 15748 3156 15750
rect 3212 15748 3236 15750
rect 1398 15736 1454 15745
rect 2916 15739 3292 15748
rect 1398 15671 1454 15680
rect 10704 15638 10732 15982
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 3656 15260 4032 15269
rect 3712 15258 3736 15260
rect 3792 15258 3816 15260
rect 3872 15258 3896 15260
rect 3952 15258 3976 15260
rect 3712 15206 3722 15258
rect 3966 15206 3976 15258
rect 3712 15204 3736 15206
rect 3792 15204 3816 15206
rect 3872 15204 3896 15206
rect 3952 15204 3976 15206
rect 3656 15195 4032 15204
rect 1400 15020 1452 15026
rect 1400 14962 1452 14968
rect 112 14952 164 14958
rect 1412 14929 1440 14962
rect 10704 14958 10732 15574
rect 10796 15162 10824 15846
rect 10916 15804 11292 15813
rect 10972 15802 10996 15804
rect 11052 15802 11076 15804
rect 11132 15802 11156 15804
rect 11212 15802 11236 15804
rect 10972 15750 10982 15802
rect 11226 15750 11236 15802
rect 10972 15748 10996 15750
rect 11052 15748 11076 15750
rect 11132 15748 11156 15750
rect 11212 15748 11236 15750
rect 10916 15739 11292 15748
rect 11348 15570 11376 17478
rect 11440 15706 11468 19246
rect 11532 17678 11560 22986
rect 11656 22876 12032 22885
rect 11712 22874 11736 22876
rect 11792 22874 11816 22876
rect 11872 22874 11896 22876
rect 11952 22874 11976 22876
rect 11712 22822 11722 22874
rect 11966 22822 11976 22874
rect 11712 22820 11736 22822
rect 11792 22820 11816 22822
rect 11872 22820 11896 22822
rect 11952 22820 11976 22822
rect 11656 22811 12032 22820
rect 12084 22574 12112 23190
rect 12176 23174 12388 23202
rect 12176 23118 12204 23174
rect 12164 23112 12216 23118
rect 12164 23054 12216 23060
rect 12072 22568 12124 22574
rect 12072 22510 12124 22516
rect 11656 21788 12032 21797
rect 11712 21786 11736 21788
rect 11792 21786 11816 21788
rect 11872 21786 11896 21788
rect 11952 21786 11976 21788
rect 11712 21734 11722 21786
rect 11966 21734 11976 21786
rect 11712 21732 11736 21734
rect 11792 21732 11816 21734
rect 11872 21732 11896 21734
rect 11952 21732 11976 21734
rect 11656 21723 12032 21732
rect 12176 21078 12204 23054
rect 12452 22642 12480 26930
rect 13280 26314 13308 26998
rect 21284 26858 21312 27406
rect 27656 27228 28032 27237
rect 27712 27226 27736 27228
rect 27792 27226 27816 27228
rect 27872 27226 27896 27228
rect 27952 27226 27976 27228
rect 27712 27174 27722 27226
rect 27966 27174 27976 27226
rect 27712 27172 27736 27174
rect 27792 27172 27816 27174
rect 27872 27172 27896 27174
rect 27952 27172 27976 27174
rect 27656 27163 28032 27172
rect 21364 26988 21416 26994
rect 21364 26930 21416 26936
rect 21272 26852 21324 26858
rect 21272 26794 21324 26800
rect 18916 26684 19292 26693
rect 18972 26682 18996 26684
rect 19052 26682 19076 26684
rect 19132 26682 19156 26684
rect 19212 26682 19236 26684
rect 18972 26630 18982 26682
rect 19226 26630 19236 26682
rect 18972 26628 18996 26630
rect 19052 26628 19076 26630
rect 19132 26628 19156 26630
rect 19212 26628 19236 26630
rect 18916 26619 19292 26628
rect 21376 26382 21404 26930
rect 28356 26920 28408 26926
rect 28356 26862 28408 26868
rect 28368 26761 28396 26862
rect 28354 26752 28410 26761
rect 26916 26684 27292 26693
rect 28354 26687 28410 26696
rect 26972 26682 26996 26684
rect 27052 26682 27076 26684
rect 27132 26682 27156 26684
rect 27212 26682 27236 26684
rect 26972 26630 26982 26682
rect 27226 26630 27236 26682
rect 26972 26628 26996 26630
rect 27052 26628 27076 26630
rect 27132 26628 27156 26630
rect 27212 26628 27236 26630
rect 26916 26619 27292 26628
rect 21364 26376 21416 26382
rect 21364 26318 21416 26324
rect 13268 26308 13320 26314
rect 13268 26250 13320 26256
rect 13544 26308 13596 26314
rect 13544 26250 13596 26256
rect 28356 26308 28408 26314
rect 28356 26250 28408 26256
rect 12992 26240 13044 26246
rect 12992 26182 13044 26188
rect 13004 25838 13032 26182
rect 13556 26042 13584 26250
rect 19656 26140 20032 26149
rect 19712 26138 19736 26140
rect 19792 26138 19816 26140
rect 19872 26138 19896 26140
rect 19952 26138 19976 26140
rect 19712 26086 19722 26138
rect 19966 26086 19976 26138
rect 19712 26084 19736 26086
rect 19792 26084 19816 26086
rect 19872 26084 19896 26086
rect 19952 26084 19976 26086
rect 19656 26075 20032 26084
rect 27656 26140 28032 26149
rect 27712 26138 27736 26140
rect 27792 26138 27816 26140
rect 27872 26138 27896 26140
rect 27952 26138 27976 26140
rect 27712 26086 27722 26138
rect 27966 26086 27976 26138
rect 27712 26084 27736 26086
rect 27792 26084 27816 26086
rect 27872 26084 27896 26086
rect 27952 26084 27976 26086
rect 27656 26075 28032 26084
rect 13544 26036 13596 26042
rect 13544 25978 13596 25984
rect 28368 25945 28396 26250
rect 28354 25936 28410 25945
rect 28354 25871 28410 25880
rect 12992 25832 13044 25838
rect 12992 25774 13044 25780
rect 18916 25596 19292 25605
rect 18972 25594 18996 25596
rect 19052 25594 19076 25596
rect 19132 25594 19156 25596
rect 19212 25594 19236 25596
rect 18972 25542 18982 25594
rect 19226 25542 19236 25594
rect 18972 25540 18996 25542
rect 19052 25540 19076 25542
rect 19132 25540 19156 25542
rect 19212 25540 19236 25542
rect 18916 25531 19292 25540
rect 26916 25596 27292 25605
rect 26972 25594 26996 25596
rect 27052 25594 27076 25596
rect 27132 25594 27156 25596
rect 27212 25594 27236 25596
rect 26972 25542 26982 25594
rect 27226 25542 27236 25594
rect 26972 25540 26996 25542
rect 27052 25540 27076 25542
rect 27132 25540 27156 25542
rect 27212 25540 27236 25542
rect 26916 25531 27292 25540
rect 28356 25220 28408 25226
rect 28356 25162 28408 25168
rect 12808 25152 12860 25158
rect 28368 25129 28396 25162
rect 12808 25094 12860 25100
rect 28354 25120 28410 25129
rect 12820 24886 12848 25094
rect 19656 25052 20032 25061
rect 19712 25050 19736 25052
rect 19792 25050 19816 25052
rect 19872 25050 19896 25052
rect 19952 25050 19976 25052
rect 19712 24998 19722 25050
rect 19966 24998 19976 25050
rect 19712 24996 19736 24998
rect 19792 24996 19816 24998
rect 19872 24996 19896 24998
rect 19952 24996 19976 24998
rect 19656 24987 20032 24996
rect 27656 25052 28032 25061
rect 28354 25055 28410 25064
rect 27712 25050 27736 25052
rect 27792 25050 27816 25052
rect 27872 25050 27896 25052
rect 27952 25050 27976 25052
rect 27712 24998 27722 25050
rect 27966 24998 27976 25050
rect 27712 24996 27736 24998
rect 27792 24996 27816 24998
rect 27872 24996 27896 24998
rect 27952 24996 27976 24998
rect 27656 24987 28032 24996
rect 12808 24880 12860 24886
rect 12808 24822 12860 24828
rect 12820 24154 12848 24822
rect 13360 24812 13412 24818
rect 13360 24754 13412 24760
rect 12992 24744 13044 24750
rect 12992 24686 13044 24692
rect 13004 24410 13032 24686
rect 12992 24404 13044 24410
rect 12992 24346 13044 24352
rect 13372 24206 13400 24754
rect 28356 24744 28408 24750
rect 28356 24686 28408 24692
rect 18916 24508 19292 24517
rect 18972 24506 18996 24508
rect 19052 24506 19076 24508
rect 19132 24506 19156 24508
rect 19212 24506 19236 24508
rect 18972 24454 18982 24506
rect 19226 24454 19236 24506
rect 18972 24452 18996 24454
rect 19052 24452 19076 24454
rect 19132 24452 19156 24454
rect 19212 24452 19236 24454
rect 18916 24443 19292 24452
rect 26916 24508 27292 24517
rect 26972 24506 26996 24508
rect 27052 24506 27076 24508
rect 27132 24506 27156 24508
rect 27212 24506 27236 24508
rect 26972 24454 26982 24506
rect 27226 24454 27236 24506
rect 26972 24452 26996 24454
rect 27052 24452 27076 24454
rect 27132 24452 27156 24454
rect 27212 24452 27236 24454
rect 26916 24443 27292 24452
rect 28368 24313 28396 24686
rect 28354 24304 28410 24313
rect 28354 24239 28410 24248
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12728 24126 12848 24154
rect 13360 24200 13412 24206
rect 13360 24142 13412 24148
rect 28080 24132 28132 24138
rect 12636 23866 12664 24074
rect 12728 24070 12756 24126
rect 28080 24074 28132 24080
rect 12716 24064 12768 24070
rect 12716 24006 12768 24012
rect 12624 23860 12676 23866
rect 12624 23802 12676 23808
rect 12624 22704 12676 22710
rect 12624 22646 12676 22652
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12164 21072 12216 21078
rect 12164 21014 12216 21020
rect 11656 20700 12032 20709
rect 11712 20698 11736 20700
rect 11792 20698 11816 20700
rect 11872 20698 11896 20700
rect 11952 20698 11976 20700
rect 11712 20646 11722 20698
rect 11966 20646 11976 20698
rect 11712 20644 11736 20646
rect 11792 20644 11816 20646
rect 11872 20644 11896 20646
rect 11952 20644 11976 20646
rect 11656 20635 12032 20644
rect 11656 19612 12032 19621
rect 11712 19610 11736 19612
rect 11792 19610 11816 19612
rect 11872 19610 11896 19612
rect 11952 19610 11976 19612
rect 11712 19558 11722 19610
rect 11966 19558 11976 19610
rect 11712 19556 11736 19558
rect 11792 19556 11816 19558
rect 11872 19556 11896 19558
rect 11952 19556 11976 19558
rect 11656 19547 12032 19556
rect 12176 19310 12204 21014
rect 12452 20602 12480 22578
rect 12636 21962 12664 22646
rect 12728 22506 12756 24006
rect 19656 23964 20032 23973
rect 19712 23962 19736 23964
rect 19792 23962 19816 23964
rect 19872 23962 19896 23964
rect 19952 23962 19976 23964
rect 19712 23910 19722 23962
rect 19966 23910 19976 23962
rect 19712 23908 19736 23910
rect 19792 23908 19816 23910
rect 19872 23908 19896 23910
rect 19952 23908 19976 23910
rect 19656 23899 20032 23908
rect 27656 23964 28032 23973
rect 27712 23962 27736 23964
rect 27792 23962 27816 23964
rect 27872 23962 27896 23964
rect 27952 23962 27976 23964
rect 27712 23910 27722 23962
rect 27966 23910 27976 23962
rect 27712 23908 27736 23910
rect 27792 23908 27816 23910
rect 27872 23908 27896 23910
rect 27952 23908 27976 23910
rect 27656 23899 28032 23908
rect 28092 23730 28120 24074
rect 14556 23724 14608 23730
rect 14556 23666 14608 23672
rect 28080 23724 28132 23730
rect 28080 23666 28132 23672
rect 14568 23186 14596 23666
rect 28356 23656 28408 23662
rect 28356 23598 28408 23604
rect 28368 23497 28396 23598
rect 28354 23488 28410 23497
rect 18916 23420 19292 23429
rect 18972 23418 18996 23420
rect 19052 23418 19076 23420
rect 19132 23418 19156 23420
rect 19212 23418 19236 23420
rect 18972 23366 18982 23418
rect 19226 23366 19236 23418
rect 18972 23364 18996 23366
rect 19052 23364 19076 23366
rect 19132 23364 19156 23366
rect 19212 23364 19236 23366
rect 18916 23355 19292 23364
rect 26916 23420 27292 23429
rect 28354 23423 28410 23432
rect 26972 23418 26996 23420
rect 27052 23418 27076 23420
rect 27132 23418 27156 23420
rect 27212 23418 27236 23420
rect 26972 23366 26982 23418
rect 27226 23366 27236 23418
rect 26972 23364 26996 23366
rect 27052 23364 27076 23366
rect 27132 23364 27156 23366
rect 27212 23364 27236 23366
rect 26916 23355 27292 23364
rect 14556 23180 14608 23186
rect 14556 23122 14608 23128
rect 14648 23180 14700 23186
rect 14648 23122 14700 23128
rect 13084 22976 13136 22982
rect 13084 22918 13136 22924
rect 13452 22976 13504 22982
rect 13452 22918 13504 22924
rect 13096 22574 13124 22918
rect 13464 22642 13492 22918
rect 13820 22704 13872 22710
rect 13740 22652 13820 22658
rect 13740 22646 13872 22652
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 13740 22630 13860 22646
rect 13084 22568 13136 22574
rect 13084 22510 13136 22516
rect 12716 22500 12768 22506
rect 12716 22442 12768 22448
rect 12728 22030 12756 22442
rect 13096 22098 13124 22510
rect 13084 22092 13136 22098
rect 13084 22034 13136 22040
rect 12716 22024 12768 22030
rect 12716 21966 12768 21972
rect 12624 21956 12676 21962
rect 12624 21898 12676 21904
rect 13096 21554 13124 22034
rect 13740 22030 13768 22630
rect 14660 22166 14688 23122
rect 14924 23112 14976 23118
rect 14924 23054 14976 23060
rect 14936 22778 14964 23054
rect 28356 23044 28408 23050
rect 28356 22986 28408 22992
rect 19656 22876 20032 22885
rect 19712 22874 19736 22876
rect 19792 22874 19816 22876
rect 19872 22874 19896 22876
rect 19952 22874 19976 22876
rect 19712 22822 19722 22874
rect 19966 22822 19976 22874
rect 19712 22820 19736 22822
rect 19792 22820 19816 22822
rect 19872 22820 19896 22822
rect 19952 22820 19976 22822
rect 19656 22811 20032 22820
rect 27656 22876 28032 22885
rect 27712 22874 27736 22876
rect 27792 22874 27816 22876
rect 27872 22874 27896 22876
rect 27952 22874 27976 22876
rect 27712 22822 27722 22874
rect 27966 22822 27976 22874
rect 27712 22820 27736 22822
rect 27792 22820 27816 22822
rect 27872 22820 27896 22822
rect 27952 22820 27976 22822
rect 27656 22811 28032 22820
rect 14924 22772 14976 22778
rect 14924 22714 14976 22720
rect 28368 22681 28396 22986
rect 28354 22672 28410 22681
rect 28354 22607 28410 22616
rect 18916 22332 19292 22341
rect 18972 22330 18996 22332
rect 19052 22330 19076 22332
rect 19132 22330 19156 22332
rect 19212 22330 19236 22332
rect 18972 22278 18982 22330
rect 19226 22278 19236 22330
rect 18972 22276 18996 22278
rect 19052 22276 19076 22278
rect 19132 22276 19156 22278
rect 19212 22276 19236 22278
rect 18916 22267 19292 22276
rect 26916 22332 27292 22341
rect 26972 22330 26996 22332
rect 27052 22330 27076 22332
rect 27132 22330 27156 22332
rect 27212 22330 27236 22332
rect 26972 22278 26982 22330
rect 27226 22278 27236 22330
rect 26972 22276 26996 22278
rect 27052 22276 27076 22278
rect 27132 22276 27156 22278
rect 27212 22276 27236 22278
rect 26916 22267 27292 22276
rect 14648 22160 14700 22166
rect 14648 22102 14700 22108
rect 13728 22024 13780 22030
rect 13728 21966 13780 21972
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13464 21554 13492 21830
rect 13740 21690 13768 21966
rect 14832 21956 14884 21962
rect 14832 21898 14884 21904
rect 17868 21956 17920 21962
rect 17868 21898 17920 21904
rect 28356 21956 28408 21962
rect 28356 21898 28408 21904
rect 14844 21690 14872 21898
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 17880 21554 17908 21898
rect 28368 21865 28396 21898
rect 28354 21856 28410 21865
rect 19656 21788 20032 21797
rect 19712 21786 19736 21788
rect 19792 21786 19816 21788
rect 19872 21786 19896 21788
rect 19952 21786 19976 21788
rect 19712 21734 19722 21786
rect 19966 21734 19976 21786
rect 19712 21732 19736 21734
rect 19792 21732 19816 21734
rect 19872 21732 19896 21734
rect 19952 21732 19976 21734
rect 19656 21723 20032 21732
rect 27656 21788 28032 21797
rect 28354 21791 28410 21800
rect 27712 21786 27736 21788
rect 27792 21786 27816 21788
rect 27872 21786 27896 21788
rect 27952 21786 27976 21788
rect 27712 21734 27722 21786
rect 27966 21734 27976 21786
rect 27712 21732 27736 21734
rect 27792 21732 27816 21734
rect 27872 21732 27896 21734
rect 27952 21732 27976 21734
rect 27656 21723 28032 21732
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 28356 21480 28408 21486
rect 28356 21422 28408 21428
rect 14556 21344 14608 21350
rect 14556 21286 14608 21292
rect 14568 21010 14596 21286
rect 18916 21244 19292 21253
rect 18972 21242 18996 21244
rect 19052 21242 19076 21244
rect 19132 21242 19156 21244
rect 19212 21242 19236 21244
rect 18972 21190 18982 21242
rect 19226 21190 19236 21242
rect 18972 21188 18996 21190
rect 19052 21188 19076 21190
rect 19132 21188 19156 21190
rect 19212 21188 19236 21190
rect 18916 21179 19292 21188
rect 26916 21244 27292 21253
rect 26972 21242 26996 21244
rect 27052 21242 27076 21244
rect 27132 21242 27156 21244
rect 27212 21242 27236 21244
rect 26972 21190 26982 21242
rect 27226 21190 27236 21242
rect 26972 21188 26996 21190
rect 27052 21188 27076 21190
rect 27132 21188 27156 21190
rect 27212 21188 27236 21190
rect 26916 21179 27292 21188
rect 28368 21049 28396 21422
rect 28354 21040 28410 21049
rect 14556 21004 14608 21010
rect 28354 20975 28410 20984
rect 14556 20946 14608 20952
rect 14648 20868 14700 20874
rect 14648 20810 14700 20816
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 12360 19922 12388 20334
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 12268 19514 12296 19790
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 12360 19378 12388 19858
rect 12452 19786 12480 20538
rect 13924 20398 13952 20742
rect 14660 20466 14688 20810
rect 19656 20700 20032 20709
rect 19712 20698 19736 20700
rect 19792 20698 19816 20700
rect 19872 20698 19896 20700
rect 19952 20698 19976 20700
rect 19712 20646 19722 20698
rect 19966 20646 19976 20698
rect 19712 20644 19736 20646
rect 19792 20644 19816 20646
rect 19872 20644 19896 20646
rect 19952 20644 19976 20646
rect 19656 20635 20032 20644
rect 27656 20700 28032 20709
rect 27712 20698 27736 20700
rect 27792 20698 27816 20700
rect 27872 20698 27896 20700
rect 27952 20698 27976 20700
rect 27712 20646 27722 20698
rect 27966 20646 27976 20698
rect 27712 20644 27736 20646
rect 27792 20644 27816 20646
rect 27872 20644 27896 20646
rect 27952 20644 27976 20646
rect 27656 20635 28032 20644
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 28356 20392 28408 20398
rect 28356 20334 28408 20340
rect 28368 20233 28396 20334
rect 28354 20224 28410 20233
rect 18916 20156 19292 20165
rect 18972 20154 18996 20156
rect 19052 20154 19076 20156
rect 19132 20154 19156 20156
rect 19212 20154 19236 20156
rect 18972 20102 18982 20154
rect 19226 20102 19236 20154
rect 18972 20100 18996 20102
rect 19052 20100 19076 20102
rect 19132 20100 19156 20102
rect 19212 20100 19236 20102
rect 18916 20091 19292 20100
rect 26916 20156 27292 20165
rect 28354 20159 28410 20168
rect 26972 20154 26996 20156
rect 27052 20154 27076 20156
rect 27132 20154 27156 20156
rect 27212 20154 27236 20156
rect 26972 20102 26982 20154
rect 27226 20102 27236 20154
rect 26972 20100 26996 20102
rect 27052 20100 27076 20102
rect 27132 20100 27156 20102
rect 27212 20100 27236 20102
rect 26916 20091 27292 20100
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 12440 19780 12492 19786
rect 12440 19722 12492 19728
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12360 18698 12388 19314
rect 12452 18850 12480 19722
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13004 19378 13032 19654
rect 13556 19514 13584 19654
rect 13544 19508 13596 19514
rect 13544 19450 13596 19456
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 12452 18822 12664 18850
rect 12348 18692 12400 18698
rect 12348 18634 12400 18640
rect 11656 18524 12032 18533
rect 11712 18522 11736 18524
rect 11792 18522 11816 18524
rect 11872 18522 11896 18524
rect 11952 18522 11976 18524
rect 11712 18470 11722 18522
rect 11966 18470 11976 18522
rect 11712 18468 11736 18470
rect 11792 18468 11816 18470
rect 11872 18468 11896 18470
rect 11952 18468 11976 18470
rect 11656 18459 12032 18468
rect 12360 18222 12388 18634
rect 12348 18216 12400 18222
rect 12348 18158 12400 18164
rect 12360 17882 12388 18158
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 11656 17436 12032 17445
rect 11712 17434 11736 17436
rect 11792 17434 11816 17436
rect 11872 17434 11896 17436
rect 11952 17434 11976 17436
rect 11712 17382 11722 17434
rect 11966 17382 11976 17434
rect 11712 17380 11736 17382
rect 11792 17380 11816 17382
rect 11872 17380 11896 17382
rect 11952 17380 11976 17382
rect 11656 17371 12032 17380
rect 11520 17128 11572 17134
rect 11520 17070 11572 17076
rect 11532 16590 11560 17070
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 11532 16114 11560 16526
rect 11656 16348 12032 16357
rect 11712 16346 11736 16348
rect 11792 16346 11816 16348
rect 11872 16346 11896 16348
rect 11952 16346 11976 16348
rect 11712 16294 11722 16346
rect 11966 16294 11976 16346
rect 11712 16292 11736 16294
rect 11792 16292 11816 16294
rect 11872 16292 11896 16294
rect 11952 16292 11976 16294
rect 11656 16283 12032 16292
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 12084 15706 12112 16526
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11440 15502 11468 15642
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11610 15464 11666 15473
rect 11610 15399 11612 15408
rect 11664 15399 11666 15408
rect 11612 15370 11664 15376
rect 11656 15260 12032 15269
rect 11712 15258 11736 15260
rect 11792 15258 11816 15260
rect 11872 15258 11896 15260
rect 11952 15258 11976 15260
rect 11712 15206 11722 15258
rect 11966 15206 11976 15258
rect 11712 15204 11736 15206
rect 11792 15204 11816 15206
rect 11872 15204 11896 15206
rect 11952 15204 11976 15206
rect 11656 15195 12032 15204
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 10692 14952 10744 14958
rect 112 14894 164 14900
rect 1398 14920 1454 14929
rect 124 1193 152 14894
rect 10692 14894 10744 14900
rect 1398 14855 1454 14864
rect 11520 14884 11572 14890
rect 11520 14826 11572 14832
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 2916 14716 3292 14725
rect 2972 14714 2996 14716
rect 3052 14714 3076 14716
rect 3132 14714 3156 14716
rect 3212 14714 3236 14716
rect 2972 14662 2982 14714
rect 3226 14662 3236 14714
rect 2972 14660 2996 14662
rect 3052 14660 3076 14662
rect 3132 14660 3156 14662
rect 3212 14660 3236 14662
rect 2916 14651 3292 14660
rect 10796 14482 10824 14758
rect 10916 14716 11292 14725
rect 10972 14714 10996 14716
rect 11052 14714 11076 14716
rect 11132 14714 11156 14716
rect 11212 14714 11236 14716
rect 10972 14662 10982 14714
rect 11226 14662 11236 14714
rect 10972 14660 10996 14662
rect 11052 14660 11076 14662
rect 11132 14660 11156 14662
rect 11212 14660 11236 14662
rect 10916 14651 11292 14660
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 1412 14113 1440 14350
rect 3656 14172 4032 14181
rect 3712 14170 3736 14172
rect 3792 14170 3816 14172
rect 3872 14170 3896 14172
rect 3952 14170 3976 14172
rect 3712 14118 3722 14170
rect 3966 14118 3976 14170
rect 3712 14116 3736 14118
rect 3792 14116 3816 14118
rect 3872 14116 3896 14118
rect 3952 14116 3976 14118
rect 1398 14104 1454 14113
rect 3656 14107 4032 14116
rect 1398 14039 1454 14048
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 2916 13628 3292 13637
rect 2972 13626 2996 13628
rect 3052 13626 3076 13628
rect 3132 13626 3156 13628
rect 3212 13626 3236 13628
rect 2972 13574 2982 13626
rect 3226 13574 3236 13626
rect 2972 13572 2996 13574
rect 3052 13572 3076 13574
rect 3132 13572 3156 13574
rect 3212 13572 3236 13574
rect 2916 13563 3292 13572
rect 1400 13320 1452 13326
rect 1398 13288 1400 13297
rect 1452 13288 1454 13297
rect 1398 13223 1454 13232
rect 3656 13084 4032 13093
rect 3712 13082 3736 13084
rect 3792 13082 3816 13084
rect 3872 13082 3896 13084
rect 3952 13082 3976 13084
rect 3712 13030 3722 13082
rect 3966 13030 3976 13082
rect 3712 13028 3736 13030
rect 3792 13028 3816 13030
rect 3872 13028 3896 13030
rect 3952 13028 3976 13030
rect 3656 13019 4032 13028
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12481 1440 12786
rect 2916 12540 3292 12549
rect 2972 12538 2996 12540
rect 3052 12538 3076 12540
rect 3132 12538 3156 12540
rect 3212 12538 3236 12540
rect 2972 12486 2982 12538
rect 3226 12486 3236 12538
rect 2972 12484 2996 12486
rect 3052 12484 3076 12486
rect 3132 12484 3156 12486
rect 3212 12484 3236 12486
rect 1398 12472 1454 12481
rect 2916 12475 3292 12484
rect 1398 12407 1454 12416
rect 3656 11996 4032 12005
rect 3712 11994 3736 11996
rect 3792 11994 3816 11996
rect 3872 11994 3896 11996
rect 3952 11994 3976 11996
rect 3712 11942 3722 11994
rect 3966 11942 3976 11994
rect 3712 11940 3736 11942
rect 3792 11940 3816 11942
rect 3872 11940 3896 11942
rect 3952 11940 3976 11942
rect 3656 11931 4032 11940
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1412 11665 1440 11698
rect 1398 11656 1454 11665
rect 1398 11591 1454 11600
rect 2916 11452 3292 11461
rect 2972 11450 2996 11452
rect 3052 11450 3076 11452
rect 3132 11450 3156 11452
rect 3212 11450 3236 11452
rect 2972 11398 2982 11450
rect 3226 11398 3236 11450
rect 2972 11396 2996 11398
rect 3052 11396 3076 11398
rect 3132 11396 3156 11398
rect 3212 11396 3236 11398
rect 2916 11387 3292 11396
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10849 1440 11086
rect 3656 10908 4032 10917
rect 3712 10906 3736 10908
rect 3792 10906 3816 10908
rect 3872 10906 3896 10908
rect 3952 10906 3976 10908
rect 3712 10854 3722 10906
rect 3966 10854 3976 10906
rect 3712 10852 3736 10854
rect 3792 10852 3816 10854
rect 3872 10852 3896 10854
rect 3952 10852 3976 10854
rect 1398 10840 1454 10849
rect 3656 10843 4032 10852
rect 1398 10775 1454 10784
rect 10336 10742 10364 13806
rect 10704 13326 10732 14350
rect 11532 14074 11560 14826
rect 11808 14414 11836 14962
rect 12176 14822 12204 17614
rect 12360 17134 12388 17818
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12452 17202 12480 17478
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12452 16182 12480 16390
rect 12440 16176 12492 16182
rect 12440 16118 12492 16124
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 12164 14272 12216 14278
rect 12164 14214 12216 14220
rect 11656 14172 12032 14181
rect 11712 14170 11736 14172
rect 11792 14170 11816 14172
rect 11872 14170 11896 14172
rect 11952 14170 11976 14172
rect 11712 14118 11722 14170
rect 11966 14118 11976 14170
rect 11712 14116 11736 14118
rect 11792 14116 11816 14118
rect 11872 14116 11896 14118
rect 11952 14116 11976 14118
rect 11656 14107 12032 14116
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 10916 13628 11292 13637
rect 10972 13626 10996 13628
rect 11052 13626 11076 13628
rect 11132 13626 11156 13628
rect 11212 13626 11236 13628
rect 10972 13574 10982 13626
rect 11226 13574 11236 13626
rect 10972 13572 10996 13574
rect 11052 13572 11076 13574
rect 11132 13572 11156 13574
rect 11212 13572 11236 13574
rect 10916 13563 11292 13572
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10704 12646 10732 13262
rect 10796 12782 10824 13466
rect 11532 13394 11560 13670
rect 12176 13394 12204 14214
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10888 12986 10916 13126
rect 11656 13084 12032 13093
rect 11712 13082 11736 13084
rect 11792 13082 11816 13084
rect 11872 13082 11896 13084
rect 11952 13082 11976 13084
rect 11712 13030 11722 13082
rect 11966 13030 11976 13082
rect 11712 13028 11736 13030
rect 11792 13028 11816 13030
rect 11872 13028 11896 13030
rect 11952 13028 11976 13030
rect 11656 13019 12032 13028
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10612 10810 10640 12582
rect 10704 12238 10732 12582
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10704 11694 10732 12174
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10704 11150 10732 11630
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 2916 10364 3292 10373
rect 2972 10362 2996 10364
rect 3052 10362 3076 10364
rect 3132 10362 3156 10364
rect 3212 10362 3236 10364
rect 2972 10310 2982 10362
rect 3226 10310 3236 10362
rect 2972 10308 2996 10310
rect 3052 10308 3076 10310
rect 3132 10308 3156 10310
rect 3212 10308 3236 10310
rect 2916 10299 3292 10308
rect 10704 10062 10732 11086
rect 10796 10606 10824 12718
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 10916 12540 11292 12549
rect 10972 12538 10996 12540
rect 11052 12538 11076 12540
rect 11132 12538 11156 12540
rect 11212 12538 11236 12540
rect 10972 12486 10982 12538
rect 11226 12486 11236 12538
rect 10972 12484 10996 12486
rect 11052 12484 11076 12486
rect 11132 12484 11156 12486
rect 11212 12484 11236 12486
rect 10916 12475 11292 12484
rect 11348 12306 11376 12582
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11992 12238 12020 12786
rect 12268 12434 12296 15438
rect 12452 14278 12480 16118
rect 12636 15366 12664 18822
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12728 18290 12756 18566
rect 13740 18358 13768 19382
rect 13832 18834 13860 19858
rect 28356 19780 28408 19786
rect 28356 19722 28408 19728
rect 19656 19612 20032 19621
rect 19712 19610 19736 19612
rect 19792 19610 19816 19612
rect 19872 19610 19896 19612
rect 19952 19610 19976 19612
rect 19712 19558 19722 19610
rect 19966 19558 19976 19610
rect 19712 19556 19736 19558
rect 19792 19556 19816 19558
rect 19872 19556 19896 19558
rect 19952 19556 19976 19558
rect 19656 19547 20032 19556
rect 27656 19612 28032 19621
rect 27712 19610 27736 19612
rect 27792 19610 27816 19612
rect 27872 19610 27896 19612
rect 27952 19610 27976 19612
rect 27712 19558 27722 19610
rect 27966 19558 27976 19610
rect 27712 19556 27736 19558
rect 27792 19556 27816 19558
rect 27872 19556 27896 19558
rect 27952 19556 27976 19558
rect 27656 19547 28032 19556
rect 28368 19417 28396 19722
rect 28354 19408 28410 19417
rect 23480 19372 23532 19378
rect 28354 19343 28410 19352
rect 23480 19314 23532 19320
rect 14556 19304 14608 19310
rect 14556 19246 14608 19252
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 14568 18766 14596 19246
rect 18916 19068 19292 19077
rect 18972 19066 18996 19068
rect 19052 19066 19076 19068
rect 19132 19066 19156 19068
rect 19212 19066 19236 19068
rect 18972 19014 18982 19066
rect 19226 19014 19236 19066
rect 18972 19012 18996 19014
rect 19052 19012 19076 19014
rect 19132 19012 19156 19014
rect 19212 19012 19236 19014
rect 18916 19003 19292 19012
rect 14648 18828 14700 18834
rect 14648 18770 14700 18776
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 13728 18352 13780 18358
rect 13728 18294 13780 18300
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 13740 17270 13768 18294
rect 14476 18290 14504 18566
rect 14556 18420 14608 18426
rect 14556 18362 14608 18368
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14568 17746 14596 18362
rect 14660 17746 14688 18770
rect 23492 18766 23520 19314
rect 26916 19068 27292 19077
rect 26972 19066 26996 19068
rect 27052 19066 27076 19068
rect 27132 19066 27156 19068
rect 27212 19066 27236 19068
rect 26972 19014 26982 19066
rect 27226 19014 27236 19066
rect 26972 19012 26996 19014
rect 27052 19012 27076 19014
rect 27132 19012 27156 19014
rect 27212 19012 27236 19014
rect 26916 19003 27292 19012
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 28356 18692 28408 18698
rect 28356 18634 28408 18640
rect 28368 18601 28396 18634
rect 28354 18592 28410 18601
rect 19656 18524 20032 18533
rect 19712 18522 19736 18524
rect 19792 18522 19816 18524
rect 19872 18522 19896 18524
rect 19952 18522 19976 18524
rect 19712 18470 19722 18522
rect 19966 18470 19976 18522
rect 19712 18468 19736 18470
rect 19792 18468 19816 18470
rect 19872 18468 19896 18470
rect 19952 18468 19976 18470
rect 19656 18459 20032 18468
rect 27656 18524 28032 18533
rect 28354 18527 28410 18536
rect 27712 18522 27736 18524
rect 27792 18522 27816 18524
rect 27872 18522 27896 18524
rect 27952 18522 27976 18524
rect 27712 18470 27722 18522
rect 27966 18470 27976 18522
rect 27712 18468 27736 18470
rect 27792 18468 27816 18470
rect 27872 18468 27896 18470
rect 27952 18468 27976 18470
rect 27656 18459 28032 18468
rect 28356 18216 28408 18222
rect 28356 18158 28408 18164
rect 18916 17980 19292 17989
rect 18972 17978 18996 17980
rect 19052 17978 19076 17980
rect 19132 17978 19156 17980
rect 19212 17978 19236 17980
rect 18972 17926 18982 17978
rect 19226 17926 19236 17978
rect 18972 17924 18996 17926
rect 19052 17924 19076 17926
rect 19132 17924 19156 17926
rect 19212 17924 19236 17926
rect 18916 17915 19292 17924
rect 26916 17980 27292 17989
rect 26972 17978 26996 17980
rect 27052 17978 27076 17980
rect 27132 17978 27156 17980
rect 27212 17978 27236 17980
rect 26972 17926 26982 17978
rect 27226 17926 27236 17978
rect 26972 17924 26996 17926
rect 27052 17924 27076 17926
rect 27132 17924 27156 17926
rect 27212 17924 27236 17926
rect 26916 17915 27292 17924
rect 28368 17785 28396 18158
rect 28354 17776 28410 17785
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 14648 17740 14700 17746
rect 28354 17711 28410 17720
rect 14648 17682 14700 17688
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 14476 17202 14504 17478
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 13004 16574 13032 17070
rect 12912 16546 13032 16574
rect 12912 16454 12940 16546
rect 12900 16448 12952 16454
rect 12900 16390 12952 16396
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13464 15434 13492 16390
rect 14660 15570 14688 17682
rect 19656 17436 20032 17445
rect 19712 17434 19736 17436
rect 19792 17434 19816 17436
rect 19872 17434 19896 17436
rect 19952 17434 19976 17436
rect 19712 17382 19722 17434
rect 19966 17382 19976 17434
rect 19712 17380 19736 17382
rect 19792 17380 19816 17382
rect 19872 17380 19896 17382
rect 19952 17380 19976 17382
rect 19656 17371 20032 17380
rect 27656 17436 28032 17445
rect 27712 17434 27736 17436
rect 27792 17434 27816 17436
rect 27872 17434 27896 17436
rect 27952 17434 27976 17436
rect 27712 17382 27722 17434
rect 27966 17382 27976 17434
rect 27712 17380 27736 17382
rect 27792 17380 27816 17382
rect 27872 17380 27896 17382
rect 27952 17380 27976 17382
rect 27656 17371 28032 17380
rect 28356 17128 28408 17134
rect 28356 17070 28408 17076
rect 28368 16969 28396 17070
rect 28354 16960 28410 16969
rect 18916 16892 19292 16901
rect 18972 16890 18996 16892
rect 19052 16890 19076 16892
rect 19132 16890 19156 16892
rect 19212 16890 19236 16892
rect 18972 16838 18982 16890
rect 19226 16838 19236 16890
rect 18972 16836 18996 16838
rect 19052 16836 19076 16838
rect 19132 16836 19156 16838
rect 19212 16836 19236 16838
rect 18916 16827 19292 16836
rect 26916 16892 27292 16901
rect 28354 16895 28410 16904
rect 26972 16890 26996 16892
rect 27052 16890 27076 16892
rect 27132 16890 27156 16892
rect 27212 16890 27236 16892
rect 26972 16838 26982 16890
rect 27226 16838 27236 16890
rect 26972 16836 26996 16838
rect 27052 16836 27076 16838
rect 27132 16836 27156 16838
rect 27212 16836 27236 16838
rect 26916 16827 27292 16836
rect 21364 16584 21416 16590
rect 21364 16526 21416 16532
rect 19656 16348 20032 16357
rect 19712 16346 19736 16348
rect 19792 16346 19816 16348
rect 19872 16346 19896 16348
rect 19952 16346 19976 16348
rect 19712 16294 19722 16346
rect 19966 16294 19976 16346
rect 19712 16292 19736 16294
rect 19792 16292 19816 16294
rect 19872 16292 19896 16294
rect 19952 16292 19976 16294
rect 19656 16283 20032 16292
rect 18916 15804 19292 15813
rect 18972 15802 18996 15804
rect 19052 15802 19076 15804
rect 19132 15802 19156 15804
rect 19212 15802 19236 15804
rect 18972 15750 18982 15802
rect 19226 15750 19236 15802
rect 18972 15748 18996 15750
rect 19052 15748 19076 15750
rect 19132 15748 19156 15750
rect 19212 15748 19236 15750
rect 18916 15739 19292 15748
rect 14648 15564 14700 15570
rect 14648 15506 14700 15512
rect 21376 15434 21404 16526
rect 28356 16516 28408 16522
rect 28356 16458 28408 16464
rect 27656 16348 28032 16357
rect 27712 16346 27736 16348
rect 27792 16346 27816 16348
rect 27872 16346 27896 16348
rect 27952 16346 27976 16348
rect 27712 16294 27722 16346
rect 27966 16294 27976 16346
rect 27712 16292 27736 16294
rect 27792 16292 27816 16294
rect 27872 16292 27896 16294
rect 27952 16292 27976 16294
rect 27656 16283 28032 16292
rect 28368 16153 28396 16458
rect 28354 16144 28410 16153
rect 28354 16079 28410 16088
rect 28080 15904 28132 15910
rect 28080 15846 28132 15852
rect 26916 15804 27292 15813
rect 26972 15802 26996 15804
rect 27052 15802 27076 15804
rect 27132 15802 27156 15804
rect 27212 15802 27236 15804
rect 26972 15750 26982 15802
rect 27226 15750 27236 15802
rect 26972 15748 26996 15750
rect 27052 15748 27076 15750
rect 27132 15748 27156 15750
rect 27212 15748 27236 15750
rect 26916 15739 27292 15748
rect 28092 15502 28120 15846
rect 28080 15496 28132 15502
rect 28080 15438 28132 15444
rect 13452 15428 13504 15434
rect 13452 15370 13504 15376
rect 21364 15428 21416 15434
rect 21364 15370 21416 15376
rect 28356 15428 28408 15434
rect 28356 15370 28408 15376
rect 12624 15360 12676 15366
rect 28368 15337 28396 15370
rect 28354 15328 28410 15337
rect 12676 15308 12756 15314
rect 12624 15302 12756 15308
rect 12636 15286 12756 15302
rect 12728 14346 12756 15286
rect 19656 15260 20032 15269
rect 19712 15258 19736 15260
rect 19792 15258 19816 15260
rect 19872 15258 19896 15260
rect 19952 15258 19976 15260
rect 19712 15206 19722 15258
rect 19966 15206 19976 15258
rect 19712 15204 19736 15206
rect 19792 15204 19816 15206
rect 19872 15204 19896 15206
rect 19952 15204 19976 15206
rect 19656 15195 20032 15204
rect 27656 15260 28032 15269
rect 28354 15263 28410 15272
rect 27712 15258 27736 15260
rect 27792 15258 27816 15260
rect 27872 15258 27896 15260
rect 27952 15258 27976 15260
rect 27712 15206 27722 15258
rect 27966 15206 27976 15258
rect 27712 15204 27736 15206
rect 27792 15204 27816 15206
rect 27872 15204 27896 15206
rect 27952 15204 27976 15206
rect 27656 15195 28032 15204
rect 28080 15020 28132 15026
rect 28080 14962 28132 14968
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12716 14340 12768 14346
rect 12716 14282 12768 14288
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12360 13530 12388 13874
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12176 12406 12296 12434
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 11656 11996 12032 12005
rect 11712 11994 11736 11996
rect 11792 11994 11816 11996
rect 11872 11994 11896 11996
rect 11952 11994 11976 11996
rect 11712 11942 11722 11994
rect 11966 11942 11976 11994
rect 11712 11940 11736 11942
rect 11792 11940 11816 11942
rect 11872 11940 11896 11942
rect 11952 11940 11976 11942
rect 11656 11931 12032 11940
rect 11704 11688 11756 11694
rect 11532 11648 11704 11676
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 10916 11452 11292 11461
rect 10972 11450 10996 11452
rect 11052 11450 11076 11452
rect 11132 11450 11156 11452
rect 11212 11450 11236 11452
rect 10972 11398 10982 11450
rect 11226 11398 11236 11450
rect 10972 11396 10996 11398
rect 11052 11396 11076 11398
rect 11132 11396 11156 11398
rect 11212 11396 11236 11398
rect 10916 11387 11292 11396
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11072 10810 11100 11086
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 11256 10554 11284 11154
rect 11348 10742 11376 11494
rect 11440 11218 11468 11562
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 1412 9897 1440 9998
rect 1584 9920 1636 9926
rect 1398 9888 1454 9897
rect 1584 9862 1636 9868
rect 1398 9823 1454 9832
rect 1596 9722 1624 9862
rect 3656 9820 4032 9829
rect 3712 9818 3736 9820
rect 3792 9818 3816 9820
rect 3872 9818 3896 9820
rect 3952 9818 3976 9820
rect 3712 9766 3722 9818
rect 3966 9766 3976 9818
rect 3712 9764 3736 9766
rect 3792 9764 3816 9766
rect 3872 9764 3896 9766
rect 3952 9764 3976 9766
rect 3656 9755 4032 9764
rect 1584 9716 1636 9722
rect 1584 9658 1636 9664
rect 10704 9654 10732 9998
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1412 9217 1440 9522
rect 10796 9518 10824 10542
rect 11256 10526 11376 10554
rect 10916 10364 11292 10373
rect 10972 10362 10996 10364
rect 11052 10362 11076 10364
rect 11132 10362 11156 10364
rect 11212 10362 11236 10364
rect 10972 10310 10982 10362
rect 11226 10310 11236 10362
rect 10972 10308 10996 10310
rect 11052 10308 11076 10310
rect 11132 10308 11156 10310
rect 11212 10308 11236 10310
rect 10916 10299 11292 10308
rect 11348 9926 11376 10526
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 2916 9276 3292 9285
rect 2972 9274 2996 9276
rect 3052 9274 3076 9276
rect 3132 9274 3156 9276
rect 3212 9274 3236 9276
rect 2972 9222 2982 9274
rect 3226 9222 3236 9274
rect 2972 9220 2996 9222
rect 3052 9220 3076 9222
rect 3132 9220 3156 9222
rect 3212 9220 3236 9222
rect 1398 9208 1454 9217
rect 2916 9211 3292 9220
rect 1398 9143 1454 9152
rect 3656 8732 4032 8741
rect 3712 8730 3736 8732
rect 3792 8730 3816 8732
rect 3872 8730 3896 8732
rect 3952 8730 3976 8732
rect 3712 8678 3722 8730
rect 3966 8678 3976 8730
rect 3712 8676 3736 8678
rect 3792 8676 3816 8678
rect 3872 8676 3896 8678
rect 3952 8676 3976 8678
rect 3656 8667 4032 8676
rect 10796 8634 10824 9318
rect 10916 9276 11292 9285
rect 10972 9274 10996 9276
rect 11052 9274 11076 9276
rect 11132 9274 11156 9276
rect 11212 9274 11236 9276
rect 10972 9222 10982 9274
rect 11226 9222 11236 9274
rect 10972 9220 10996 9222
rect 11052 9220 11076 9222
rect 11132 9220 11156 9222
rect 11212 9220 11236 9222
rect 10916 9211 11292 9220
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 1412 8401 1440 8434
rect 1398 8392 1454 8401
rect 1398 8327 1454 8336
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 2916 8188 3292 8197
rect 2972 8186 2996 8188
rect 3052 8186 3076 8188
rect 3132 8186 3156 8188
rect 3212 8186 3236 8188
rect 2972 8134 2982 8186
rect 3226 8134 3236 8186
rect 2972 8132 2996 8134
rect 3052 8132 3076 8134
rect 3132 8132 3156 8134
rect 3212 8132 3236 8134
rect 2916 8123 3292 8132
rect 10704 7954 10732 8230
rect 10916 8188 11292 8197
rect 10972 8186 10996 8188
rect 11052 8186 11076 8188
rect 11132 8186 11156 8188
rect 11212 8186 11236 8188
rect 10972 8134 10982 8186
rect 11226 8134 11236 8186
rect 10972 8132 10996 8134
rect 11052 8132 11076 8134
rect 11132 8132 11156 8134
rect 11212 8132 11236 8134
rect 10916 8123 11292 8132
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 7585 1440 7822
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 3656 7644 4032 7653
rect 3712 7642 3736 7644
rect 3792 7642 3816 7644
rect 3872 7642 3896 7644
rect 3952 7642 3976 7644
rect 3712 7590 3722 7642
rect 3966 7590 3976 7642
rect 3712 7588 3736 7590
rect 3792 7588 3816 7590
rect 3872 7588 3896 7590
rect 3952 7588 3976 7590
rect 1398 7576 1454 7585
rect 3656 7579 4032 7588
rect 1398 7511 1454 7520
rect 2916 7100 3292 7109
rect 2972 7098 2996 7100
rect 3052 7098 3076 7100
rect 3132 7098 3156 7100
rect 3212 7098 3236 7100
rect 2972 7046 2982 7098
rect 3226 7046 3236 7098
rect 2972 7044 2996 7046
rect 3052 7044 3076 7046
rect 3132 7044 3156 7046
rect 3212 7044 3236 7046
rect 2916 7035 3292 7044
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6497 1440 6734
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 3656 6556 4032 6565
rect 3712 6554 3736 6556
rect 3792 6554 3816 6556
rect 3872 6554 3896 6556
rect 3952 6554 3976 6556
rect 3712 6502 3722 6554
rect 3966 6502 3976 6554
rect 3712 6500 3736 6502
rect 3792 6500 3816 6502
rect 3872 6500 3896 6502
rect 3952 6500 3976 6502
rect 1398 6488 1454 6497
rect 3656 6491 4032 6500
rect 10060 6458 10088 6598
rect 10152 6458 10180 7686
rect 10704 6866 10732 7890
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10980 7546 11008 7754
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 11348 7478 11376 8434
rect 11440 8430 11468 10610
rect 11532 10538 11560 11648
rect 11704 11630 11756 11636
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 11656 10908 12032 10917
rect 11712 10906 11736 10908
rect 11792 10906 11816 10908
rect 11872 10906 11896 10908
rect 11952 10906 11976 10908
rect 11712 10854 11722 10906
rect 11966 10854 11976 10906
rect 11712 10852 11736 10854
rect 11792 10852 11816 10854
rect 11872 10852 11896 10854
rect 11952 10852 11976 10854
rect 11656 10843 12032 10852
rect 12084 10810 12112 11154
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 11520 10532 11572 10538
rect 11520 10474 11572 10480
rect 12072 10464 12124 10470
rect 11518 10432 11574 10441
rect 12072 10406 12124 10412
rect 11518 10367 11574 10376
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11336 7472 11388 7478
rect 11336 7414 11388 7420
rect 11440 7342 11468 8366
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 10916 7100 11292 7109
rect 10972 7098 10996 7100
rect 11052 7098 11076 7100
rect 11132 7098 11156 7100
rect 11212 7098 11236 7100
rect 10972 7046 10982 7098
rect 11226 7046 11236 7098
rect 10972 7044 10996 7046
rect 11052 7044 11076 7046
rect 11132 7044 11156 7046
rect 11212 7044 11236 7046
rect 10916 7035 11292 7044
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 1398 6423 1454 6432
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10704 6390 10732 6802
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 1412 5953 1440 6258
rect 2916 6012 3292 6021
rect 2972 6010 2996 6012
rect 3052 6010 3076 6012
rect 3132 6010 3156 6012
rect 3212 6010 3236 6012
rect 2972 5958 2982 6010
rect 3226 5958 3236 6010
rect 2972 5956 2996 5958
rect 3052 5956 3076 5958
rect 3132 5956 3156 5958
rect 3212 5956 3236 5958
rect 1398 5944 1454 5953
rect 2916 5947 3292 5956
rect 10152 5914 10180 6258
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 1398 5879 1454 5888
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 3656 5468 4032 5477
rect 3712 5466 3736 5468
rect 3792 5466 3816 5468
rect 3872 5466 3896 5468
rect 3952 5466 3976 5468
rect 3712 5414 3722 5466
rect 3966 5414 3976 5466
rect 3712 5412 3736 5414
rect 3792 5412 3816 5414
rect 3872 5412 3896 5414
rect 3952 5412 3976 5414
rect 3656 5403 4032 5412
rect 10428 5370 10456 6122
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10520 5846 10548 6054
rect 10508 5840 10560 5846
rect 10508 5782 10560 5788
rect 10704 5778 10732 6326
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10704 5658 10732 5714
rect 10612 5630 10732 5658
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 1398 5264 1454 5273
rect 1398 5199 1400 5208
rect 1452 5199 1454 5208
rect 1400 5170 1452 5176
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 2916 4924 3292 4933
rect 2972 4922 2996 4924
rect 3052 4922 3076 4924
rect 3132 4922 3156 4924
rect 3212 4922 3236 4924
rect 2972 4870 2982 4922
rect 3226 4870 3236 4922
rect 2972 4868 2996 4870
rect 3052 4868 3076 4870
rect 3132 4868 3156 4870
rect 3212 4868 3236 4870
rect 2916 4859 3292 4868
rect 7576 4826 7604 4966
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 10612 4690 10640 5630
rect 10796 5166 10824 6190
rect 10916 6012 11292 6021
rect 10972 6010 10996 6012
rect 11052 6010 11076 6012
rect 11132 6010 11156 6012
rect 11212 6010 11236 6012
rect 10972 5958 10982 6010
rect 11226 5958 11236 6010
rect 10972 5956 10996 5958
rect 11052 5956 11076 5958
rect 11132 5956 11156 5958
rect 11212 5956 11236 5958
rect 10916 5947 11292 5956
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1412 4321 1440 4558
rect 3656 4380 4032 4389
rect 3712 4378 3736 4380
rect 3792 4378 3816 4380
rect 3872 4378 3896 4380
rect 3952 4378 3976 4380
rect 3712 4326 3722 4378
rect 3966 4326 3976 4378
rect 3712 4324 3736 4326
rect 3792 4324 3816 4326
rect 3872 4324 3896 4326
rect 3952 4324 3976 4326
rect 1398 4312 1454 4321
rect 3656 4315 4032 4324
rect 1398 4247 1454 4256
rect 10612 4078 10640 4626
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 2916 3836 3292 3845
rect 2972 3834 2996 3836
rect 3052 3834 3076 3836
rect 3132 3834 3156 3836
rect 3212 3834 3236 3836
rect 2972 3782 2982 3834
rect 3226 3782 3236 3834
rect 2972 3780 2996 3782
rect 3052 3780 3076 3782
rect 3132 3780 3156 3782
rect 3212 3780 3236 3782
rect 2916 3771 3292 3780
rect 10612 3602 10640 4014
rect 10796 3754 10824 5102
rect 10916 4924 11292 4933
rect 10972 4922 10996 4924
rect 11052 4922 11076 4924
rect 11132 4922 11156 4924
rect 11212 4922 11236 4924
rect 10972 4870 10982 4922
rect 11226 4870 11236 4922
rect 10972 4868 10996 4870
rect 11052 4868 11076 4870
rect 11132 4868 11156 4870
rect 11212 4868 11236 4870
rect 10916 4859 11292 4868
rect 11440 4146 11468 7278
rect 11532 5114 11560 10367
rect 11656 9820 12032 9829
rect 11712 9818 11736 9820
rect 11792 9818 11816 9820
rect 11872 9818 11896 9820
rect 11952 9818 11976 9820
rect 11712 9766 11722 9818
rect 11966 9766 11976 9818
rect 11712 9764 11736 9766
rect 11792 9764 11816 9766
rect 11872 9764 11896 9766
rect 11952 9764 11976 9766
rect 11656 9755 12032 9764
rect 12084 8974 12112 10406
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 11656 8732 12032 8741
rect 11712 8730 11736 8732
rect 11792 8730 11816 8732
rect 11872 8730 11896 8732
rect 11952 8730 11976 8732
rect 11712 8678 11722 8730
rect 11966 8678 11976 8730
rect 11712 8676 11736 8678
rect 11792 8676 11816 8678
rect 11872 8676 11896 8678
rect 11952 8676 11976 8678
rect 11656 8667 12032 8676
rect 12084 8566 12112 8910
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 12084 7886 12112 8502
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 11656 7644 12032 7653
rect 11712 7642 11736 7644
rect 11792 7642 11816 7644
rect 11872 7642 11896 7644
rect 11952 7642 11976 7644
rect 11712 7590 11722 7642
rect 11966 7590 11976 7642
rect 11712 7588 11736 7590
rect 11792 7588 11816 7590
rect 11872 7588 11896 7590
rect 11952 7588 11976 7590
rect 11656 7579 12032 7588
rect 11656 6556 12032 6565
rect 11712 6554 11736 6556
rect 11792 6554 11816 6556
rect 11872 6554 11896 6556
rect 11952 6554 11976 6556
rect 11712 6502 11722 6554
rect 11966 6502 11976 6554
rect 11712 6500 11736 6502
rect 11792 6500 11816 6502
rect 11872 6500 11896 6502
rect 11952 6500 11976 6502
rect 11656 6491 12032 6500
rect 11656 5468 12032 5477
rect 11712 5466 11736 5468
rect 11792 5466 11816 5468
rect 11872 5466 11896 5468
rect 11952 5466 11976 5468
rect 11712 5414 11722 5466
rect 11966 5414 11976 5466
rect 11712 5412 11736 5414
rect 11792 5412 11816 5414
rect 11872 5412 11896 5414
rect 11952 5412 11976 5414
rect 11656 5403 12032 5412
rect 11532 5086 11652 5114
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11532 4690 11560 4966
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11624 4468 11652 5086
rect 11532 4440 11652 4468
rect 11532 4214 11560 4440
rect 11656 4380 12032 4389
rect 11712 4378 11736 4380
rect 11792 4378 11816 4380
rect 11872 4378 11896 4380
rect 11952 4378 11976 4380
rect 11712 4326 11722 4378
rect 11966 4326 11976 4378
rect 11712 4324 11736 4326
rect 11792 4324 11816 4326
rect 11872 4324 11896 4326
rect 11952 4324 11976 4326
rect 11656 4315 12032 4324
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 10916 3836 11292 3845
rect 10972 3834 10996 3836
rect 11052 3834 11076 3836
rect 11132 3834 11156 3836
rect 11212 3834 11236 3836
rect 10972 3782 10982 3834
rect 11226 3782 11236 3834
rect 10972 3780 10996 3782
rect 11052 3780 11076 3782
rect 11132 3780 11156 3782
rect 11212 3780 11236 3782
rect 10916 3771 11292 3780
rect 10704 3738 10824 3754
rect 10692 3732 10824 3738
rect 10744 3726 10824 3732
rect 10692 3674 10744 3680
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 1400 3528 1452 3534
rect 1398 3496 1400 3505
rect 1452 3496 1454 3505
rect 1398 3431 1454 3440
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 3656 3292 4032 3301
rect 3712 3290 3736 3292
rect 3792 3290 3816 3292
rect 3872 3290 3896 3292
rect 3952 3290 3976 3292
rect 3712 3238 3722 3290
rect 3966 3238 3976 3290
rect 3712 3236 3736 3238
rect 3792 3236 3816 3238
rect 3872 3236 3896 3238
rect 3952 3236 3976 3238
rect 3656 3227 4032 3236
rect 10244 3194 10272 3334
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10612 3126 10640 3538
rect 10600 3120 10652 3126
rect 10600 3062 10652 3068
rect 848 3052 900 3058
rect 848 2994 900 3000
rect 860 2689 888 2994
rect 10704 2990 10732 3674
rect 11440 3482 11468 4082
rect 11164 3466 11468 3482
rect 11152 3460 11468 3466
rect 11204 3454 11468 3460
rect 11152 3402 11204 3408
rect 11532 3194 11560 4150
rect 12176 3398 12204 12406
rect 12360 12322 12388 13194
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12268 12294 12388 12322
rect 12268 10470 12296 12294
rect 12452 12186 12480 12854
rect 12636 12782 12664 13126
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12360 12170 12480 12186
rect 12348 12164 12480 12170
rect 12400 12158 12480 12164
rect 12348 12106 12400 12112
rect 12452 11830 12480 12158
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12452 11234 12480 11766
rect 12820 11694 12848 14758
rect 18916 14716 19292 14725
rect 18972 14714 18996 14716
rect 19052 14714 19076 14716
rect 19132 14714 19156 14716
rect 19212 14714 19236 14716
rect 18972 14662 18982 14714
rect 19226 14662 19236 14714
rect 18972 14660 18996 14662
rect 19052 14660 19076 14662
rect 19132 14660 19156 14662
rect 19212 14660 19236 14662
rect 18916 14651 19292 14660
rect 26916 14716 27292 14725
rect 26972 14714 26996 14716
rect 27052 14714 27076 14716
rect 27132 14714 27156 14716
rect 27212 14714 27236 14716
rect 26972 14662 26982 14714
rect 27226 14662 27236 14714
rect 26972 14660 26996 14662
rect 27052 14660 27076 14662
rect 27132 14660 27156 14662
rect 27212 14660 27236 14662
rect 26916 14651 27292 14660
rect 28092 14278 28120 14962
rect 28356 14952 28408 14958
rect 28356 14894 28408 14900
rect 28368 14521 28396 14894
rect 28354 14512 28410 14521
rect 28354 14447 28410 14456
rect 28080 14272 28132 14278
rect 28080 14214 28132 14220
rect 19656 14172 20032 14181
rect 19712 14170 19736 14172
rect 19792 14170 19816 14172
rect 19872 14170 19896 14172
rect 19952 14170 19976 14172
rect 19712 14118 19722 14170
rect 19966 14118 19976 14170
rect 19712 14116 19736 14118
rect 19792 14116 19816 14118
rect 19872 14116 19896 14118
rect 19952 14116 19976 14118
rect 19656 14107 20032 14116
rect 27656 14172 28032 14181
rect 27712 14170 27736 14172
rect 27792 14170 27816 14172
rect 27872 14170 27896 14172
rect 27952 14170 27976 14172
rect 27712 14118 27722 14170
rect 27966 14118 27976 14170
rect 27712 14116 27736 14118
rect 27792 14116 27816 14118
rect 27872 14116 27896 14118
rect 27952 14116 27976 14118
rect 27656 14107 28032 14116
rect 28356 13864 28408 13870
rect 28356 13806 28408 13812
rect 28368 13705 28396 13806
rect 28354 13696 28410 13705
rect 18916 13628 19292 13637
rect 18972 13626 18996 13628
rect 19052 13626 19076 13628
rect 19132 13626 19156 13628
rect 19212 13626 19236 13628
rect 18972 13574 18982 13626
rect 19226 13574 19236 13626
rect 18972 13572 18996 13574
rect 19052 13572 19076 13574
rect 19132 13572 19156 13574
rect 19212 13572 19236 13574
rect 18916 13563 19292 13572
rect 26916 13628 27292 13637
rect 28354 13631 28410 13640
rect 26972 13626 26996 13628
rect 27052 13626 27076 13628
rect 27132 13626 27156 13628
rect 27212 13626 27236 13628
rect 26972 13574 26982 13626
rect 27226 13574 27236 13626
rect 26972 13572 26996 13574
rect 27052 13572 27076 13574
rect 27132 13572 27156 13574
rect 27212 13572 27236 13574
rect 26916 13563 27292 13572
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13372 12986 13400 13262
rect 28356 13252 28408 13258
rect 28356 13194 28408 13200
rect 19656 13084 20032 13093
rect 19712 13082 19736 13084
rect 19792 13082 19816 13084
rect 19872 13082 19896 13084
rect 19952 13082 19976 13084
rect 19712 13030 19722 13082
rect 19966 13030 19976 13082
rect 19712 13028 19736 13030
rect 19792 13028 19816 13030
rect 19872 13028 19896 13030
rect 19952 13028 19976 13030
rect 19656 13019 20032 13028
rect 27656 13084 28032 13093
rect 27712 13082 27736 13084
rect 27792 13082 27816 13084
rect 27872 13082 27896 13084
rect 27952 13082 27976 13084
rect 27712 13030 27722 13082
rect 27966 13030 27976 13082
rect 27712 13028 27736 13030
rect 27792 13028 27816 13030
rect 27872 13028 27896 13030
rect 27952 13028 27976 13030
rect 27656 13019 28032 13028
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 28368 12889 28396 13194
rect 28354 12880 28410 12889
rect 28354 12815 28410 12824
rect 18916 12540 19292 12549
rect 18972 12538 18996 12540
rect 19052 12538 19076 12540
rect 19132 12538 19156 12540
rect 19212 12538 19236 12540
rect 18972 12486 18982 12538
rect 19226 12486 19236 12538
rect 18972 12484 18996 12486
rect 19052 12484 19076 12486
rect 19132 12484 19156 12486
rect 19212 12484 19236 12486
rect 18916 12475 19292 12484
rect 26916 12540 27292 12549
rect 26972 12538 26996 12540
rect 27052 12538 27076 12540
rect 27132 12538 27156 12540
rect 27212 12538 27236 12540
rect 26972 12486 26982 12538
rect 27226 12486 27236 12538
rect 26972 12484 26996 12486
rect 27052 12484 27076 12486
rect 27132 12484 27156 12486
rect 27212 12484 27236 12486
rect 26916 12475 27292 12484
rect 28356 12164 28408 12170
rect 28356 12106 28408 12112
rect 28368 12073 28396 12106
rect 28354 12064 28410 12073
rect 19656 11996 20032 12005
rect 19712 11994 19736 11996
rect 19792 11994 19816 11996
rect 19872 11994 19896 11996
rect 19952 11994 19976 11996
rect 19712 11942 19722 11994
rect 19966 11942 19976 11994
rect 19712 11940 19736 11942
rect 19792 11940 19816 11942
rect 19872 11940 19896 11942
rect 19952 11940 19976 11942
rect 19656 11931 20032 11940
rect 27656 11996 28032 12005
rect 28354 11999 28410 12008
rect 27712 11994 27736 11996
rect 27792 11994 27816 11996
rect 27872 11994 27896 11996
rect 27952 11994 27976 11996
rect 27712 11942 27722 11994
rect 27966 11942 27976 11994
rect 27712 11940 27736 11942
rect 27792 11940 27816 11942
rect 27872 11940 27896 11942
rect 27952 11940 27976 11942
rect 27656 11931 28032 11940
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 28356 11688 28408 11694
rect 28356 11630 28408 11636
rect 12360 11206 12480 11234
rect 12360 11082 12388 11206
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12360 9994 12388 11018
rect 12452 10674 12480 11018
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 12360 9874 12388 9930
rect 12268 9846 12388 9874
rect 12268 9654 12296 9846
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 12268 9178 12296 9590
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 12268 5642 12296 6326
rect 12256 5636 12308 5642
rect 12256 5578 12308 5584
rect 12268 4690 12296 5578
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12268 4214 12296 4626
rect 12256 4208 12308 4214
rect 12256 4150 12308 4156
rect 12268 3466 12296 4150
rect 12360 3466 12388 7822
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 12452 7546 12480 7686
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12820 6798 12848 11630
rect 18916 11452 19292 11461
rect 18972 11450 18996 11452
rect 19052 11450 19076 11452
rect 19132 11450 19156 11452
rect 19212 11450 19236 11452
rect 18972 11398 18982 11450
rect 19226 11398 19236 11450
rect 18972 11396 18996 11398
rect 19052 11396 19076 11398
rect 19132 11396 19156 11398
rect 19212 11396 19236 11398
rect 18916 11387 19292 11396
rect 26916 11452 27292 11461
rect 26972 11450 26996 11452
rect 27052 11450 27076 11452
rect 27132 11450 27156 11452
rect 27212 11450 27236 11452
rect 26972 11398 26982 11450
rect 27226 11398 27236 11450
rect 26972 11396 26996 11398
rect 27052 11396 27076 11398
rect 27132 11396 27156 11398
rect 27212 11396 27236 11398
rect 26916 11387 27292 11396
rect 28368 11257 28396 11630
rect 28354 11248 28410 11257
rect 28354 11183 28410 11192
rect 19656 10908 20032 10917
rect 19712 10906 19736 10908
rect 19792 10906 19816 10908
rect 19872 10906 19896 10908
rect 19952 10906 19976 10908
rect 19712 10854 19722 10906
rect 19966 10854 19976 10906
rect 19712 10852 19736 10854
rect 19792 10852 19816 10854
rect 19872 10852 19896 10854
rect 19952 10852 19976 10854
rect 19656 10843 20032 10852
rect 27656 10908 28032 10917
rect 27712 10906 27736 10908
rect 27792 10906 27816 10908
rect 27872 10906 27896 10908
rect 27952 10906 27976 10908
rect 27712 10854 27722 10906
rect 27966 10854 27976 10906
rect 27712 10852 27736 10854
rect 27792 10852 27816 10854
rect 27872 10852 27896 10854
rect 27952 10852 27976 10854
rect 27656 10843 28032 10852
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 28356 10600 28408 10606
rect 28356 10542 28408 10548
rect 13188 10130 13216 10542
rect 28368 10441 28396 10542
rect 28354 10432 28410 10441
rect 18916 10364 19292 10373
rect 18972 10362 18996 10364
rect 19052 10362 19076 10364
rect 19132 10362 19156 10364
rect 19212 10362 19236 10364
rect 18972 10310 18982 10362
rect 19226 10310 19236 10362
rect 18972 10308 18996 10310
rect 19052 10308 19076 10310
rect 19132 10308 19156 10310
rect 19212 10308 19236 10310
rect 18916 10299 19292 10308
rect 26916 10364 27292 10373
rect 28354 10367 28410 10376
rect 26972 10362 26996 10364
rect 27052 10362 27076 10364
rect 27132 10362 27156 10364
rect 27212 10362 27236 10364
rect 26972 10310 26982 10362
rect 27226 10310 27236 10362
rect 26972 10308 26996 10310
rect 27052 10308 27076 10310
rect 27132 10308 27156 10310
rect 27212 10308 27236 10310
rect 26916 10299 27292 10308
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 28356 9988 28408 9994
rect 28356 9930 28408 9936
rect 19656 9820 20032 9829
rect 19712 9818 19736 9820
rect 19792 9818 19816 9820
rect 19872 9818 19896 9820
rect 19952 9818 19976 9820
rect 19712 9766 19722 9818
rect 19966 9766 19976 9818
rect 19712 9764 19736 9766
rect 19792 9764 19816 9766
rect 19872 9764 19896 9766
rect 19952 9764 19976 9766
rect 19656 9755 20032 9764
rect 27656 9820 28032 9829
rect 27712 9818 27736 9820
rect 27792 9818 27816 9820
rect 27872 9818 27896 9820
rect 27952 9818 27976 9820
rect 27712 9766 27722 9818
rect 27966 9766 27976 9818
rect 27712 9764 27736 9766
rect 27792 9764 27816 9766
rect 27872 9764 27896 9766
rect 27952 9764 27976 9766
rect 27656 9755 28032 9764
rect 28368 9625 28396 9930
rect 28354 9616 28410 9625
rect 28354 9551 28410 9560
rect 28080 9376 28132 9382
rect 28080 9318 28132 9324
rect 18916 9276 19292 9285
rect 18972 9274 18996 9276
rect 19052 9274 19076 9276
rect 19132 9274 19156 9276
rect 19212 9274 19236 9276
rect 18972 9222 18982 9274
rect 19226 9222 19236 9274
rect 18972 9220 18996 9222
rect 19052 9220 19076 9222
rect 19132 9220 19156 9222
rect 19212 9220 19236 9222
rect 18916 9211 19292 9220
rect 26916 9276 27292 9285
rect 26972 9274 26996 9276
rect 27052 9274 27076 9276
rect 27132 9274 27156 9276
rect 27212 9274 27236 9276
rect 26972 9222 26982 9274
rect 27226 9222 27236 9274
rect 26972 9220 26996 9222
rect 27052 9220 27076 9222
rect 27132 9220 27156 9222
rect 27212 9220 27236 9222
rect 26916 9211 27292 9220
rect 28092 8974 28120 9318
rect 28080 8968 28132 8974
rect 28080 8910 28132 8916
rect 28356 8900 28408 8906
rect 28356 8842 28408 8848
rect 28368 8809 28396 8842
rect 28354 8800 28410 8809
rect 19656 8732 20032 8741
rect 19712 8730 19736 8732
rect 19792 8730 19816 8732
rect 19872 8730 19896 8732
rect 19952 8730 19976 8732
rect 19712 8678 19722 8730
rect 19966 8678 19976 8730
rect 19712 8676 19736 8678
rect 19792 8676 19816 8678
rect 19872 8676 19896 8678
rect 19952 8676 19976 8678
rect 19656 8667 20032 8676
rect 27656 8732 28032 8741
rect 28354 8735 28410 8744
rect 27712 8730 27736 8732
rect 27792 8730 27816 8732
rect 27872 8730 27896 8732
rect 27952 8730 27976 8732
rect 27712 8678 27722 8730
rect 27966 8678 27976 8730
rect 27712 8676 27736 8678
rect 27792 8676 27816 8678
rect 27872 8676 27896 8678
rect 27952 8676 27976 8678
rect 27656 8667 28032 8676
rect 28356 8424 28408 8430
rect 28356 8366 28408 8372
rect 18916 8188 19292 8197
rect 18972 8186 18996 8188
rect 19052 8186 19076 8188
rect 19132 8186 19156 8188
rect 19212 8186 19236 8188
rect 18972 8134 18982 8186
rect 19226 8134 19236 8186
rect 18972 8132 18996 8134
rect 19052 8132 19076 8134
rect 19132 8132 19156 8134
rect 19212 8132 19236 8134
rect 18916 8123 19292 8132
rect 26916 8188 27292 8197
rect 26972 8186 26996 8188
rect 27052 8186 27076 8188
rect 27132 8186 27156 8188
rect 27212 8186 27236 8188
rect 26972 8134 26982 8186
rect 27226 8134 27236 8186
rect 26972 8132 26996 8134
rect 27052 8132 27076 8134
rect 27132 8132 27156 8134
rect 27212 8132 27236 8134
rect 26916 8123 27292 8132
rect 28368 7993 28396 8366
rect 28354 7984 28410 7993
rect 28354 7919 28410 7928
rect 28080 7744 28132 7750
rect 28080 7686 28132 7692
rect 19656 7644 20032 7653
rect 19712 7642 19736 7644
rect 19792 7642 19816 7644
rect 19872 7642 19896 7644
rect 19952 7642 19976 7644
rect 19712 7590 19722 7642
rect 19966 7590 19976 7642
rect 19712 7588 19736 7590
rect 19792 7588 19816 7590
rect 19872 7588 19896 7590
rect 19952 7588 19976 7590
rect 19656 7579 20032 7588
rect 27656 7644 28032 7653
rect 27712 7642 27736 7644
rect 27792 7642 27816 7644
rect 27872 7642 27896 7644
rect 27952 7642 27976 7644
rect 27712 7590 27722 7642
rect 27966 7590 27976 7642
rect 27712 7588 27736 7590
rect 27792 7588 27816 7590
rect 27872 7588 27896 7590
rect 27952 7588 27976 7590
rect 27656 7579 28032 7588
rect 28092 7410 28120 7686
rect 28080 7404 28132 7410
rect 28080 7346 28132 7352
rect 28356 7336 28408 7342
rect 28356 7278 28408 7284
rect 28368 7177 28396 7278
rect 28354 7168 28410 7177
rect 18916 7100 19292 7109
rect 18972 7098 18996 7100
rect 19052 7098 19076 7100
rect 19132 7098 19156 7100
rect 19212 7098 19236 7100
rect 18972 7046 18982 7098
rect 19226 7046 19236 7098
rect 18972 7044 18996 7046
rect 19052 7044 19076 7046
rect 19132 7044 19156 7046
rect 19212 7044 19236 7046
rect 18916 7035 19292 7044
rect 26916 7100 27292 7109
rect 28354 7103 28410 7112
rect 26972 7098 26996 7100
rect 27052 7098 27076 7100
rect 27132 7098 27156 7100
rect 27212 7098 27236 7100
rect 26972 7046 26982 7098
rect 27226 7046 27236 7098
rect 26972 7044 26996 7046
rect 27052 7044 27076 7046
rect 27132 7044 27156 7046
rect 27212 7044 27236 7046
rect 26916 7035 27292 7044
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 28080 6792 28132 6798
rect 28080 6734 28132 6740
rect 19656 6556 20032 6565
rect 19712 6554 19736 6556
rect 19792 6554 19816 6556
rect 19872 6554 19896 6556
rect 19952 6554 19976 6556
rect 19712 6502 19722 6554
rect 19966 6502 19976 6554
rect 19712 6500 19736 6502
rect 19792 6500 19816 6502
rect 19872 6500 19896 6502
rect 19952 6500 19976 6502
rect 19656 6491 20032 6500
rect 27656 6556 28032 6565
rect 27712 6554 27736 6556
rect 27792 6554 27816 6556
rect 27872 6554 27896 6556
rect 27952 6554 27976 6556
rect 27712 6502 27722 6554
rect 27966 6502 27976 6554
rect 27712 6500 27736 6502
rect 27792 6500 27816 6502
rect 27872 6500 27896 6502
rect 27952 6500 27976 6502
rect 27656 6491 28032 6500
rect 28092 6118 28120 6734
rect 28356 6724 28408 6730
rect 28356 6666 28408 6672
rect 28368 6361 28396 6666
rect 28354 6352 28410 6361
rect 28354 6287 28410 6296
rect 28080 6112 28132 6118
rect 28080 6054 28132 6060
rect 18916 6012 19292 6021
rect 18972 6010 18996 6012
rect 19052 6010 19076 6012
rect 19132 6010 19156 6012
rect 19212 6010 19236 6012
rect 18972 5958 18982 6010
rect 19226 5958 19236 6010
rect 18972 5956 18996 5958
rect 19052 5956 19076 5958
rect 19132 5956 19156 5958
rect 19212 5956 19236 5958
rect 18916 5947 19292 5956
rect 26916 6012 27292 6021
rect 26972 6010 26996 6012
rect 27052 6010 27076 6012
rect 27132 6010 27156 6012
rect 27212 6010 27236 6012
rect 26972 5958 26982 6010
rect 27226 5958 27236 6010
rect 26972 5956 26996 5958
rect 27052 5956 27076 5958
rect 27132 5956 27156 5958
rect 27212 5956 27236 5958
rect 26916 5947 27292 5956
rect 28356 5636 28408 5642
rect 28356 5578 28408 5584
rect 28368 5545 28396 5578
rect 28354 5536 28410 5545
rect 19656 5468 20032 5477
rect 19712 5466 19736 5468
rect 19792 5466 19816 5468
rect 19872 5466 19896 5468
rect 19952 5466 19976 5468
rect 19712 5414 19722 5466
rect 19966 5414 19976 5466
rect 19712 5412 19736 5414
rect 19792 5412 19816 5414
rect 19872 5412 19896 5414
rect 19952 5412 19976 5414
rect 19656 5403 20032 5412
rect 27656 5468 28032 5477
rect 28354 5471 28410 5480
rect 27712 5466 27736 5468
rect 27792 5466 27816 5468
rect 27872 5466 27896 5468
rect 27952 5466 27976 5468
rect 27712 5414 27722 5466
rect 27966 5414 27976 5466
rect 27712 5412 27736 5414
rect 27792 5412 27816 5414
rect 27872 5412 27896 5414
rect 27952 5412 27976 5414
rect 27656 5403 28032 5412
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 28080 5228 28132 5234
rect 28080 5170 28132 5176
rect 12544 4554 12572 5170
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 13004 4690 13032 5102
rect 18916 4924 19292 4933
rect 18972 4922 18996 4924
rect 19052 4922 19076 4924
rect 19132 4922 19156 4924
rect 19212 4922 19236 4924
rect 18972 4870 18982 4922
rect 19226 4870 19236 4922
rect 18972 4868 18996 4870
rect 19052 4868 19076 4870
rect 19132 4868 19156 4870
rect 19212 4868 19236 4870
rect 18916 4859 19292 4868
rect 26916 4924 27292 4933
rect 26972 4922 26996 4924
rect 27052 4922 27076 4924
rect 27132 4922 27156 4924
rect 27212 4922 27236 4924
rect 26972 4870 26982 4922
rect 27226 4870 27236 4922
rect 26972 4868 26996 4870
rect 27052 4868 27076 4870
rect 27132 4868 27156 4870
rect 27212 4868 27236 4870
rect 26916 4859 27292 4868
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12532 4548 12584 4554
rect 12532 4490 12584 4496
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12452 4078 12480 4422
rect 12544 4282 12572 4490
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12728 3602 12756 4558
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12820 4078 12848 4422
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 13004 3602 13032 4626
rect 19656 4380 20032 4389
rect 19712 4378 19736 4380
rect 19792 4378 19816 4380
rect 19872 4378 19896 4380
rect 19952 4378 19976 4380
rect 19712 4326 19722 4378
rect 19966 4326 19976 4378
rect 19712 4324 19736 4326
rect 19792 4324 19816 4326
rect 19872 4324 19896 4326
rect 19952 4324 19976 4326
rect 19656 4315 20032 4324
rect 27656 4380 28032 4389
rect 27712 4378 27736 4380
rect 27792 4378 27816 4380
rect 27872 4378 27896 4380
rect 27952 4378 27976 4380
rect 27712 4326 27722 4378
rect 27966 4326 27976 4378
rect 27712 4324 27736 4326
rect 27792 4324 27816 4326
rect 27872 4324 27896 4326
rect 27952 4324 27976 4326
rect 27656 4315 28032 4324
rect 28092 4282 28120 5170
rect 28356 5160 28408 5166
rect 28356 5102 28408 5108
rect 28368 4729 28396 5102
rect 28354 4720 28410 4729
rect 28354 4655 28410 4664
rect 28080 4276 28132 4282
rect 28080 4218 28132 4224
rect 28356 4072 28408 4078
rect 28356 4014 28408 4020
rect 28368 3913 28396 4014
rect 28354 3904 28410 3913
rect 18916 3836 19292 3845
rect 18972 3834 18996 3836
rect 19052 3834 19076 3836
rect 19132 3834 19156 3836
rect 19212 3834 19236 3836
rect 18972 3782 18982 3834
rect 19226 3782 19236 3834
rect 18972 3780 18996 3782
rect 19052 3780 19076 3782
rect 19132 3780 19156 3782
rect 19212 3780 19236 3782
rect 18916 3771 19292 3780
rect 26916 3836 27292 3845
rect 28354 3839 28410 3848
rect 26972 3834 26996 3836
rect 27052 3834 27076 3836
rect 27132 3834 27156 3836
rect 27212 3834 27236 3836
rect 26972 3782 26982 3834
rect 27226 3782 27236 3834
rect 26972 3780 26996 3782
rect 27052 3780 27076 3782
rect 27132 3780 27156 3782
rect 27212 3780 27236 3782
rect 26916 3771 27292 3780
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 12256 3460 12308 3466
rect 12256 3402 12308 3408
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 28356 3460 28408 3466
rect 28356 3402 28408 3408
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 11656 3292 12032 3301
rect 11712 3290 11736 3292
rect 11792 3290 11816 3292
rect 11872 3290 11896 3292
rect 11952 3290 11976 3292
rect 11712 3238 11722 3290
rect 11966 3238 11976 3290
rect 11712 3236 11736 3238
rect 11792 3236 11816 3238
rect 11872 3236 11896 3238
rect 11952 3236 11976 3238
rect 11656 3227 12032 3236
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 10692 2984 10744 2990
rect 11072 2938 11100 3130
rect 10692 2926 10744 2932
rect 10888 2910 11100 2938
rect 10888 2854 10916 2910
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 2916 2748 3292 2757
rect 2972 2746 2996 2748
rect 3052 2746 3076 2748
rect 3132 2746 3156 2748
rect 3212 2746 3236 2748
rect 2972 2694 2982 2746
rect 3226 2694 3236 2746
rect 2972 2692 2996 2694
rect 3052 2692 3076 2694
rect 3132 2692 3156 2694
rect 3212 2692 3236 2694
rect 846 2680 902 2689
rect 2916 2683 3292 2692
rect 10916 2748 11292 2757
rect 10972 2746 10996 2748
rect 11052 2746 11076 2748
rect 11132 2746 11156 2748
rect 11212 2746 11236 2748
rect 10972 2694 10982 2746
rect 11226 2694 11236 2746
rect 10972 2692 10996 2694
rect 11052 2692 11076 2694
rect 11132 2692 11156 2694
rect 11212 2692 11236 2694
rect 10916 2683 11292 2692
rect 846 2615 902 2624
rect 848 2440 900 2446
rect 848 2382 900 2388
rect 860 1873 888 2382
rect 12176 2310 12204 3334
rect 12268 3126 12296 3402
rect 12256 3120 12308 3126
rect 12256 3062 12308 3068
rect 12268 2650 12296 3062
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12360 2446 12388 3402
rect 19656 3292 20032 3301
rect 19712 3290 19736 3292
rect 19792 3290 19816 3292
rect 19872 3290 19896 3292
rect 19952 3290 19976 3292
rect 19712 3238 19722 3290
rect 19966 3238 19976 3290
rect 19712 3236 19736 3238
rect 19792 3236 19816 3238
rect 19872 3236 19896 3238
rect 19952 3236 19976 3238
rect 19656 3227 20032 3236
rect 27656 3292 28032 3301
rect 27712 3290 27736 3292
rect 27792 3290 27816 3292
rect 27872 3290 27896 3292
rect 27952 3290 27976 3292
rect 27712 3238 27722 3290
rect 27966 3238 27976 3290
rect 27712 3236 27736 3238
rect 27792 3236 27816 3238
rect 27872 3236 27896 3238
rect 27952 3236 27976 3238
rect 27656 3227 28032 3236
rect 28368 3097 28396 3402
rect 28354 3088 28410 3097
rect 28354 3023 28410 3032
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 18916 2748 19292 2757
rect 18972 2746 18996 2748
rect 19052 2746 19076 2748
rect 19132 2746 19156 2748
rect 19212 2746 19236 2748
rect 18972 2694 18982 2746
rect 19226 2694 19236 2746
rect 18972 2692 18996 2694
rect 19052 2692 19076 2694
rect 19132 2692 19156 2694
rect 19212 2692 19236 2694
rect 18916 2683 19292 2692
rect 20640 2446 20668 2790
rect 26916 2748 27292 2757
rect 26972 2746 26996 2748
rect 27052 2746 27076 2748
rect 27132 2746 27156 2748
rect 27212 2746 27236 2748
rect 26972 2694 26982 2746
rect 27226 2694 27236 2746
rect 26972 2692 26996 2694
rect 27052 2692 27076 2694
rect 27132 2692 27156 2694
rect 27212 2692 27236 2694
rect 26916 2683 27292 2692
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 28356 2372 28408 2378
rect 28356 2314 28408 2320
rect 12164 2304 12216 2310
rect 28368 2281 28396 2314
rect 12164 2246 12216 2252
rect 28354 2272 28410 2281
rect 3656 2204 4032 2213
rect 3712 2202 3736 2204
rect 3792 2202 3816 2204
rect 3872 2202 3896 2204
rect 3952 2202 3976 2204
rect 3712 2150 3722 2202
rect 3966 2150 3976 2202
rect 3712 2148 3736 2150
rect 3792 2148 3816 2150
rect 3872 2148 3896 2150
rect 3952 2148 3976 2150
rect 3656 2139 4032 2148
rect 11656 2204 12032 2213
rect 11712 2202 11736 2204
rect 11792 2202 11816 2204
rect 11872 2202 11896 2204
rect 11952 2202 11976 2204
rect 11712 2150 11722 2202
rect 11966 2150 11976 2202
rect 11712 2148 11736 2150
rect 11792 2148 11816 2150
rect 11872 2148 11896 2150
rect 11952 2148 11976 2150
rect 11656 2139 12032 2148
rect 19656 2204 20032 2213
rect 19712 2202 19736 2204
rect 19792 2202 19816 2204
rect 19872 2202 19896 2204
rect 19952 2202 19976 2204
rect 19712 2150 19722 2202
rect 19966 2150 19976 2202
rect 19712 2148 19736 2150
rect 19792 2148 19816 2150
rect 19872 2148 19896 2150
rect 19952 2148 19976 2150
rect 19656 2139 20032 2148
rect 27656 2204 28032 2213
rect 28354 2207 28410 2216
rect 27712 2202 27736 2204
rect 27792 2202 27816 2204
rect 27872 2202 27896 2204
rect 27952 2202 27976 2204
rect 27712 2150 27722 2202
rect 27966 2150 27976 2202
rect 27712 2148 27736 2150
rect 27792 2148 27816 2150
rect 27872 2148 27896 2150
rect 27952 2148 27976 2150
rect 27656 2139 28032 2148
rect 846 1864 902 1873
rect 846 1799 902 1808
rect 110 1184 166 1193
rect 110 1119 166 1128
<< via2 >>
rect 1030 28600 1086 28656
rect 938 27784 994 27840
rect 2916 27770 2972 27772
rect 2996 27770 3052 27772
rect 3076 27770 3132 27772
rect 3156 27770 3212 27772
rect 3236 27770 3292 27772
rect 2916 27718 2918 27770
rect 2918 27718 2970 27770
rect 2970 27718 2972 27770
rect 2996 27718 3034 27770
rect 3034 27718 3046 27770
rect 3046 27718 3052 27770
rect 3076 27718 3098 27770
rect 3098 27718 3110 27770
rect 3110 27718 3132 27770
rect 3156 27718 3162 27770
rect 3162 27718 3174 27770
rect 3174 27718 3212 27770
rect 3236 27718 3238 27770
rect 3238 27718 3290 27770
rect 3290 27718 3292 27770
rect 2916 27716 2972 27718
rect 2996 27716 3052 27718
rect 3076 27716 3132 27718
rect 3156 27716 3212 27718
rect 3236 27716 3292 27718
rect 10916 27770 10972 27772
rect 10996 27770 11052 27772
rect 11076 27770 11132 27772
rect 11156 27770 11212 27772
rect 11236 27770 11292 27772
rect 10916 27718 10918 27770
rect 10918 27718 10970 27770
rect 10970 27718 10972 27770
rect 10996 27718 11034 27770
rect 11034 27718 11046 27770
rect 11046 27718 11052 27770
rect 11076 27718 11098 27770
rect 11098 27718 11110 27770
rect 11110 27718 11132 27770
rect 11156 27718 11162 27770
rect 11162 27718 11174 27770
rect 11174 27718 11212 27770
rect 11236 27718 11238 27770
rect 11238 27718 11290 27770
rect 11290 27718 11292 27770
rect 10916 27716 10972 27718
rect 10996 27716 11052 27718
rect 11076 27716 11132 27718
rect 11156 27716 11212 27718
rect 11236 27716 11292 27718
rect 18916 27770 18972 27772
rect 18996 27770 19052 27772
rect 19076 27770 19132 27772
rect 19156 27770 19212 27772
rect 19236 27770 19292 27772
rect 18916 27718 18918 27770
rect 18918 27718 18970 27770
rect 18970 27718 18972 27770
rect 18996 27718 19034 27770
rect 19034 27718 19046 27770
rect 19046 27718 19052 27770
rect 19076 27718 19098 27770
rect 19098 27718 19110 27770
rect 19110 27718 19132 27770
rect 19156 27718 19162 27770
rect 19162 27718 19174 27770
rect 19174 27718 19212 27770
rect 19236 27718 19238 27770
rect 19238 27718 19290 27770
rect 19290 27718 19292 27770
rect 18916 27716 18972 27718
rect 18996 27716 19052 27718
rect 19076 27716 19132 27718
rect 19156 27716 19212 27718
rect 19236 27716 19292 27718
rect 26916 27770 26972 27772
rect 26996 27770 27052 27772
rect 27076 27770 27132 27772
rect 27156 27770 27212 27772
rect 27236 27770 27292 27772
rect 26916 27718 26918 27770
rect 26918 27718 26970 27770
rect 26970 27718 26972 27770
rect 26996 27718 27034 27770
rect 27034 27718 27046 27770
rect 27046 27718 27052 27770
rect 27076 27718 27098 27770
rect 27098 27718 27110 27770
rect 27110 27718 27132 27770
rect 27156 27718 27162 27770
rect 27162 27718 27174 27770
rect 27174 27718 27212 27770
rect 27236 27718 27238 27770
rect 27238 27718 27290 27770
rect 27290 27718 27292 27770
rect 26916 27716 26972 27718
rect 26996 27716 27052 27718
rect 27076 27716 27132 27718
rect 27156 27716 27212 27718
rect 27236 27716 27292 27718
rect 846 27104 902 27160
rect 3656 27226 3712 27228
rect 3736 27226 3792 27228
rect 3816 27226 3872 27228
rect 3896 27226 3952 27228
rect 3976 27226 4032 27228
rect 3656 27174 3658 27226
rect 3658 27174 3710 27226
rect 3710 27174 3712 27226
rect 3736 27174 3774 27226
rect 3774 27174 3786 27226
rect 3786 27174 3792 27226
rect 3816 27174 3838 27226
rect 3838 27174 3850 27226
rect 3850 27174 3872 27226
rect 3896 27174 3902 27226
rect 3902 27174 3914 27226
rect 3914 27174 3952 27226
rect 3976 27174 3978 27226
rect 3978 27174 4030 27226
rect 4030 27174 4032 27226
rect 3656 27172 3712 27174
rect 3736 27172 3792 27174
rect 3816 27172 3872 27174
rect 3896 27172 3952 27174
rect 3976 27172 4032 27174
rect 28354 27532 28410 27568
rect 28354 27512 28356 27532
rect 28356 27512 28408 27532
rect 28408 27512 28410 27532
rect 11656 27226 11712 27228
rect 11736 27226 11792 27228
rect 11816 27226 11872 27228
rect 11896 27226 11952 27228
rect 11976 27226 12032 27228
rect 11656 27174 11658 27226
rect 11658 27174 11710 27226
rect 11710 27174 11712 27226
rect 11736 27174 11774 27226
rect 11774 27174 11786 27226
rect 11786 27174 11792 27226
rect 11816 27174 11838 27226
rect 11838 27174 11850 27226
rect 11850 27174 11872 27226
rect 11896 27174 11902 27226
rect 11902 27174 11914 27226
rect 11914 27174 11952 27226
rect 11976 27174 11978 27226
rect 11978 27174 12030 27226
rect 12030 27174 12032 27226
rect 11656 27172 11712 27174
rect 11736 27172 11792 27174
rect 11816 27172 11872 27174
rect 11896 27172 11952 27174
rect 11976 27172 12032 27174
rect 2916 26682 2972 26684
rect 2996 26682 3052 26684
rect 3076 26682 3132 26684
rect 3156 26682 3212 26684
rect 3236 26682 3292 26684
rect 2916 26630 2918 26682
rect 2918 26630 2970 26682
rect 2970 26630 2972 26682
rect 2996 26630 3034 26682
rect 3034 26630 3046 26682
rect 3046 26630 3052 26682
rect 3076 26630 3098 26682
rect 3098 26630 3110 26682
rect 3110 26630 3132 26682
rect 3156 26630 3162 26682
rect 3162 26630 3174 26682
rect 3174 26630 3212 26682
rect 3236 26630 3238 26682
rect 3238 26630 3290 26682
rect 3290 26630 3292 26682
rect 2916 26628 2972 26630
rect 2996 26628 3052 26630
rect 3076 26628 3132 26630
rect 3156 26628 3212 26630
rect 3236 26628 3292 26630
rect 10916 26682 10972 26684
rect 10996 26682 11052 26684
rect 11076 26682 11132 26684
rect 11156 26682 11212 26684
rect 11236 26682 11292 26684
rect 10916 26630 10918 26682
rect 10918 26630 10970 26682
rect 10970 26630 10972 26682
rect 10996 26630 11034 26682
rect 11034 26630 11046 26682
rect 11046 26630 11052 26682
rect 11076 26630 11098 26682
rect 11098 26630 11110 26682
rect 11110 26630 11132 26682
rect 11156 26630 11162 26682
rect 11162 26630 11174 26682
rect 11174 26630 11212 26682
rect 11236 26630 11238 26682
rect 11238 26630 11290 26682
rect 11290 26630 11292 26682
rect 10916 26628 10972 26630
rect 10996 26628 11052 26630
rect 11076 26628 11132 26630
rect 11156 26628 11212 26630
rect 11236 26628 11292 26630
rect 3656 26138 3712 26140
rect 3736 26138 3792 26140
rect 3816 26138 3872 26140
rect 3896 26138 3952 26140
rect 3976 26138 4032 26140
rect 3656 26086 3658 26138
rect 3658 26086 3710 26138
rect 3710 26086 3712 26138
rect 3736 26086 3774 26138
rect 3774 26086 3786 26138
rect 3786 26086 3792 26138
rect 3816 26086 3838 26138
rect 3838 26086 3850 26138
rect 3850 26086 3872 26138
rect 3896 26086 3902 26138
rect 3902 26086 3914 26138
rect 3914 26086 3952 26138
rect 3976 26086 3978 26138
rect 3978 26086 4030 26138
rect 4030 26086 4032 26138
rect 3656 26084 3712 26086
rect 3736 26084 3792 26086
rect 3816 26084 3872 26086
rect 3896 26084 3952 26086
rect 3976 26084 4032 26086
rect 846 26016 902 26072
rect 11656 26138 11712 26140
rect 11736 26138 11792 26140
rect 11816 26138 11872 26140
rect 11896 26138 11952 26140
rect 11976 26138 12032 26140
rect 11656 26086 11658 26138
rect 11658 26086 11710 26138
rect 11710 26086 11712 26138
rect 11736 26086 11774 26138
rect 11774 26086 11786 26138
rect 11786 26086 11792 26138
rect 11816 26086 11838 26138
rect 11838 26086 11850 26138
rect 11850 26086 11872 26138
rect 11896 26086 11902 26138
rect 11902 26086 11914 26138
rect 11914 26086 11952 26138
rect 11976 26086 11978 26138
rect 11978 26086 12030 26138
rect 12030 26086 12032 26138
rect 11656 26084 11712 26086
rect 11736 26084 11792 26086
rect 11816 26084 11872 26086
rect 11896 26084 11952 26086
rect 11976 26084 12032 26086
rect 2916 25594 2972 25596
rect 2996 25594 3052 25596
rect 3076 25594 3132 25596
rect 3156 25594 3212 25596
rect 3236 25594 3292 25596
rect 2916 25542 2918 25594
rect 2918 25542 2970 25594
rect 2970 25542 2972 25594
rect 2996 25542 3034 25594
rect 3034 25542 3046 25594
rect 3046 25542 3052 25594
rect 3076 25542 3098 25594
rect 3098 25542 3110 25594
rect 3110 25542 3132 25594
rect 3156 25542 3162 25594
rect 3162 25542 3174 25594
rect 3174 25542 3212 25594
rect 3236 25542 3238 25594
rect 3238 25542 3290 25594
rect 3290 25542 3292 25594
rect 2916 25540 2972 25542
rect 2996 25540 3052 25542
rect 3076 25540 3132 25542
rect 3156 25540 3212 25542
rect 3236 25540 3292 25542
rect 846 25472 902 25528
rect 3656 25050 3712 25052
rect 3736 25050 3792 25052
rect 3816 25050 3872 25052
rect 3896 25050 3952 25052
rect 3976 25050 4032 25052
rect 3656 24998 3658 25050
rect 3658 24998 3710 25050
rect 3710 24998 3712 25050
rect 3736 24998 3774 25050
rect 3774 24998 3786 25050
rect 3786 24998 3792 25050
rect 3816 24998 3838 25050
rect 3838 24998 3850 25050
rect 3850 24998 3872 25050
rect 3896 24998 3902 25050
rect 3902 24998 3914 25050
rect 3914 24998 3952 25050
rect 3976 24998 3978 25050
rect 3978 24998 4030 25050
rect 4030 24998 4032 25050
rect 3656 24996 3712 24998
rect 3736 24996 3792 24998
rect 3816 24996 3872 24998
rect 3896 24996 3952 24998
rect 3976 24996 4032 24998
rect 846 24656 902 24712
rect 2916 24506 2972 24508
rect 2996 24506 3052 24508
rect 3076 24506 3132 24508
rect 3156 24506 3212 24508
rect 3236 24506 3292 24508
rect 2916 24454 2918 24506
rect 2918 24454 2970 24506
rect 2970 24454 2972 24506
rect 2996 24454 3034 24506
rect 3034 24454 3046 24506
rect 3046 24454 3052 24506
rect 3076 24454 3098 24506
rect 3098 24454 3110 24506
rect 3110 24454 3132 24506
rect 3156 24454 3162 24506
rect 3162 24454 3174 24506
rect 3174 24454 3212 24506
rect 3236 24454 3238 24506
rect 3238 24454 3290 24506
rect 3290 24454 3292 24506
rect 2916 24452 2972 24454
rect 2996 24452 3052 24454
rect 3076 24452 3132 24454
rect 3156 24452 3212 24454
rect 3236 24452 3292 24454
rect 10916 25594 10972 25596
rect 10996 25594 11052 25596
rect 11076 25594 11132 25596
rect 11156 25594 11212 25596
rect 11236 25594 11292 25596
rect 10916 25542 10918 25594
rect 10918 25542 10970 25594
rect 10970 25542 10972 25594
rect 10996 25542 11034 25594
rect 11034 25542 11046 25594
rect 11046 25542 11052 25594
rect 11076 25542 11098 25594
rect 11098 25542 11110 25594
rect 11110 25542 11132 25594
rect 11156 25542 11162 25594
rect 11162 25542 11174 25594
rect 11174 25542 11212 25594
rect 11236 25542 11238 25594
rect 11238 25542 11290 25594
rect 11290 25542 11292 25594
rect 10916 25540 10972 25542
rect 10996 25540 11052 25542
rect 11076 25540 11132 25542
rect 11156 25540 11212 25542
rect 11236 25540 11292 25542
rect 11656 25050 11712 25052
rect 11736 25050 11792 25052
rect 11816 25050 11872 25052
rect 11896 25050 11952 25052
rect 11976 25050 12032 25052
rect 11656 24998 11658 25050
rect 11658 24998 11710 25050
rect 11710 24998 11712 25050
rect 11736 24998 11774 25050
rect 11774 24998 11786 25050
rect 11786 24998 11792 25050
rect 11816 24998 11838 25050
rect 11838 24998 11850 25050
rect 11850 24998 11872 25050
rect 11896 24998 11902 25050
rect 11902 24998 11914 25050
rect 11914 24998 11952 25050
rect 11976 24998 11978 25050
rect 11978 24998 12030 25050
rect 12030 24998 12032 25050
rect 11656 24996 11712 24998
rect 11736 24996 11792 24998
rect 11816 24996 11872 24998
rect 11896 24996 11952 24998
rect 11976 24996 12032 24998
rect 10916 24506 10972 24508
rect 10996 24506 11052 24508
rect 11076 24506 11132 24508
rect 11156 24506 11212 24508
rect 11236 24506 11292 24508
rect 10916 24454 10918 24506
rect 10918 24454 10970 24506
rect 10970 24454 10972 24506
rect 10996 24454 11034 24506
rect 11034 24454 11046 24506
rect 11046 24454 11052 24506
rect 11076 24454 11098 24506
rect 11098 24454 11110 24506
rect 11110 24454 11132 24506
rect 11156 24454 11162 24506
rect 11162 24454 11174 24506
rect 11174 24454 11212 24506
rect 11236 24454 11238 24506
rect 11238 24454 11290 24506
rect 11290 24454 11292 24506
rect 10916 24452 10972 24454
rect 10996 24452 11052 24454
rect 11076 24452 11132 24454
rect 11156 24452 11212 24454
rect 11236 24452 11292 24454
rect 846 23840 902 23896
rect 3656 23962 3712 23964
rect 3736 23962 3792 23964
rect 3816 23962 3872 23964
rect 3896 23962 3952 23964
rect 3976 23962 4032 23964
rect 3656 23910 3658 23962
rect 3658 23910 3710 23962
rect 3710 23910 3712 23962
rect 3736 23910 3774 23962
rect 3774 23910 3786 23962
rect 3786 23910 3792 23962
rect 3816 23910 3838 23962
rect 3838 23910 3850 23962
rect 3850 23910 3872 23962
rect 3896 23910 3902 23962
rect 3902 23910 3914 23962
rect 3914 23910 3952 23962
rect 3976 23910 3978 23962
rect 3978 23910 4030 23962
rect 4030 23910 4032 23962
rect 3656 23908 3712 23910
rect 3736 23908 3792 23910
rect 3816 23908 3872 23910
rect 3896 23908 3952 23910
rect 3976 23908 4032 23910
rect 2916 23418 2972 23420
rect 2996 23418 3052 23420
rect 3076 23418 3132 23420
rect 3156 23418 3212 23420
rect 3236 23418 3292 23420
rect 2916 23366 2918 23418
rect 2918 23366 2970 23418
rect 2970 23366 2972 23418
rect 2996 23366 3034 23418
rect 3034 23366 3046 23418
rect 3046 23366 3052 23418
rect 3076 23366 3098 23418
rect 3098 23366 3110 23418
rect 3110 23366 3132 23418
rect 3156 23366 3162 23418
rect 3162 23366 3174 23418
rect 3174 23366 3212 23418
rect 3236 23366 3238 23418
rect 3238 23366 3290 23418
rect 3290 23366 3292 23418
rect 2916 23364 2972 23366
rect 2996 23364 3052 23366
rect 3076 23364 3132 23366
rect 3156 23364 3212 23366
rect 3236 23364 3292 23366
rect 10916 23418 10972 23420
rect 10996 23418 11052 23420
rect 11076 23418 11132 23420
rect 11156 23418 11212 23420
rect 11236 23418 11292 23420
rect 10916 23366 10918 23418
rect 10918 23366 10970 23418
rect 10970 23366 10972 23418
rect 10996 23366 11034 23418
rect 11034 23366 11046 23418
rect 11046 23366 11052 23418
rect 11076 23366 11098 23418
rect 11098 23366 11110 23418
rect 11110 23366 11132 23418
rect 11156 23366 11162 23418
rect 11162 23366 11174 23418
rect 11174 23366 11212 23418
rect 11236 23366 11238 23418
rect 11238 23366 11290 23418
rect 11290 23366 11292 23418
rect 10916 23364 10972 23366
rect 10996 23364 11052 23366
rect 11076 23364 11132 23366
rect 11156 23364 11212 23366
rect 11236 23364 11292 23366
rect 846 23060 848 23080
rect 848 23060 900 23080
rect 900 23060 902 23080
rect 846 23024 902 23060
rect 3656 22874 3712 22876
rect 3736 22874 3792 22876
rect 3816 22874 3872 22876
rect 3896 22874 3952 22876
rect 3976 22874 4032 22876
rect 3656 22822 3658 22874
rect 3658 22822 3710 22874
rect 3710 22822 3712 22874
rect 3736 22822 3774 22874
rect 3774 22822 3786 22874
rect 3786 22822 3792 22874
rect 3816 22822 3838 22874
rect 3838 22822 3850 22874
rect 3850 22822 3872 22874
rect 3896 22822 3902 22874
rect 3902 22822 3914 22874
rect 3914 22822 3952 22874
rect 3976 22822 3978 22874
rect 3978 22822 4030 22874
rect 4030 22822 4032 22874
rect 3656 22820 3712 22822
rect 3736 22820 3792 22822
rect 3816 22820 3872 22822
rect 3896 22820 3952 22822
rect 3976 22820 4032 22822
rect 846 22208 902 22264
rect 2916 22330 2972 22332
rect 2996 22330 3052 22332
rect 3076 22330 3132 22332
rect 3156 22330 3212 22332
rect 3236 22330 3292 22332
rect 2916 22278 2918 22330
rect 2918 22278 2970 22330
rect 2970 22278 2972 22330
rect 2996 22278 3034 22330
rect 3034 22278 3046 22330
rect 3046 22278 3052 22330
rect 3076 22278 3098 22330
rect 3098 22278 3110 22330
rect 3110 22278 3132 22330
rect 3156 22278 3162 22330
rect 3162 22278 3174 22330
rect 3174 22278 3212 22330
rect 3236 22278 3238 22330
rect 3238 22278 3290 22330
rect 3290 22278 3292 22330
rect 2916 22276 2972 22278
rect 2996 22276 3052 22278
rect 3076 22276 3132 22278
rect 3156 22276 3212 22278
rect 3236 22276 3292 22278
rect 10916 22330 10972 22332
rect 10996 22330 11052 22332
rect 11076 22330 11132 22332
rect 11156 22330 11212 22332
rect 11236 22330 11292 22332
rect 10916 22278 10918 22330
rect 10918 22278 10970 22330
rect 10970 22278 10972 22330
rect 10996 22278 11034 22330
rect 11034 22278 11046 22330
rect 11046 22278 11052 22330
rect 11076 22278 11098 22330
rect 11098 22278 11110 22330
rect 11110 22278 11132 22330
rect 11156 22278 11162 22330
rect 11162 22278 11174 22330
rect 11174 22278 11212 22330
rect 11236 22278 11238 22330
rect 11238 22278 11290 22330
rect 11290 22278 11292 22330
rect 10916 22276 10972 22278
rect 10996 22276 11052 22278
rect 11076 22276 11132 22278
rect 11156 22276 11212 22278
rect 11236 22276 11292 22278
rect 11656 23962 11712 23964
rect 11736 23962 11792 23964
rect 11816 23962 11872 23964
rect 11896 23962 11952 23964
rect 11976 23962 12032 23964
rect 11656 23910 11658 23962
rect 11658 23910 11710 23962
rect 11710 23910 11712 23962
rect 11736 23910 11774 23962
rect 11774 23910 11786 23962
rect 11786 23910 11792 23962
rect 11816 23910 11838 23962
rect 11838 23910 11850 23962
rect 11850 23910 11872 23962
rect 11896 23910 11902 23962
rect 11902 23910 11914 23962
rect 11914 23910 11952 23962
rect 11976 23910 11978 23962
rect 11978 23910 12030 23962
rect 12030 23910 12032 23962
rect 11656 23908 11712 23910
rect 11736 23908 11792 23910
rect 11816 23908 11872 23910
rect 11896 23908 11952 23910
rect 11976 23908 12032 23910
rect 19656 27226 19712 27228
rect 19736 27226 19792 27228
rect 19816 27226 19872 27228
rect 19896 27226 19952 27228
rect 19976 27226 20032 27228
rect 19656 27174 19658 27226
rect 19658 27174 19710 27226
rect 19710 27174 19712 27226
rect 19736 27174 19774 27226
rect 19774 27174 19786 27226
rect 19786 27174 19792 27226
rect 19816 27174 19838 27226
rect 19838 27174 19850 27226
rect 19850 27174 19872 27226
rect 19896 27174 19902 27226
rect 19902 27174 19914 27226
rect 19914 27174 19952 27226
rect 19976 27174 19978 27226
rect 19978 27174 20030 27226
rect 20030 27174 20032 27226
rect 19656 27172 19712 27174
rect 19736 27172 19792 27174
rect 19816 27172 19872 27174
rect 19896 27172 19952 27174
rect 19976 27172 20032 27174
rect 3656 21786 3712 21788
rect 3736 21786 3792 21788
rect 3816 21786 3872 21788
rect 3896 21786 3952 21788
rect 3976 21786 4032 21788
rect 3656 21734 3658 21786
rect 3658 21734 3710 21786
rect 3710 21734 3712 21786
rect 3736 21734 3774 21786
rect 3774 21734 3786 21786
rect 3786 21734 3792 21786
rect 3816 21734 3838 21786
rect 3838 21734 3850 21786
rect 3850 21734 3872 21786
rect 3896 21734 3902 21786
rect 3902 21734 3914 21786
rect 3914 21734 3952 21786
rect 3976 21734 3978 21786
rect 3978 21734 4030 21786
rect 4030 21734 4032 21786
rect 3656 21732 3712 21734
rect 3736 21732 3792 21734
rect 3816 21732 3872 21734
rect 3896 21732 3952 21734
rect 3976 21732 4032 21734
rect 1398 21392 1454 21448
rect 2916 21242 2972 21244
rect 2996 21242 3052 21244
rect 3076 21242 3132 21244
rect 3156 21242 3212 21244
rect 3236 21242 3292 21244
rect 2916 21190 2918 21242
rect 2918 21190 2970 21242
rect 2970 21190 2972 21242
rect 2996 21190 3034 21242
rect 3034 21190 3046 21242
rect 3046 21190 3052 21242
rect 3076 21190 3098 21242
rect 3098 21190 3110 21242
rect 3110 21190 3132 21242
rect 3156 21190 3162 21242
rect 3162 21190 3174 21242
rect 3174 21190 3212 21242
rect 3236 21190 3238 21242
rect 3238 21190 3290 21242
rect 3290 21190 3292 21242
rect 2916 21188 2972 21190
rect 2996 21188 3052 21190
rect 3076 21188 3132 21190
rect 3156 21188 3212 21190
rect 3236 21188 3292 21190
rect 10916 21242 10972 21244
rect 10996 21242 11052 21244
rect 11076 21242 11132 21244
rect 11156 21242 11212 21244
rect 11236 21242 11292 21244
rect 10916 21190 10918 21242
rect 10918 21190 10970 21242
rect 10970 21190 10972 21242
rect 10996 21190 11034 21242
rect 11034 21190 11046 21242
rect 11046 21190 11052 21242
rect 11076 21190 11098 21242
rect 11098 21190 11110 21242
rect 11110 21190 11132 21242
rect 11156 21190 11162 21242
rect 11162 21190 11174 21242
rect 11174 21190 11212 21242
rect 11236 21190 11238 21242
rect 11238 21190 11290 21242
rect 11290 21190 11292 21242
rect 10916 21188 10972 21190
rect 10996 21188 11052 21190
rect 11076 21188 11132 21190
rect 11156 21188 11212 21190
rect 11236 21188 11292 21190
rect 3656 20698 3712 20700
rect 3736 20698 3792 20700
rect 3816 20698 3872 20700
rect 3896 20698 3952 20700
rect 3976 20698 4032 20700
rect 3656 20646 3658 20698
rect 3658 20646 3710 20698
rect 3710 20646 3712 20698
rect 3736 20646 3774 20698
rect 3774 20646 3786 20698
rect 3786 20646 3792 20698
rect 3816 20646 3838 20698
rect 3838 20646 3850 20698
rect 3850 20646 3872 20698
rect 3896 20646 3902 20698
rect 3902 20646 3914 20698
rect 3914 20646 3952 20698
rect 3976 20646 3978 20698
rect 3978 20646 4030 20698
rect 4030 20646 4032 20698
rect 3656 20644 3712 20646
rect 3736 20644 3792 20646
rect 3816 20644 3872 20646
rect 3896 20644 3952 20646
rect 3976 20644 4032 20646
rect 1398 20576 1454 20632
rect 2916 20154 2972 20156
rect 2996 20154 3052 20156
rect 3076 20154 3132 20156
rect 3156 20154 3212 20156
rect 3236 20154 3292 20156
rect 2916 20102 2918 20154
rect 2918 20102 2970 20154
rect 2970 20102 2972 20154
rect 2996 20102 3034 20154
rect 3034 20102 3046 20154
rect 3046 20102 3052 20154
rect 3076 20102 3098 20154
rect 3098 20102 3110 20154
rect 3110 20102 3132 20154
rect 3156 20102 3162 20154
rect 3162 20102 3174 20154
rect 3174 20102 3212 20154
rect 3236 20102 3238 20154
rect 3238 20102 3290 20154
rect 3290 20102 3292 20154
rect 2916 20100 2972 20102
rect 2996 20100 3052 20102
rect 3076 20100 3132 20102
rect 3156 20100 3212 20102
rect 3236 20100 3292 20102
rect 10916 20154 10972 20156
rect 10996 20154 11052 20156
rect 11076 20154 11132 20156
rect 11156 20154 11212 20156
rect 11236 20154 11292 20156
rect 10916 20102 10918 20154
rect 10918 20102 10970 20154
rect 10970 20102 10972 20154
rect 10996 20102 11034 20154
rect 11034 20102 11046 20154
rect 11046 20102 11052 20154
rect 11076 20102 11098 20154
rect 11098 20102 11110 20154
rect 11110 20102 11132 20154
rect 11156 20102 11162 20154
rect 11162 20102 11174 20154
rect 11174 20102 11212 20154
rect 11236 20102 11238 20154
rect 11238 20102 11290 20154
rect 11290 20102 11292 20154
rect 10916 20100 10972 20102
rect 10996 20100 11052 20102
rect 11076 20100 11132 20102
rect 11156 20100 11212 20102
rect 11236 20100 11292 20102
rect 1398 19796 1400 19816
rect 1400 19796 1452 19816
rect 1452 19796 1454 19816
rect 1398 19760 1454 19796
rect 3656 19610 3712 19612
rect 3736 19610 3792 19612
rect 3816 19610 3872 19612
rect 3896 19610 3952 19612
rect 3976 19610 4032 19612
rect 3656 19558 3658 19610
rect 3658 19558 3710 19610
rect 3710 19558 3712 19610
rect 3736 19558 3774 19610
rect 3774 19558 3786 19610
rect 3786 19558 3792 19610
rect 3816 19558 3838 19610
rect 3838 19558 3850 19610
rect 3850 19558 3872 19610
rect 3896 19558 3902 19610
rect 3902 19558 3914 19610
rect 3914 19558 3952 19610
rect 3976 19558 3978 19610
rect 3978 19558 4030 19610
rect 4030 19558 4032 19610
rect 3656 19556 3712 19558
rect 3736 19556 3792 19558
rect 3816 19556 3872 19558
rect 3896 19556 3952 19558
rect 3976 19556 4032 19558
rect 2916 19066 2972 19068
rect 2996 19066 3052 19068
rect 3076 19066 3132 19068
rect 3156 19066 3212 19068
rect 3236 19066 3292 19068
rect 2916 19014 2918 19066
rect 2918 19014 2970 19066
rect 2970 19014 2972 19066
rect 2996 19014 3034 19066
rect 3034 19014 3046 19066
rect 3046 19014 3052 19066
rect 3076 19014 3098 19066
rect 3098 19014 3110 19066
rect 3110 19014 3132 19066
rect 3156 19014 3162 19066
rect 3162 19014 3174 19066
rect 3174 19014 3212 19066
rect 3236 19014 3238 19066
rect 3238 19014 3290 19066
rect 3290 19014 3292 19066
rect 2916 19012 2972 19014
rect 2996 19012 3052 19014
rect 3076 19012 3132 19014
rect 3156 19012 3212 19014
rect 3236 19012 3292 19014
rect 10916 19066 10972 19068
rect 10996 19066 11052 19068
rect 11076 19066 11132 19068
rect 11156 19066 11212 19068
rect 11236 19066 11292 19068
rect 10916 19014 10918 19066
rect 10918 19014 10970 19066
rect 10970 19014 10972 19066
rect 10996 19014 11034 19066
rect 11034 19014 11046 19066
rect 11046 19014 11052 19066
rect 11076 19014 11098 19066
rect 11098 19014 11110 19066
rect 11110 19014 11132 19066
rect 11156 19014 11162 19066
rect 11162 19014 11174 19066
rect 11174 19014 11212 19066
rect 11236 19014 11238 19066
rect 11238 19014 11290 19066
rect 11290 19014 11292 19066
rect 10916 19012 10972 19014
rect 10996 19012 11052 19014
rect 11076 19012 11132 19014
rect 11156 19012 11212 19014
rect 11236 19012 11292 19014
rect 846 18944 902 19000
rect 3656 18522 3712 18524
rect 3736 18522 3792 18524
rect 3816 18522 3872 18524
rect 3896 18522 3952 18524
rect 3976 18522 4032 18524
rect 3656 18470 3658 18522
rect 3658 18470 3710 18522
rect 3710 18470 3712 18522
rect 3736 18470 3774 18522
rect 3774 18470 3786 18522
rect 3786 18470 3792 18522
rect 3816 18470 3838 18522
rect 3838 18470 3850 18522
rect 3850 18470 3872 18522
rect 3896 18470 3902 18522
rect 3902 18470 3914 18522
rect 3914 18470 3952 18522
rect 3976 18470 3978 18522
rect 3978 18470 4030 18522
rect 4030 18470 4032 18522
rect 3656 18468 3712 18470
rect 3736 18468 3792 18470
rect 3816 18468 3872 18470
rect 3896 18468 3952 18470
rect 3976 18468 4032 18470
rect 1398 17992 1454 18048
rect 2916 17978 2972 17980
rect 2996 17978 3052 17980
rect 3076 17978 3132 17980
rect 3156 17978 3212 17980
rect 3236 17978 3292 17980
rect 2916 17926 2918 17978
rect 2918 17926 2970 17978
rect 2970 17926 2972 17978
rect 2996 17926 3034 17978
rect 3034 17926 3046 17978
rect 3046 17926 3052 17978
rect 3076 17926 3098 17978
rect 3098 17926 3110 17978
rect 3110 17926 3132 17978
rect 3156 17926 3162 17978
rect 3162 17926 3174 17978
rect 3174 17926 3212 17978
rect 3236 17926 3238 17978
rect 3238 17926 3290 17978
rect 3290 17926 3292 17978
rect 2916 17924 2972 17926
rect 2996 17924 3052 17926
rect 3076 17924 3132 17926
rect 3156 17924 3212 17926
rect 3236 17924 3292 17926
rect 10916 17978 10972 17980
rect 10996 17978 11052 17980
rect 11076 17978 11132 17980
rect 11156 17978 11212 17980
rect 11236 17978 11292 17980
rect 10916 17926 10918 17978
rect 10918 17926 10970 17978
rect 10970 17926 10972 17978
rect 10996 17926 11034 17978
rect 11034 17926 11046 17978
rect 11046 17926 11052 17978
rect 11076 17926 11098 17978
rect 11098 17926 11110 17978
rect 11110 17926 11132 17978
rect 11156 17926 11162 17978
rect 11162 17926 11174 17978
rect 11174 17926 11212 17978
rect 11236 17926 11238 17978
rect 11238 17926 11290 17978
rect 11290 17926 11292 17978
rect 10916 17924 10972 17926
rect 10996 17924 11052 17926
rect 11076 17924 11132 17926
rect 11156 17924 11212 17926
rect 11236 17924 11292 17926
rect 3656 17434 3712 17436
rect 3736 17434 3792 17436
rect 3816 17434 3872 17436
rect 3896 17434 3952 17436
rect 3976 17434 4032 17436
rect 3656 17382 3658 17434
rect 3658 17382 3710 17434
rect 3710 17382 3712 17434
rect 3736 17382 3774 17434
rect 3774 17382 3786 17434
rect 3786 17382 3792 17434
rect 3816 17382 3838 17434
rect 3838 17382 3850 17434
rect 3850 17382 3872 17434
rect 3896 17382 3902 17434
rect 3902 17382 3914 17434
rect 3914 17382 3952 17434
rect 3976 17382 3978 17434
rect 3978 17382 4030 17434
rect 4030 17382 4032 17434
rect 3656 17380 3712 17382
rect 3736 17380 3792 17382
rect 3816 17380 3872 17382
rect 3896 17380 3952 17382
rect 3976 17380 4032 17382
rect 1398 17312 1454 17368
rect 2916 16890 2972 16892
rect 2996 16890 3052 16892
rect 3076 16890 3132 16892
rect 3156 16890 3212 16892
rect 3236 16890 3292 16892
rect 2916 16838 2918 16890
rect 2918 16838 2970 16890
rect 2970 16838 2972 16890
rect 2996 16838 3034 16890
rect 3034 16838 3046 16890
rect 3046 16838 3052 16890
rect 3076 16838 3098 16890
rect 3098 16838 3110 16890
rect 3110 16838 3132 16890
rect 3156 16838 3162 16890
rect 3162 16838 3174 16890
rect 3174 16838 3212 16890
rect 3236 16838 3238 16890
rect 3238 16838 3290 16890
rect 3290 16838 3292 16890
rect 2916 16836 2972 16838
rect 2996 16836 3052 16838
rect 3076 16836 3132 16838
rect 3156 16836 3212 16838
rect 3236 16836 3292 16838
rect 10916 16890 10972 16892
rect 10996 16890 11052 16892
rect 11076 16890 11132 16892
rect 11156 16890 11212 16892
rect 11236 16890 11292 16892
rect 10916 16838 10918 16890
rect 10918 16838 10970 16890
rect 10970 16838 10972 16890
rect 10996 16838 11034 16890
rect 11034 16838 11046 16890
rect 11046 16838 11052 16890
rect 11076 16838 11098 16890
rect 11098 16838 11110 16890
rect 11110 16838 11132 16890
rect 11156 16838 11162 16890
rect 11162 16838 11174 16890
rect 11174 16838 11212 16890
rect 11236 16838 11238 16890
rect 11238 16838 11290 16890
rect 11290 16838 11292 16890
rect 10916 16836 10972 16838
rect 10996 16836 11052 16838
rect 11076 16836 11132 16838
rect 11156 16836 11212 16838
rect 11236 16836 11292 16838
rect 1398 16532 1400 16552
rect 1400 16532 1452 16552
rect 1452 16532 1454 16552
rect 1398 16496 1454 16532
rect 3656 16346 3712 16348
rect 3736 16346 3792 16348
rect 3816 16346 3872 16348
rect 3896 16346 3952 16348
rect 3976 16346 4032 16348
rect 3656 16294 3658 16346
rect 3658 16294 3710 16346
rect 3710 16294 3712 16346
rect 3736 16294 3774 16346
rect 3774 16294 3786 16346
rect 3786 16294 3792 16346
rect 3816 16294 3838 16346
rect 3838 16294 3850 16346
rect 3850 16294 3872 16346
rect 3896 16294 3902 16346
rect 3902 16294 3914 16346
rect 3914 16294 3952 16346
rect 3976 16294 3978 16346
rect 3978 16294 4030 16346
rect 4030 16294 4032 16346
rect 3656 16292 3712 16294
rect 3736 16292 3792 16294
rect 3816 16292 3872 16294
rect 3896 16292 3952 16294
rect 3976 16292 4032 16294
rect 2916 15802 2972 15804
rect 2996 15802 3052 15804
rect 3076 15802 3132 15804
rect 3156 15802 3212 15804
rect 3236 15802 3292 15804
rect 2916 15750 2918 15802
rect 2918 15750 2970 15802
rect 2970 15750 2972 15802
rect 2996 15750 3034 15802
rect 3034 15750 3046 15802
rect 3046 15750 3052 15802
rect 3076 15750 3098 15802
rect 3098 15750 3110 15802
rect 3110 15750 3132 15802
rect 3156 15750 3162 15802
rect 3162 15750 3174 15802
rect 3174 15750 3212 15802
rect 3236 15750 3238 15802
rect 3238 15750 3290 15802
rect 3290 15750 3292 15802
rect 2916 15748 2972 15750
rect 2996 15748 3052 15750
rect 3076 15748 3132 15750
rect 3156 15748 3212 15750
rect 3236 15748 3292 15750
rect 1398 15680 1454 15736
rect 3656 15258 3712 15260
rect 3736 15258 3792 15260
rect 3816 15258 3872 15260
rect 3896 15258 3952 15260
rect 3976 15258 4032 15260
rect 3656 15206 3658 15258
rect 3658 15206 3710 15258
rect 3710 15206 3712 15258
rect 3736 15206 3774 15258
rect 3774 15206 3786 15258
rect 3786 15206 3792 15258
rect 3816 15206 3838 15258
rect 3838 15206 3850 15258
rect 3850 15206 3872 15258
rect 3896 15206 3902 15258
rect 3902 15206 3914 15258
rect 3914 15206 3952 15258
rect 3976 15206 3978 15258
rect 3978 15206 4030 15258
rect 4030 15206 4032 15258
rect 3656 15204 3712 15206
rect 3736 15204 3792 15206
rect 3816 15204 3872 15206
rect 3896 15204 3952 15206
rect 3976 15204 4032 15206
rect 10916 15802 10972 15804
rect 10996 15802 11052 15804
rect 11076 15802 11132 15804
rect 11156 15802 11212 15804
rect 11236 15802 11292 15804
rect 10916 15750 10918 15802
rect 10918 15750 10970 15802
rect 10970 15750 10972 15802
rect 10996 15750 11034 15802
rect 11034 15750 11046 15802
rect 11046 15750 11052 15802
rect 11076 15750 11098 15802
rect 11098 15750 11110 15802
rect 11110 15750 11132 15802
rect 11156 15750 11162 15802
rect 11162 15750 11174 15802
rect 11174 15750 11212 15802
rect 11236 15750 11238 15802
rect 11238 15750 11290 15802
rect 11290 15750 11292 15802
rect 10916 15748 10972 15750
rect 10996 15748 11052 15750
rect 11076 15748 11132 15750
rect 11156 15748 11212 15750
rect 11236 15748 11292 15750
rect 11656 22874 11712 22876
rect 11736 22874 11792 22876
rect 11816 22874 11872 22876
rect 11896 22874 11952 22876
rect 11976 22874 12032 22876
rect 11656 22822 11658 22874
rect 11658 22822 11710 22874
rect 11710 22822 11712 22874
rect 11736 22822 11774 22874
rect 11774 22822 11786 22874
rect 11786 22822 11792 22874
rect 11816 22822 11838 22874
rect 11838 22822 11850 22874
rect 11850 22822 11872 22874
rect 11896 22822 11902 22874
rect 11902 22822 11914 22874
rect 11914 22822 11952 22874
rect 11976 22822 11978 22874
rect 11978 22822 12030 22874
rect 12030 22822 12032 22874
rect 11656 22820 11712 22822
rect 11736 22820 11792 22822
rect 11816 22820 11872 22822
rect 11896 22820 11952 22822
rect 11976 22820 12032 22822
rect 11656 21786 11712 21788
rect 11736 21786 11792 21788
rect 11816 21786 11872 21788
rect 11896 21786 11952 21788
rect 11976 21786 12032 21788
rect 11656 21734 11658 21786
rect 11658 21734 11710 21786
rect 11710 21734 11712 21786
rect 11736 21734 11774 21786
rect 11774 21734 11786 21786
rect 11786 21734 11792 21786
rect 11816 21734 11838 21786
rect 11838 21734 11850 21786
rect 11850 21734 11872 21786
rect 11896 21734 11902 21786
rect 11902 21734 11914 21786
rect 11914 21734 11952 21786
rect 11976 21734 11978 21786
rect 11978 21734 12030 21786
rect 12030 21734 12032 21786
rect 11656 21732 11712 21734
rect 11736 21732 11792 21734
rect 11816 21732 11872 21734
rect 11896 21732 11952 21734
rect 11976 21732 12032 21734
rect 27656 27226 27712 27228
rect 27736 27226 27792 27228
rect 27816 27226 27872 27228
rect 27896 27226 27952 27228
rect 27976 27226 28032 27228
rect 27656 27174 27658 27226
rect 27658 27174 27710 27226
rect 27710 27174 27712 27226
rect 27736 27174 27774 27226
rect 27774 27174 27786 27226
rect 27786 27174 27792 27226
rect 27816 27174 27838 27226
rect 27838 27174 27850 27226
rect 27850 27174 27872 27226
rect 27896 27174 27902 27226
rect 27902 27174 27914 27226
rect 27914 27174 27952 27226
rect 27976 27174 27978 27226
rect 27978 27174 28030 27226
rect 28030 27174 28032 27226
rect 27656 27172 27712 27174
rect 27736 27172 27792 27174
rect 27816 27172 27872 27174
rect 27896 27172 27952 27174
rect 27976 27172 28032 27174
rect 18916 26682 18972 26684
rect 18996 26682 19052 26684
rect 19076 26682 19132 26684
rect 19156 26682 19212 26684
rect 19236 26682 19292 26684
rect 18916 26630 18918 26682
rect 18918 26630 18970 26682
rect 18970 26630 18972 26682
rect 18996 26630 19034 26682
rect 19034 26630 19046 26682
rect 19046 26630 19052 26682
rect 19076 26630 19098 26682
rect 19098 26630 19110 26682
rect 19110 26630 19132 26682
rect 19156 26630 19162 26682
rect 19162 26630 19174 26682
rect 19174 26630 19212 26682
rect 19236 26630 19238 26682
rect 19238 26630 19290 26682
rect 19290 26630 19292 26682
rect 18916 26628 18972 26630
rect 18996 26628 19052 26630
rect 19076 26628 19132 26630
rect 19156 26628 19212 26630
rect 19236 26628 19292 26630
rect 28354 26696 28410 26752
rect 26916 26682 26972 26684
rect 26996 26682 27052 26684
rect 27076 26682 27132 26684
rect 27156 26682 27212 26684
rect 27236 26682 27292 26684
rect 26916 26630 26918 26682
rect 26918 26630 26970 26682
rect 26970 26630 26972 26682
rect 26996 26630 27034 26682
rect 27034 26630 27046 26682
rect 27046 26630 27052 26682
rect 27076 26630 27098 26682
rect 27098 26630 27110 26682
rect 27110 26630 27132 26682
rect 27156 26630 27162 26682
rect 27162 26630 27174 26682
rect 27174 26630 27212 26682
rect 27236 26630 27238 26682
rect 27238 26630 27290 26682
rect 27290 26630 27292 26682
rect 26916 26628 26972 26630
rect 26996 26628 27052 26630
rect 27076 26628 27132 26630
rect 27156 26628 27212 26630
rect 27236 26628 27292 26630
rect 19656 26138 19712 26140
rect 19736 26138 19792 26140
rect 19816 26138 19872 26140
rect 19896 26138 19952 26140
rect 19976 26138 20032 26140
rect 19656 26086 19658 26138
rect 19658 26086 19710 26138
rect 19710 26086 19712 26138
rect 19736 26086 19774 26138
rect 19774 26086 19786 26138
rect 19786 26086 19792 26138
rect 19816 26086 19838 26138
rect 19838 26086 19850 26138
rect 19850 26086 19872 26138
rect 19896 26086 19902 26138
rect 19902 26086 19914 26138
rect 19914 26086 19952 26138
rect 19976 26086 19978 26138
rect 19978 26086 20030 26138
rect 20030 26086 20032 26138
rect 19656 26084 19712 26086
rect 19736 26084 19792 26086
rect 19816 26084 19872 26086
rect 19896 26084 19952 26086
rect 19976 26084 20032 26086
rect 27656 26138 27712 26140
rect 27736 26138 27792 26140
rect 27816 26138 27872 26140
rect 27896 26138 27952 26140
rect 27976 26138 28032 26140
rect 27656 26086 27658 26138
rect 27658 26086 27710 26138
rect 27710 26086 27712 26138
rect 27736 26086 27774 26138
rect 27774 26086 27786 26138
rect 27786 26086 27792 26138
rect 27816 26086 27838 26138
rect 27838 26086 27850 26138
rect 27850 26086 27872 26138
rect 27896 26086 27902 26138
rect 27902 26086 27914 26138
rect 27914 26086 27952 26138
rect 27976 26086 27978 26138
rect 27978 26086 28030 26138
rect 28030 26086 28032 26138
rect 27656 26084 27712 26086
rect 27736 26084 27792 26086
rect 27816 26084 27872 26086
rect 27896 26084 27952 26086
rect 27976 26084 28032 26086
rect 28354 25880 28410 25936
rect 18916 25594 18972 25596
rect 18996 25594 19052 25596
rect 19076 25594 19132 25596
rect 19156 25594 19212 25596
rect 19236 25594 19292 25596
rect 18916 25542 18918 25594
rect 18918 25542 18970 25594
rect 18970 25542 18972 25594
rect 18996 25542 19034 25594
rect 19034 25542 19046 25594
rect 19046 25542 19052 25594
rect 19076 25542 19098 25594
rect 19098 25542 19110 25594
rect 19110 25542 19132 25594
rect 19156 25542 19162 25594
rect 19162 25542 19174 25594
rect 19174 25542 19212 25594
rect 19236 25542 19238 25594
rect 19238 25542 19290 25594
rect 19290 25542 19292 25594
rect 18916 25540 18972 25542
rect 18996 25540 19052 25542
rect 19076 25540 19132 25542
rect 19156 25540 19212 25542
rect 19236 25540 19292 25542
rect 26916 25594 26972 25596
rect 26996 25594 27052 25596
rect 27076 25594 27132 25596
rect 27156 25594 27212 25596
rect 27236 25594 27292 25596
rect 26916 25542 26918 25594
rect 26918 25542 26970 25594
rect 26970 25542 26972 25594
rect 26996 25542 27034 25594
rect 27034 25542 27046 25594
rect 27046 25542 27052 25594
rect 27076 25542 27098 25594
rect 27098 25542 27110 25594
rect 27110 25542 27132 25594
rect 27156 25542 27162 25594
rect 27162 25542 27174 25594
rect 27174 25542 27212 25594
rect 27236 25542 27238 25594
rect 27238 25542 27290 25594
rect 27290 25542 27292 25594
rect 26916 25540 26972 25542
rect 26996 25540 27052 25542
rect 27076 25540 27132 25542
rect 27156 25540 27212 25542
rect 27236 25540 27292 25542
rect 28354 25064 28410 25120
rect 19656 25050 19712 25052
rect 19736 25050 19792 25052
rect 19816 25050 19872 25052
rect 19896 25050 19952 25052
rect 19976 25050 20032 25052
rect 19656 24998 19658 25050
rect 19658 24998 19710 25050
rect 19710 24998 19712 25050
rect 19736 24998 19774 25050
rect 19774 24998 19786 25050
rect 19786 24998 19792 25050
rect 19816 24998 19838 25050
rect 19838 24998 19850 25050
rect 19850 24998 19872 25050
rect 19896 24998 19902 25050
rect 19902 24998 19914 25050
rect 19914 24998 19952 25050
rect 19976 24998 19978 25050
rect 19978 24998 20030 25050
rect 20030 24998 20032 25050
rect 19656 24996 19712 24998
rect 19736 24996 19792 24998
rect 19816 24996 19872 24998
rect 19896 24996 19952 24998
rect 19976 24996 20032 24998
rect 27656 25050 27712 25052
rect 27736 25050 27792 25052
rect 27816 25050 27872 25052
rect 27896 25050 27952 25052
rect 27976 25050 28032 25052
rect 27656 24998 27658 25050
rect 27658 24998 27710 25050
rect 27710 24998 27712 25050
rect 27736 24998 27774 25050
rect 27774 24998 27786 25050
rect 27786 24998 27792 25050
rect 27816 24998 27838 25050
rect 27838 24998 27850 25050
rect 27850 24998 27872 25050
rect 27896 24998 27902 25050
rect 27902 24998 27914 25050
rect 27914 24998 27952 25050
rect 27976 24998 27978 25050
rect 27978 24998 28030 25050
rect 28030 24998 28032 25050
rect 27656 24996 27712 24998
rect 27736 24996 27792 24998
rect 27816 24996 27872 24998
rect 27896 24996 27952 24998
rect 27976 24996 28032 24998
rect 18916 24506 18972 24508
rect 18996 24506 19052 24508
rect 19076 24506 19132 24508
rect 19156 24506 19212 24508
rect 19236 24506 19292 24508
rect 18916 24454 18918 24506
rect 18918 24454 18970 24506
rect 18970 24454 18972 24506
rect 18996 24454 19034 24506
rect 19034 24454 19046 24506
rect 19046 24454 19052 24506
rect 19076 24454 19098 24506
rect 19098 24454 19110 24506
rect 19110 24454 19132 24506
rect 19156 24454 19162 24506
rect 19162 24454 19174 24506
rect 19174 24454 19212 24506
rect 19236 24454 19238 24506
rect 19238 24454 19290 24506
rect 19290 24454 19292 24506
rect 18916 24452 18972 24454
rect 18996 24452 19052 24454
rect 19076 24452 19132 24454
rect 19156 24452 19212 24454
rect 19236 24452 19292 24454
rect 26916 24506 26972 24508
rect 26996 24506 27052 24508
rect 27076 24506 27132 24508
rect 27156 24506 27212 24508
rect 27236 24506 27292 24508
rect 26916 24454 26918 24506
rect 26918 24454 26970 24506
rect 26970 24454 26972 24506
rect 26996 24454 27034 24506
rect 27034 24454 27046 24506
rect 27046 24454 27052 24506
rect 27076 24454 27098 24506
rect 27098 24454 27110 24506
rect 27110 24454 27132 24506
rect 27156 24454 27162 24506
rect 27162 24454 27174 24506
rect 27174 24454 27212 24506
rect 27236 24454 27238 24506
rect 27238 24454 27290 24506
rect 27290 24454 27292 24506
rect 26916 24452 26972 24454
rect 26996 24452 27052 24454
rect 27076 24452 27132 24454
rect 27156 24452 27212 24454
rect 27236 24452 27292 24454
rect 28354 24248 28410 24304
rect 11656 20698 11712 20700
rect 11736 20698 11792 20700
rect 11816 20698 11872 20700
rect 11896 20698 11952 20700
rect 11976 20698 12032 20700
rect 11656 20646 11658 20698
rect 11658 20646 11710 20698
rect 11710 20646 11712 20698
rect 11736 20646 11774 20698
rect 11774 20646 11786 20698
rect 11786 20646 11792 20698
rect 11816 20646 11838 20698
rect 11838 20646 11850 20698
rect 11850 20646 11872 20698
rect 11896 20646 11902 20698
rect 11902 20646 11914 20698
rect 11914 20646 11952 20698
rect 11976 20646 11978 20698
rect 11978 20646 12030 20698
rect 12030 20646 12032 20698
rect 11656 20644 11712 20646
rect 11736 20644 11792 20646
rect 11816 20644 11872 20646
rect 11896 20644 11952 20646
rect 11976 20644 12032 20646
rect 11656 19610 11712 19612
rect 11736 19610 11792 19612
rect 11816 19610 11872 19612
rect 11896 19610 11952 19612
rect 11976 19610 12032 19612
rect 11656 19558 11658 19610
rect 11658 19558 11710 19610
rect 11710 19558 11712 19610
rect 11736 19558 11774 19610
rect 11774 19558 11786 19610
rect 11786 19558 11792 19610
rect 11816 19558 11838 19610
rect 11838 19558 11850 19610
rect 11850 19558 11872 19610
rect 11896 19558 11902 19610
rect 11902 19558 11914 19610
rect 11914 19558 11952 19610
rect 11976 19558 11978 19610
rect 11978 19558 12030 19610
rect 12030 19558 12032 19610
rect 11656 19556 11712 19558
rect 11736 19556 11792 19558
rect 11816 19556 11872 19558
rect 11896 19556 11952 19558
rect 11976 19556 12032 19558
rect 19656 23962 19712 23964
rect 19736 23962 19792 23964
rect 19816 23962 19872 23964
rect 19896 23962 19952 23964
rect 19976 23962 20032 23964
rect 19656 23910 19658 23962
rect 19658 23910 19710 23962
rect 19710 23910 19712 23962
rect 19736 23910 19774 23962
rect 19774 23910 19786 23962
rect 19786 23910 19792 23962
rect 19816 23910 19838 23962
rect 19838 23910 19850 23962
rect 19850 23910 19872 23962
rect 19896 23910 19902 23962
rect 19902 23910 19914 23962
rect 19914 23910 19952 23962
rect 19976 23910 19978 23962
rect 19978 23910 20030 23962
rect 20030 23910 20032 23962
rect 19656 23908 19712 23910
rect 19736 23908 19792 23910
rect 19816 23908 19872 23910
rect 19896 23908 19952 23910
rect 19976 23908 20032 23910
rect 27656 23962 27712 23964
rect 27736 23962 27792 23964
rect 27816 23962 27872 23964
rect 27896 23962 27952 23964
rect 27976 23962 28032 23964
rect 27656 23910 27658 23962
rect 27658 23910 27710 23962
rect 27710 23910 27712 23962
rect 27736 23910 27774 23962
rect 27774 23910 27786 23962
rect 27786 23910 27792 23962
rect 27816 23910 27838 23962
rect 27838 23910 27850 23962
rect 27850 23910 27872 23962
rect 27896 23910 27902 23962
rect 27902 23910 27914 23962
rect 27914 23910 27952 23962
rect 27976 23910 27978 23962
rect 27978 23910 28030 23962
rect 28030 23910 28032 23962
rect 27656 23908 27712 23910
rect 27736 23908 27792 23910
rect 27816 23908 27872 23910
rect 27896 23908 27952 23910
rect 27976 23908 28032 23910
rect 28354 23432 28410 23488
rect 18916 23418 18972 23420
rect 18996 23418 19052 23420
rect 19076 23418 19132 23420
rect 19156 23418 19212 23420
rect 19236 23418 19292 23420
rect 18916 23366 18918 23418
rect 18918 23366 18970 23418
rect 18970 23366 18972 23418
rect 18996 23366 19034 23418
rect 19034 23366 19046 23418
rect 19046 23366 19052 23418
rect 19076 23366 19098 23418
rect 19098 23366 19110 23418
rect 19110 23366 19132 23418
rect 19156 23366 19162 23418
rect 19162 23366 19174 23418
rect 19174 23366 19212 23418
rect 19236 23366 19238 23418
rect 19238 23366 19290 23418
rect 19290 23366 19292 23418
rect 18916 23364 18972 23366
rect 18996 23364 19052 23366
rect 19076 23364 19132 23366
rect 19156 23364 19212 23366
rect 19236 23364 19292 23366
rect 26916 23418 26972 23420
rect 26996 23418 27052 23420
rect 27076 23418 27132 23420
rect 27156 23418 27212 23420
rect 27236 23418 27292 23420
rect 26916 23366 26918 23418
rect 26918 23366 26970 23418
rect 26970 23366 26972 23418
rect 26996 23366 27034 23418
rect 27034 23366 27046 23418
rect 27046 23366 27052 23418
rect 27076 23366 27098 23418
rect 27098 23366 27110 23418
rect 27110 23366 27132 23418
rect 27156 23366 27162 23418
rect 27162 23366 27174 23418
rect 27174 23366 27212 23418
rect 27236 23366 27238 23418
rect 27238 23366 27290 23418
rect 27290 23366 27292 23418
rect 26916 23364 26972 23366
rect 26996 23364 27052 23366
rect 27076 23364 27132 23366
rect 27156 23364 27212 23366
rect 27236 23364 27292 23366
rect 19656 22874 19712 22876
rect 19736 22874 19792 22876
rect 19816 22874 19872 22876
rect 19896 22874 19952 22876
rect 19976 22874 20032 22876
rect 19656 22822 19658 22874
rect 19658 22822 19710 22874
rect 19710 22822 19712 22874
rect 19736 22822 19774 22874
rect 19774 22822 19786 22874
rect 19786 22822 19792 22874
rect 19816 22822 19838 22874
rect 19838 22822 19850 22874
rect 19850 22822 19872 22874
rect 19896 22822 19902 22874
rect 19902 22822 19914 22874
rect 19914 22822 19952 22874
rect 19976 22822 19978 22874
rect 19978 22822 20030 22874
rect 20030 22822 20032 22874
rect 19656 22820 19712 22822
rect 19736 22820 19792 22822
rect 19816 22820 19872 22822
rect 19896 22820 19952 22822
rect 19976 22820 20032 22822
rect 27656 22874 27712 22876
rect 27736 22874 27792 22876
rect 27816 22874 27872 22876
rect 27896 22874 27952 22876
rect 27976 22874 28032 22876
rect 27656 22822 27658 22874
rect 27658 22822 27710 22874
rect 27710 22822 27712 22874
rect 27736 22822 27774 22874
rect 27774 22822 27786 22874
rect 27786 22822 27792 22874
rect 27816 22822 27838 22874
rect 27838 22822 27850 22874
rect 27850 22822 27872 22874
rect 27896 22822 27902 22874
rect 27902 22822 27914 22874
rect 27914 22822 27952 22874
rect 27976 22822 27978 22874
rect 27978 22822 28030 22874
rect 28030 22822 28032 22874
rect 27656 22820 27712 22822
rect 27736 22820 27792 22822
rect 27816 22820 27872 22822
rect 27896 22820 27952 22822
rect 27976 22820 28032 22822
rect 28354 22616 28410 22672
rect 18916 22330 18972 22332
rect 18996 22330 19052 22332
rect 19076 22330 19132 22332
rect 19156 22330 19212 22332
rect 19236 22330 19292 22332
rect 18916 22278 18918 22330
rect 18918 22278 18970 22330
rect 18970 22278 18972 22330
rect 18996 22278 19034 22330
rect 19034 22278 19046 22330
rect 19046 22278 19052 22330
rect 19076 22278 19098 22330
rect 19098 22278 19110 22330
rect 19110 22278 19132 22330
rect 19156 22278 19162 22330
rect 19162 22278 19174 22330
rect 19174 22278 19212 22330
rect 19236 22278 19238 22330
rect 19238 22278 19290 22330
rect 19290 22278 19292 22330
rect 18916 22276 18972 22278
rect 18996 22276 19052 22278
rect 19076 22276 19132 22278
rect 19156 22276 19212 22278
rect 19236 22276 19292 22278
rect 26916 22330 26972 22332
rect 26996 22330 27052 22332
rect 27076 22330 27132 22332
rect 27156 22330 27212 22332
rect 27236 22330 27292 22332
rect 26916 22278 26918 22330
rect 26918 22278 26970 22330
rect 26970 22278 26972 22330
rect 26996 22278 27034 22330
rect 27034 22278 27046 22330
rect 27046 22278 27052 22330
rect 27076 22278 27098 22330
rect 27098 22278 27110 22330
rect 27110 22278 27132 22330
rect 27156 22278 27162 22330
rect 27162 22278 27174 22330
rect 27174 22278 27212 22330
rect 27236 22278 27238 22330
rect 27238 22278 27290 22330
rect 27290 22278 27292 22330
rect 26916 22276 26972 22278
rect 26996 22276 27052 22278
rect 27076 22276 27132 22278
rect 27156 22276 27212 22278
rect 27236 22276 27292 22278
rect 28354 21800 28410 21856
rect 19656 21786 19712 21788
rect 19736 21786 19792 21788
rect 19816 21786 19872 21788
rect 19896 21786 19952 21788
rect 19976 21786 20032 21788
rect 19656 21734 19658 21786
rect 19658 21734 19710 21786
rect 19710 21734 19712 21786
rect 19736 21734 19774 21786
rect 19774 21734 19786 21786
rect 19786 21734 19792 21786
rect 19816 21734 19838 21786
rect 19838 21734 19850 21786
rect 19850 21734 19872 21786
rect 19896 21734 19902 21786
rect 19902 21734 19914 21786
rect 19914 21734 19952 21786
rect 19976 21734 19978 21786
rect 19978 21734 20030 21786
rect 20030 21734 20032 21786
rect 19656 21732 19712 21734
rect 19736 21732 19792 21734
rect 19816 21732 19872 21734
rect 19896 21732 19952 21734
rect 19976 21732 20032 21734
rect 27656 21786 27712 21788
rect 27736 21786 27792 21788
rect 27816 21786 27872 21788
rect 27896 21786 27952 21788
rect 27976 21786 28032 21788
rect 27656 21734 27658 21786
rect 27658 21734 27710 21786
rect 27710 21734 27712 21786
rect 27736 21734 27774 21786
rect 27774 21734 27786 21786
rect 27786 21734 27792 21786
rect 27816 21734 27838 21786
rect 27838 21734 27850 21786
rect 27850 21734 27872 21786
rect 27896 21734 27902 21786
rect 27902 21734 27914 21786
rect 27914 21734 27952 21786
rect 27976 21734 27978 21786
rect 27978 21734 28030 21786
rect 28030 21734 28032 21786
rect 27656 21732 27712 21734
rect 27736 21732 27792 21734
rect 27816 21732 27872 21734
rect 27896 21732 27952 21734
rect 27976 21732 28032 21734
rect 18916 21242 18972 21244
rect 18996 21242 19052 21244
rect 19076 21242 19132 21244
rect 19156 21242 19212 21244
rect 19236 21242 19292 21244
rect 18916 21190 18918 21242
rect 18918 21190 18970 21242
rect 18970 21190 18972 21242
rect 18996 21190 19034 21242
rect 19034 21190 19046 21242
rect 19046 21190 19052 21242
rect 19076 21190 19098 21242
rect 19098 21190 19110 21242
rect 19110 21190 19132 21242
rect 19156 21190 19162 21242
rect 19162 21190 19174 21242
rect 19174 21190 19212 21242
rect 19236 21190 19238 21242
rect 19238 21190 19290 21242
rect 19290 21190 19292 21242
rect 18916 21188 18972 21190
rect 18996 21188 19052 21190
rect 19076 21188 19132 21190
rect 19156 21188 19212 21190
rect 19236 21188 19292 21190
rect 26916 21242 26972 21244
rect 26996 21242 27052 21244
rect 27076 21242 27132 21244
rect 27156 21242 27212 21244
rect 27236 21242 27292 21244
rect 26916 21190 26918 21242
rect 26918 21190 26970 21242
rect 26970 21190 26972 21242
rect 26996 21190 27034 21242
rect 27034 21190 27046 21242
rect 27046 21190 27052 21242
rect 27076 21190 27098 21242
rect 27098 21190 27110 21242
rect 27110 21190 27132 21242
rect 27156 21190 27162 21242
rect 27162 21190 27174 21242
rect 27174 21190 27212 21242
rect 27236 21190 27238 21242
rect 27238 21190 27290 21242
rect 27290 21190 27292 21242
rect 26916 21188 26972 21190
rect 26996 21188 27052 21190
rect 27076 21188 27132 21190
rect 27156 21188 27212 21190
rect 27236 21188 27292 21190
rect 28354 20984 28410 21040
rect 19656 20698 19712 20700
rect 19736 20698 19792 20700
rect 19816 20698 19872 20700
rect 19896 20698 19952 20700
rect 19976 20698 20032 20700
rect 19656 20646 19658 20698
rect 19658 20646 19710 20698
rect 19710 20646 19712 20698
rect 19736 20646 19774 20698
rect 19774 20646 19786 20698
rect 19786 20646 19792 20698
rect 19816 20646 19838 20698
rect 19838 20646 19850 20698
rect 19850 20646 19872 20698
rect 19896 20646 19902 20698
rect 19902 20646 19914 20698
rect 19914 20646 19952 20698
rect 19976 20646 19978 20698
rect 19978 20646 20030 20698
rect 20030 20646 20032 20698
rect 19656 20644 19712 20646
rect 19736 20644 19792 20646
rect 19816 20644 19872 20646
rect 19896 20644 19952 20646
rect 19976 20644 20032 20646
rect 27656 20698 27712 20700
rect 27736 20698 27792 20700
rect 27816 20698 27872 20700
rect 27896 20698 27952 20700
rect 27976 20698 28032 20700
rect 27656 20646 27658 20698
rect 27658 20646 27710 20698
rect 27710 20646 27712 20698
rect 27736 20646 27774 20698
rect 27774 20646 27786 20698
rect 27786 20646 27792 20698
rect 27816 20646 27838 20698
rect 27838 20646 27850 20698
rect 27850 20646 27872 20698
rect 27896 20646 27902 20698
rect 27902 20646 27914 20698
rect 27914 20646 27952 20698
rect 27976 20646 27978 20698
rect 27978 20646 28030 20698
rect 28030 20646 28032 20698
rect 27656 20644 27712 20646
rect 27736 20644 27792 20646
rect 27816 20644 27872 20646
rect 27896 20644 27952 20646
rect 27976 20644 28032 20646
rect 28354 20168 28410 20224
rect 18916 20154 18972 20156
rect 18996 20154 19052 20156
rect 19076 20154 19132 20156
rect 19156 20154 19212 20156
rect 19236 20154 19292 20156
rect 18916 20102 18918 20154
rect 18918 20102 18970 20154
rect 18970 20102 18972 20154
rect 18996 20102 19034 20154
rect 19034 20102 19046 20154
rect 19046 20102 19052 20154
rect 19076 20102 19098 20154
rect 19098 20102 19110 20154
rect 19110 20102 19132 20154
rect 19156 20102 19162 20154
rect 19162 20102 19174 20154
rect 19174 20102 19212 20154
rect 19236 20102 19238 20154
rect 19238 20102 19290 20154
rect 19290 20102 19292 20154
rect 18916 20100 18972 20102
rect 18996 20100 19052 20102
rect 19076 20100 19132 20102
rect 19156 20100 19212 20102
rect 19236 20100 19292 20102
rect 26916 20154 26972 20156
rect 26996 20154 27052 20156
rect 27076 20154 27132 20156
rect 27156 20154 27212 20156
rect 27236 20154 27292 20156
rect 26916 20102 26918 20154
rect 26918 20102 26970 20154
rect 26970 20102 26972 20154
rect 26996 20102 27034 20154
rect 27034 20102 27046 20154
rect 27046 20102 27052 20154
rect 27076 20102 27098 20154
rect 27098 20102 27110 20154
rect 27110 20102 27132 20154
rect 27156 20102 27162 20154
rect 27162 20102 27174 20154
rect 27174 20102 27212 20154
rect 27236 20102 27238 20154
rect 27238 20102 27290 20154
rect 27290 20102 27292 20154
rect 26916 20100 26972 20102
rect 26996 20100 27052 20102
rect 27076 20100 27132 20102
rect 27156 20100 27212 20102
rect 27236 20100 27292 20102
rect 11656 18522 11712 18524
rect 11736 18522 11792 18524
rect 11816 18522 11872 18524
rect 11896 18522 11952 18524
rect 11976 18522 12032 18524
rect 11656 18470 11658 18522
rect 11658 18470 11710 18522
rect 11710 18470 11712 18522
rect 11736 18470 11774 18522
rect 11774 18470 11786 18522
rect 11786 18470 11792 18522
rect 11816 18470 11838 18522
rect 11838 18470 11850 18522
rect 11850 18470 11872 18522
rect 11896 18470 11902 18522
rect 11902 18470 11914 18522
rect 11914 18470 11952 18522
rect 11976 18470 11978 18522
rect 11978 18470 12030 18522
rect 12030 18470 12032 18522
rect 11656 18468 11712 18470
rect 11736 18468 11792 18470
rect 11816 18468 11872 18470
rect 11896 18468 11952 18470
rect 11976 18468 12032 18470
rect 11656 17434 11712 17436
rect 11736 17434 11792 17436
rect 11816 17434 11872 17436
rect 11896 17434 11952 17436
rect 11976 17434 12032 17436
rect 11656 17382 11658 17434
rect 11658 17382 11710 17434
rect 11710 17382 11712 17434
rect 11736 17382 11774 17434
rect 11774 17382 11786 17434
rect 11786 17382 11792 17434
rect 11816 17382 11838 17434
rect 11838 17382 11850 17434
rect 11850 17382 11872 17434
rect 11896 17382 11902 17434
rect 11902 17382 11914 17434
rect 11914 17382 11952 17434
rect 11976 17382 11978 17434
rect 11978 17382 12030 17434
rect 12030 17382 12032 17434
rect 11656 17380 11712 17382
rect 11736 17380 11792 17382
rect 11816 17380 11872 17382
rect 11896 17380 11952 17382
rect 11976 17380 12032 17382
rect 11656 16346 11712 16348
rect 11736 16346 11792 16348
rect 11816 16346 11872 16348
rect 11896 16346 11952 16348
rect 11976 16346 12032 16348
rect 11656 16294 11658 16346
rect 11658 16294 11710 16346
rect 11710 16294 11712 16346
rect 11736 16294 11774 16346
rect 11774 16294 11786 16346
rect 11786 16294 11792 16346
rect 11816 16294 11838 16346
rect 11838 16294 11850 16346
rect 11850 16294 11872 16346
rect 11896 16294 11902 16346
rect 11902 16294 11914 16346
rect 11914 16294 11952 16346
rect 11976 16294 11978 16346
rect 11978 16294 12030 16346
rect 12030 16294 12032 16346
rect 11656 16292 11712 16294
rect 11736 16292 11792 16294
rect 11816 16292 11872 16294
rect 11896 16292 11952 16294
rect 11976 16292 12032 16294
rect 11610 15428 11666 15464
rect 11610 15408 11612 15428
rect 11612 15408 11664 15428
rect 11664 15408 11666 15428
rect 11656 15258 11712 15260
rect 11736 15258 11792 15260
rect 11816 15258 11872 15260
rect 11896 15258 11952 15260
rect 11976 15258 12032 15260
rect 11656 15206 11658 15258
rect 11658 15206 11710 15258
rect 11710 15206 11712 15258
rect 11736 15206 11774 15258
rect 11774 15206 11786 15258
rect 11786 15206 11792 15258
rect 11816 15206 11838 15258
rect 11838 15206 11850 15258
rect 11850 15206 11872 15258
rect 11896 15206 11902 15258
rect 11902 15206 11914 15258
rect 11914 15206 11952 15258
rect 11976 15206 11978 15258
rect 11978 15206 12030 15258
rect 12030 15206 12032 15258
rect 11656 15204 11712 15206
rect 11736 15204 11792 15206
rect 11816 15204 11872 15206
rect 11896 15204 11952 15206
rect 11976 15204 12032 15206
rect 1398 14864 1454 14920
rect 2916 14714 2972 14716
rect 2996 14714 3052 14716
rect 3076 14714 3132 14716
rect 3156 14714 3212 14716
rect 3236 14714 3292 14716
rect 2916 14662 2918 14714
rect 2918 14662 2970 14714
rect 2970 14662 2972 14714
rect 2996 14662 3034 14714
rect 3034 14662 3046 14714
rect 3046 14662 3052 14714
rect 3076 14662 3098 14714
rect 3098 14662 3110 14714
rect 3110 14662 3132 14714
rect 3156 14662 3162 14714
rect 3162 14662 3174 14714
rect 3174 14662 3212 14714
rect 3236 14662 3238 14714
rect 3238 14662 3290 14714
rect 3290 14662 3292 14714
rect 2916 14660 2972 14662
rect 2996 14660 3052 14662
rect 3076 14660 3132 14662
rect 3156 14660 3212 14662
rect 3236 14660 3292 14662
rect 10916 14714 10972 14716
rect 10996 14714 11052 14716
rect 11076 14714 11132 14716
rect 11156 14714 11212 14716
rect 11236 14714 11292 14716
rect 10916 14662 10918 14714
rect 10918 14662 10970 14714
rect 10970 14662 10972 14714
rect 10996 14662 11034 14714
rect 11034 14662 11046 14714
rect 11046 14662 11052 14714
rect 11076 14662 11098 14714
rect 11098 14662 11110 14714
rect 11110 14662 11132 14714
rect 11156 14662 11162 14714
rect 11162 14662 11174 14714
rect 11174 14662 11212 14714
rect 11236 14662 11238 14714
rect 11238 14662 11290 14714
rect 11290 14662 11292 14714
rect 10916 14660 10972 14662
rect 10996 14660 11052 14662
rect 11076 14660 11132 14662
rect 11156 14660 11212 14662
rect 11236 14660 11292 14662
rect 3656 14170 3712 14172
rect 3736 14170 3792 14172
rect 3816 14170 3872 14172
rect 3896 14170 3952 14172
rect 3976 14170 4032 14172
rect 3656 14118 3658 14170
rect 3658 14118 3710 14170
rect 3710 14118 3712 14170
rect 3736 14118 3774 14170
rect 3774 14118 3786 14170
rect 3786 14118 3792 14170
rect 3816 14118 3838 14170
rect 3838 14118 3850 14170
rect 3850 14118 3872 14170
rect 3896 14118 3902 14170
rect 3902 14118 3914 14170
rect 3914 14118 3952 14170
rect 3976 14118 3978 14170
rect 3978 14118 4030 14170
rect 4030 14118 4032 14170
rect 3656 14116 3712 14118
rect 3736 14116 3792 14118
rect 3816 14116 3872 14118
rect 3896 14116 3952 14118
rect 3976 14116 4032 14118
rect 1398 14048 1454 14104
rect 2916 13626 2972 13628
rect 2996 13626 3052 13628
rect 3076 13626 3132 13628
rect 3156 13626 3212 13628
rect 3236 13626 3292 13628
rect 2916 13574 2918 13626
rect 2918 13574 2970 13626
rect 2970 13574 2972 13626
rect 2996 13574 3034 13626
rect 3034 13574 3046 13626
rect 3046 13574 3052 13626
rect 3076 13574 3098 13626
rect 3098 13574 3110 13626
rect 3110 13574 3132 13626
rect 3156 13574 3162 13626
rect 3162 13574 3174 13626
rect 3174 13574 3212 13626
rect 3236 13574 3238 13626
rect 3238 13574 3290 13626
rect 3290 13574 3292 13626
rect 2916 13572 2972 13574
rect 2996 13572 3052 13574
rect 3076 13572 3132 13574
rect 3156 13572 3212 13574
rect 3236 13572 3292 13574
rect 1398 13268 1400 13288
rect 1400 13268 1452 13288
rect 1452 13268 1454 13288
rect 1398 13232 1454 13268
rect 3656 13082 3712 13084
rect 3736 13082 3792 13084
rect 3816 13082 3872 13084
rect 3896 13082 3952 13084
rect 3976 13082 4032 13084
rect 3656 13030 3658 13082
rect 3658 13030 3710 13082
rect 3710 13030 3712 13082
rect 3736 13030 3774 13082
rect 3774 13030 3786 13082
rect 3786 13030 3792 13082
rect 3816 13030 3838 13082
rect 3838 13030 3850 13082
rect 3850 13030 3872 13082
rect 3896 13030 3902 13082
rect 3902 13030 3914 13082
rect 3914 13030 3952 13082
rect 3976 13030 3978 13082
rect 3978 13030 4030 13082
rect 4030 13030 4032 13082
rect 3656 13028 3712 13030
rect 3736 13028 3792 13030
rect 3816 13028 3872 13030
rect 3896 13028 3952 13030
rect 3976 13028 4032 13030
rect 2916 12538 2972 12540
rect 2996 12538 3052 12540
rect 3076 12538 3132 12540
rect 3156 12538 3212 12540
rect 3236 12538 3292 12540
rect 2916 12486 2918 12538
rect 2918 12486 2970 12538
rect 2970 12486 2972 12538
rect 2996 12486 3034 12538
rect 3034 12486 3046 12538
rect 3046 12486 3052 12538
rect 3076 12486 3098 12538
rect 3098 12486 3110 12538
rect 3110 12486 3132 12538
rect 3156 12486 3162 12538
rect 3162 12486 3174 12538
rect 3174 12486 3212 12538
rect 3236 12486 3238 12538
rect 3238 12486 3290 12538
rect 3290 12486 3292 12538
rect 2916 12484 2972 12486
rect 2996 12484 3052 12486
rect 3076 12484 3132 12486
rect 3156 12484 3212 12486
rect 3236 12484 3292 12486
rect 1398 12416 1454 12472
rect 3656 11994 3712 11996
rect 3736 11994 3792 11996
rect 3816 11994 3872 11996
rect 3896 11994 3952 11996
rect 3976 11994 4032 11996
rect 3656 11942 3658 11994
rect 3658 11942 3710 11994
rect 3710 11942 3712 11994
rect 3736 11942 3774 11994
rect 3774 11942 3786 11994
rect 3786 11942 3792 11994
rect 3816 11942 3838 11994
rect 3838 11942 3850 11994
rect 3850 11942 3872 11994
rect 3896 11942 3902 11994
rect 3902 11942 3914 11994
rect 3914 11942 3952 11994
rect 3976 11942 3978 11994
rect 3978 11942 4030 11994
rect 4030 11942 4032 11994
rect 3656 11940 3712 11942
rect 3736 11940 3792 11942
rect 3816 11940 3872 11942
rect 3896 11940 3952 11942
rect 3976 11940 4032 11942
rect 1398 11600 1454 11656
rect 2916 11450 2972 11452
rect 2996 11450 3052 11452
rect 3076 11450 3132 11452
rect 3156 11450 3212 11452
rect 3236 11450 3292 11452
rect 2916 11398 2918 11450
rect 2918 11398 2970 11450
rect 2970 11398 2972 11450
rect 2996 11398 3034 11450
rect 3034 11398 3046 11450
rect 3046 11398 3052 11450
rect 3076 11398 3098 11450
rect 3098 11398 3110 11450
rect 3110 11398 3132 11450
rect 3156 11398 3162 11450
rect 3162 11398 3174 11450
rect 3174 11398 3212 11450
rect 3236 11398 3238 11450
rect 3238 11398 3290 11450
rect 3290 11398 3292 11450
rect 2916 11396 2972 11398
rect 2996 11396 3052 11398
rect 3076 11396 3132 11398
rect 3156 11396 3212 11398
rect 3236 11396 3292 11398
rect 3656 10906 3712 10908
rect 3736 10906 3792 10908
rect 3816 10906 3872 10908
rect 3896 10906 3952 10908
rect 3976 10906 4032 10908
rect 3656 10854 3658 10906
rect 3658 10854 3710 10906
rect 3710 10854 3712 10906
rect 3736 10854 3774 10906
rect 3774 10854 3786 10906
rect 3786 10854 3792 10906
rect 3816 10854 3838 10906
rect 3838 10854 3850 10906
rect 3850 10854 3872 10906
rect 3896 10854 3902 10906
rect 3902 10854 3914 10906
rect 3914 10854 3952 10906
rect 3976 10854 3978 10906
rect 3978 10854 4030 10906
rect 4030 10854 4032 10906
rect 3656 10852 3712 10854
rect 3736 10852 3792 10854
rect 3816 10852 3872 10854
rect 3896 10852 3952 10854
rect 3976 10852 4032 10854
rect 1398 10784 1454 10840
rect 11656 14170 11712 14172
rect 11736 14170 11792 14172
rect 11816 14170 11872 14172
rect 11896 14170 11952 14172
rect 11976 14170 12032 14172
rect 11656 14118 11658 14170
rect 11658 14118 11710 14170
rect 11710 14118 11712 14170
rect 11736 14118 11774 14170
rect 11774 14118 11786 14170
rect 11786 14118 11792 14170
rect 11816 14118 11838 14170
rect 11838 14118 11850 14170
rect 11850 14118 11872 14170
rect 11896 14118 11902 14170
rect 11902 14118 11914 14170
rect 11914 14118 11952 14170
rect 11976 14118 11978 14170
rect 11978 14118 12030 14170
rect 12030 14118 12032 14170
rect 11656 14116 11712 14118
rect 11736 14116 11792 14118
rect 11816 14116 11872 14118
rect 11896 14116 11952 14118
rect 11976 14116 12032 14118
rect 10916 13626 10972 13628
rect 10996 13626 11052 13628
rect 11076 13626 11132 13628
rect 11156 13626 11212 13628
rect 11236 13626 11292 13628
rect 10916 13574 10918 13626
rect 10918 13574 10970 13626
rect 10970 13574 10972 13626
rect 10996 13574 11034 13626
rect 11034 13574 11046 13626
rect 11046 13574 11052 13626
rect 11076 13574 11098 13626
rect 11098 13574 11110 13626
rect 11110 13574 11132 13626
rect 11156 13574 11162 13626
rect 11162 13574 11174 13626
rect 11174 13574 11212 13626
rect 11236 13574 11238 13626
rect 11238 13574 11290 13626
rect 11290 13574 11292 13626
rect 10916 13572 10972 13574
rect 10996 13572 11052 13574
rect 11076 13572 11132 13574
rect 11156 13572 11212 13574
rect 11236 13572 11292 13574
rect 11656 13082 11712 13084
rect 11736 13082 11792 13084
rect 11816 13082 11872 13084
rect 11896 13082 11952 13084
rect 11976 13082 12032 13084
rect 11656 13030 11658 13082
rect 11658 13030 11710 13082
rect 11710 13030 11712 13082
rect 11736 13030 11774 13082
rect 11774 13030 11786 13082
rect 11786 13030 11792 13082
rect 11816 13030 11838 13082
rect 11838 13030 11850 13082
rect 11850 13030 11872 13082
rect 11896 13030 11902 13082
rect 11902 13030 11914 13082
rect 11914 13030 11952 13082
rect 11976 13030 11978 13082
rect 11978 13030 12030 13082
rect 12030 13030 12032 13082
rect 11656 13028 11712 13030
rect 11736 13028 11792 13030
rect 11816 13028 11872 13030
rect 11896 13028 11952 13030
rect 11976 13028 12032 13030
rect 2916 10362 2972 10364
rect 2996 10362 3052 10364
rect 3076 10362 3132 10364
rect 3156 10362 3212 10364
rect 3236 10362 3292 10364
rect 2916 10310 2918 10362
rect 2918 10310 2970 10362
rect 2970 10310 2972 10362
rect 2996 10310 3034 10362
rect 3034 10310 3046 10362
rect 3046 10310 3052 10362
rect 3076 10310 3098 10362
rect 3098 10310 3110 10362
rect 3110 10310 3132 10362
rect 3156 10310 3162 10362
rect 3162 10310 3174 10362
rect 3174 10310 3212 10362
rect 3236 10310 3238 10362
rect 3238 10310 3290 10362
rect 3290 10310 3292 10362
rect 2916 10308 2972 10310
rect 2996 10308 3052 10310
rect 3076 10308 3132 10310
rect 3156 10308 3212 10310
rect 3236 10308 3292 10310
rect 10916 12538 10972 12540
rect 10996 12538 11052 12540
rect 11076 12538 11132 12540
rect 11156 12538 11212 12540
rect 11236 12538 11292 12540
rect 10916 12486 10918 12538
rect 10918 12486 10970 12538
rect 10970 12486 10972 12538
rect 10996 12486 11034 12538
rect 11034 12486 11046 12538
rect 11046 12486 11052 12538
rect 11076 12486 11098 12538
rect 11098 12486 11110 12538
rect 11110 12486 11132 12538
rect 11156 12486 11162 12538
rect 11162 12486 11174 12538
rect 11174 12486 11212 12538
rect 11236 12486 11238 12538
rect 11238 12486 11290 12538
rect 11290 12486 11292 12538
rect 10916 12484 10972 12486
rect 10996 12484 11052 12486
rect 11076 12484 11132 12486
rect 11156 12484 11212 12486
rect 11236 12484 11292 12486
rect 19656 19610 19712 19612
rect 19736 19610 19792 19612
rect 19816 19610 19872 19612
rect 19896 19610 19952 19612
rect 19976 19610 20032 19612
rect 19656 19558 19658 19610
rect 19658 19558 19710 19610
rect 19710 19558 19712 19610
rect 19736 19558 19774 19610
rect 19774 19558 19786 19610
rect 19786 19558 19792 19610
rect 19816 19558 19838 19610
rect 19838 19558 19850 19610
rect 19850 19558 19872 19610
rect 19896 19558 19902 19610
rect 19902 19558 19914 19610
rect 19914 19558 19952 19610
rect 19976 19558 19978 19610
rect 19978 19558 20030 19610
rect 20030 19558 20032 19610
rect 19656 19556 19712 19558
rect 19736 19556 19792 19558
rect 19816 19556 19872 19558
rect 19896 19556 19952 19558
rect 19976 19556 20032 19558
rect 27656 19610 27712 19612
rect 27736 19610 27792 19612
rect 27816 19610 27872 19612
rect 27896 19610 27952 19612
rect 27976 19610 28032 19612
rect 27656 19558 27658 19610
rect 27658 19558 27710 19610
rect 27710 19558 27712 19610
rect 27736 19558 27774 19610
rect 27774 19558 27786 19610
rect 27786 19558 27792 19610
rect 27816 19558 27838 19610
rect 27838 19558 27850 19610
rect 27850 19558 27872 19610
rect 27896 19558 27902 19610
rect 27902 19558 27914 19610
rect 27914 19558 27952 19610
rect 27976 19558 27978 19610
rect 27978 19558 28030 19610
rect 28030 19558 28032 19610
rect 27656 19556 27712 19558
rect 27736 19556 27792 19558
rect 27816 19556 27872 19558
rect 27896 19556 27952 19558
rect 27976 19556 28032 19558
rect 28354 19352 28410 19408
rect 18916 19066 18972 19068
rect 18996 19066 19052 19068
rect 19076 19066 19132 19068
rect 19156 19066 19212 19068
rect 19236 19066 19292 19068
rect 18916 19014 18918 19066
rect 18918 19014 18970 19066
rect 18970 19014 18972 19066
rect 18996 19014 19034 19066
rect 19034 19014 19046 19066
rect 19046 19014 19052 19066
rect 19076 19014 19098 19066
rect 19098 19014 19110 19066
rect 19110 19014 19132 19066
rect 19156 19014 19162 19066
rect 19162 19014 19174 19066
rect 19174 19014 19212 19066
rect 19236 19014 19238 19066
rect 19238 19014 19290 19066
rect 19290 19014 19292 19066
rect 18916 19012 18972 19014
rect 18996 19012 19052 19014
rect 19076 19012 19132 19014
rect 19156 19012 19212 19014
rect 19236 19012 19292 19014
rect 26916 19066 26972 19068
rect 26996 19066 27052 19068
rect 27076 19066 27132 19068
rect 27156 19066 27212 19068
rect 27236 19066 27292 19068
rect 26916 19014 26918 19066
rect 26918 19014 26970 19066
rect 26970 19014 26972 19066
rect 26996 19014 27034 19066
rect 27034 19014 27046 19066
rect 27046 19014 27052 19066
rect 27076 19014 27098 19066
rect 27098 19014 27110 19066
rect 27110 19014 27132 19066
rect 27156 19014 27162 19066
rect 27162 19014 27174 19066
rect 27174 19014 27212 19066
rect 27236 19014 27238 19066
rect 27238 19014 27290 19066
rect 27290 19014 27292 19066
rect 26916 19012 26972 19014
rect 26996 19012 27052 19014
rect 27076 19012 27132 19014
rect 27156 19012 27212 19014
rect 27236 19012 27292 19014
rect 28354 18536 28410 18592
rect 19656 18522 19712 18524
rect 19736 18522 19792 18524
rect 19816 18522 19872 18524
rect 19896 18522 19952 18524
rect 19976 18522 20032 18524
rect 19656 18470 19658 18522
rect 19658 18470 19710 18522
rect 19710 18470 19712 18522
rect 19736 18470 19774 18522
rect 19774 18470 19786 18522
rect 19786 18470 19792 18522
rect 19816 18470 19838 18522
rect 19838 18470 19850 18522
rect 19850 18470 19872 18522
rect 19896 18470 19902 18522
rect 19902 18470 19914 18522
rect 19914 18470 19952 18522
rect 19976 18470 19978 18522
rect 19978 18470 20030 18522
rect 20030 18470 20032 18522
rect 19656 18468 19712 18470
rect 19736 18468 19792 18470
rect 19816 18468 19872 18470
rect 19896 18468 19952 18470
rect 19976 18468 20032 18470
rect 27656 18522 27712 18524
rect 27736 18522 27792 18524
rect 27816 18522 27872 18524
rect 27896 18522 27952 18524
rect 27976 18522 28032 18524
rect 27656 18470 27658 18522
rect 27658 18470 27710 18522
rect 27710 18470 27712 18522
rect 27736 18470 27774 18522
rect 27774 18470 27786 18522
rect 27786 18470 27792 18522
rect 27816 18470 27838 18522
rect 27838 18470 27850 18522
rect 27850 18470 27872 18522
rect 27896 18470 27902 18522
rect 27902 18470 27914 18522
rect 27914 18470 27952 18522
rect 27976 18470 27978 18522
rect 27978 18470 28030 18522
rect 28030 18470 28032 18522
rect 27656 18468 27712 18470
rect 27736 18468 27792 18470
rect 27816 18468 27872 18470
rect 27896 18468 27952 18470
rect 27976 18468 28032 18470
rect 18916 17978 18972 17980
rect 18996 17978 19052 17980
rect 19076 17978 19132 17980
rect 19156 17978 19212 17980
rect 19236 17978 19292 17980
rect 18916 17926 18918 17978
rect 18918 17926 18970 17978
rect 18970 17926 18972 17978
rect 18996 17926 19034 17978
rect 19034 17926 19046 17978
rect 19046 17926 19052 17978
rect 19076 17926 19098 17978
rect 19098 17926 19110 17978
rect 19110 17926 19132 17978
rect 19156 17926 19162 17978
rect 19162 17926 19174 17978
rect 19174 17926 19212 17978
rect 19236 17926 19238 17978
rect 19238 17926 19290 17978
rect 19290 17926 19292 17978
rect 18916 17924 18972 17926
rect 18996 17924 19052 17926
rect 19076 17924 19132 17926
rect 19156 17924 19212 17926
rect 19236 17924 19292 17926
rect 26916 17978 26972 17980
rect 26996 17978 27052 17980
rect 27076 17978 27132 17980
rect 27156 17978 27212 17980
rect 27236 17978 27292 17980
rect 26916 17926 26918 17978
rect 26918 17926 26970 17978
rect 26970 17926 26972 17978
rect 26996 17926 27034 17978
rect 27034 17926 27046 17978
rect 27046 17926 27052 17978
rect 27076 17926 27098 17978
rect 27098 17926 27110 17978
rect 27110 17926 27132 17978
rect 27156 17926 27162 17978
rect 27162 17926 27174 17978
rect 27174 17926 27212 17978
rect 27236 17926 27238 17978
rect 27238 17926 27290 17978
rect 27290 17926 27292 17978
rect 26916 17924 26972 17926
rect 26996 17924 27052 17926
rect 27076 17924 27132 17926
rect 27156 17924 27212 17926
rect 27236 17924 27292 17926
rect 28354 17720 28410 17776
rect 19656 17434 19712 17436
rect 19736 17434 19792 17436
rect 19816 17434 19872 17436
rect 19896 17434 19952 17436
rect 19976 17434 20032 17436
rect 19656 17382 19658 17434
rect 19658 17382 19710 17434
rect 19710 17382 19712 17434
rect 19736 17382 19774 17434
rect 19774 17382 19786 17434
rect 19786 17382 19792 17434
rect 19816 17382 19838 17434
rect 19838 17382 19850 17434
rect 19850 17382 19872 17434
rect 19896 17382 19902 17434
rect 19902 17382 19914 17434
rect 19914 17382 19952 17434
rect 19976 17382 19978 17434
rect 19978 17382 20030 17434
rect 20030 17382 20032 17434
rect 19656 17380 19712 17382
rect 19736 17380 19792 17382
rect 19816 17380 19872 17382
rect 19896 17380 19952 17382
rect 19976 17380 20032 17382
rect 27656 17434 27712 17436
rect 27736 17434 27792 17436
rect 27816 17434 27872 17436
rect 27896 17434 27952 17436
rect 27976 17434 28032 17436
rect 27656 17382 27658 17434
rect 27658 17382 27710 17434
rect 27710 17382 27712 17434
rect 27736 17382 27774 17434
rect 27774 17382 27786 17434
rect 27786 17382 27792 17434
rect 27816 17382 27838 17434
rect 27838 17382 27850 17434
rect 27850 17382 27872 17434
rect 27896 17382 27902 17434
rect 27902 17382 27914 17434
rect 27914 17382 27952 17434
rect 27976 17382 27978 17434
rect 27978 17382 28030 17434
rect 28030 17382 28032 17434
rect 27656 17380 27712 17382
rect 27736 17380 27792 17382
rect 27816 17380 27872 17382
rect 27896 17380 27952 17382
rect 27976 17380 28032 17382
rect 28354 16904 28410 16960
rect 18916 16890 18972 16892
rect 18996 16890 19052 16892
rect 19076 16890 19132 16892
rect 19156 16890 19212 16892
rect 19236 16890 19292 16892
rect 18916 16838 18918 16890
rect 18918 16838 18970 16890
rect 18970 16838 18972 16890
rect 18996 16838 19034 16890
rect 19034 16838 19046 16890
rect 19046 16838 19052 16890
rect 19076 16838 19098 16890
rect 19098 16838 19110 16890
rect 19110 16838 19132 16890
rect 19156 16838 19162 16890
rect 19162 16838 19174 16890
rect 19174 16838 19212 16890
rect 19236 16838 19238 16890
rect 19238 16838 19290 16890
rect 19290 16838 19292 16890
rect 18916 16836 18972 16838
rect 18996 16836 19052 16838
rect 19076 16836 19132 16838
rect 19156 16836 19212 16838
rect 19236 16836 19292 16838
rect 26916 16890 26972 16892
rect 26996 16890 27052 16892
rect 27076 16890 27132 16892
rect 27156 16890 27212 16892
rect 27236 16890 27292 16892
rect 26916 16838 26918 16890
rect 26918 16838 26970 16890
rect 26970 16838 26972 16890
rect 26996 16838 27034 16890
rect 27034 16838 27046 16890
rect 27046 16838 27052 16890
rect 27076 16838 27098 16890
rect 27098 16838 27110 16890
rect 27110 16838 27132 16890
rect 27156 16838 27162 16890
rect 27162 16838 27174 16890
rect 27174 16838 27212 16890
rect 27236 16838 27238 16890
rect 27238 16838 27290 16890
rect 27290 16838 27292 16890
rect 26916 16836 26972 16838
rect 26996 16836 27052 16838
rect 27076 16836 27132 16838
rect 27156 16836 27212 16838
rect 27236 16836 27292 16838
rect 19656 16346 19712 16348
rect 19736 16346 19792 16348
rect 19816 16346 19872 16348
rect 19896 16346 19952 16348
rect 19976 16346 20032 16348
rect 19656 16294 19658 16346
rect 19658 16294 19710 16346
rect 19710 16294 19712 16346
rect 19736 16294 19774 16346
rect 19774 16294 19786 16346
rect 19786 16294 19792 16346
rect 19816 16294 19838 16346
rect 19838 16294 19850 16346
rect 19850 16294 19872 16346
rect 19896 16294 19902 16346
rect 19902 16294 19914 16346
rect 19914 16294 19952 16346
rect 19976 16294 19978 16346
rect 19978 16294 20030 16346
rect 20030 16294 20032 16346
rect 19656 16292 19712 16294
rect 19736 16292 19792 16294
rect 19816 16292 19872 16294
rect 19896 16292 19952 16294
rect 19976 16292 20032 16294
rect 18916 15802 18972 15804
rect 18996 15802 19052 15804
rect 19076 15802 19132 15804
rect 19156 15802 19212 15804
rect 19236 15802 19292 15804
rect 18916 15750 18918 15802
rect 18918 15750 18970 15802
rect 18970 15750 18972 15802
rect 18996 15750 19034 15802
rect 19034 15750 19046 15802
rect 19046 15750 19052 15802
rect 19076 15750 19098 15802
rect 19098 15750 19110 15802
rect 19110 15750 19132 15802
rect 19156 15750 19162 15802
rect 19162 15750 19174 15802
rect 19174 15750 19212 15802
rect 19236 15750 19238 15802
rect 19238 15750 19290 15802
rect 19290 15750 19292 15802
rect 18916 15748 18972 15750
rect 18996 15748 19052 15750
rect 19076 15748 19132 15750
rect 19156 15748 19212 15750
rect 19236 15748 19292 15750
rect 27656 16346 27712 16348
rect 27736 16346 27792 16348
rect 27816 16346 27872 16348
rect 27896 16346 27952 16348
rect 27976 16346 28032 16348
rect 27656 16294 27658 16346
rect 27658 16294 27710 16346
rect 27710 16294 27712 16346
rect 27736 16294 27774 16346
rect 27774 16294 27786 16346
rect 27786 16294 27792 16346
rect 27816 16294 27838 16346
rect 27838 16294 27850 16346
rect 27850 16294 27872 16346
rect 27896 16294 27902 16346
rect 27902 16294 27914 16346
rect 27914 16294 27952 16346
rect 27976 16294 27978 16346
rect 27978 16294 28030 16346
rect 28030 16294 28032 16346
rect 27656 16292 27712 16294
rect 27736 16292 27792 16294
rect 27816 16292 27872 16294
rect 27896 16292 27952 16294
rect 27976 16292 28032 16294
rect 28354 16088 28410 16144
rect 26916 15802 26972 15804
rect 26996 15802 27052 15804
rect 27076 15802 27132 15804
rect 27156 15802 27212 15804
rect 27236 15802 27292 15804
rect 26916 15750 26918 15802
rect 26918 15750 26970 15802
rect 26970 15750 26972 15802
rect 26996 15750 27034 15802
rect 27034 15750 27046 15802
rect 27046 15750 27052 15802
rect 27076 15750 27098 15802
rect 27098 15750 27110 15802
rect 27110 15750 27132 15802
rect 27156 15750 27162 15802
rect 27162 15750 27174 15802
rect 27174 15750 27212 15802
rect 27236 15750 27238 15802
rect 27238 15750 27290 15802
rect 27290 15750 27292 15802
rect 26916 15748 26972 15750
rect 26996 15748 27052 15750
rect 27076 15748 27132 15750
rect 27156 15748 27212 15750
rect 27236 15748 27292 15750
rect 28354 15272 28410 15328
rect 19656 15258 19712 15260
rect 19736 15258 19792 15260
rect 19816 15258 19872 15260
rect 19896 15258 19952 15260
rect 19976 15258 20032 15260
rect 19656 15206 19658 15258
rect 19658 15206 19710 15258
rect 19710 15206 19712 15258
rect 19736 15206 19774 15258
rect 19774 15206 19786 15258
rect 19786 15206 19792 15258
rect 19816 15206 19838 15258
rect 19838 15206 19850 15258
rect 19850 15206 19872 15258
rect 19896 15206 19902 15258
rect 19902 15206 19914 15258
rect 19914 15206 19952 15258
rect 19976 15206 19978 15258
rect 19978 15206 20030 15258
rect 20030 15206 20032 15258
rect 19656 15204 19712 15206
rect 19736 15204 19792 15206
rect 19816 15204 19872 15206
rect 19896 15204 19952 15206
rect 19976 15204 20032 15206
rect 27656 15258 27712 15260
rect 27736 15258 27792 15260
rect 27816 15258 27872 15260
rect 27896 15258 27952 15260
rect 27976 15258 28032 15260
rect 27656 15206 27658 15258
rect 27658 15206 27710 15258
rect 27710 15206 27712 15258
rect 27736 15206 27774 15258
rect 27774 15206 27786 15258
rect 27786 15206 27792 15258
rect 27816 15206 27838 15258
rect 27838 15206 27850 15258
rect 27850 15206 27872 15258
rect 27896 15206 27902 15258
rect 27902 15206 27914 15258
rect 27914 15206 27952 15258
rect 27976 15206 27978 15258
rect 27978 15206 28030 15258
rect 28030 15206 28032 15258
rect 27656 15204 27712 15206
rect 27736 15204 27792 15206
rect 27816 15204 27872 15206
rect 27896 15204 27952 15206
rect 27976 15204 28032 15206
rect 11656 11994 11712 11996
rect 11736 11994 11792 11996
rect 11816 11994 11872 11996
rect 11896 11994 11952 11996
rect 11976 11994 12032 11996
rect 11656 11942 11658 11994
rect 11658 11942 11710 11994
rect 11710 11942 11712 11994
rect 11736 11942 11774 11994
rect 11774 11942 11786 11994
rect 11786 11942 11792 11994
rect 11816 11942 11838 11994
rect 11838 11942 11850 11994
rect 11850 11942 11872 11994
rect 11896 11942 11902 11994
rect 11902 11942 11914 11994
rect 11914 11942 11952 11994
rect 11976 11942 11978 11994
rect 11978 11942 12030 11994
rect 12030 11942 12032 11994
rect 11656 11940 11712 11942
rect 11736 11940 11792 11942
rect 11816 11940 11872 11942
rect 11896 11940 11952 11942
rect 11976 11940 12032 11942
rect 10916 11450 10972 11452
rect 10996 11450 11052 11452
rect 11076 11450 11132 11452
rect 11156 11450 11212 11452
rect 11236 11450 11292 11452
rect 10916 11398 10918 11450
rect 10918 11398 10970 11450
rect 10970 11398 10972 11450
rect 10996 11398 11034 11450
rect 11034 11398 11046 11450
rect 11046 11398 11052 11450
rect 11076 11398 11098 11450
rect 11098 11398 11110 11450
rect 11110 11398 11132 11450
rect 11156 11398 11162 11450
rect 11162 11398 11174 11450
rect 11174 11398 11212 11450
rect 11236 11398 11238 11450
rect 11238 11398 11290 11450
rect 11290 11398 11292 11450
rect 10916 11396 10972 11398
rect 10996 11396 11052 11398
rect 11076 11396 11132 11398
rect 11156 11396 11212 11398
rect 11236 11396 11292 11398
rect 1398 9832 1454 9888
rect 3656 9818 3712 9820
rect 3736 9818 3792 9820
rect 3816 9818 3872 9820
rect 3896 9818 3952 9820
rect 3976 9818 4032 9820
rect 3656 9766 3658 9818
rect 3658 9766 3710 9818
rect 3710 9766 3712 9818
rect 3736 9766 3774 9818
rect 3774 9766 3786 9818
rect 3786 9766 3792 9818
rect 3816 9766 3838 9818
rect 3838 9766 3850 9818
rect 3850 9766 3872 9818
rect 3896 9766 3902 9818
rect 3902 9766 3914 9818
rect 3914 9766 3952 9818
rect 3976 9766 3978 9818
rect 3978 9766 4030 9818
rect 4030 9766 4032 9818
rect 3656 9764 3712 9766
rect 3736 9764 3792 9766
rect 3816 9764 3872 9766
rect 3896 9764 3952 9766
rect 3976 9764 4032 9766
rect 10916 10362 10972 10364
rect 10996 10362 11052 10364
rect 11076 10362 11132 10364
rect 11156 10362 11212 10364
rect 11236 10362 11292 10364
rect 10916 10310 10918 10362
rect 10918 10310 10970 10362
rect 10970 10310 10972 10362
rect 10996 10310 11034 10362
rect 11034 10310 11046 10362
rect 11046 10310 11052 10362
rect 11076 10310 11098 10362
rect 11098 10310 11110 10362
rect 11110 10310 11132 10362
rect 11156 10310 11162 10362
rect 11162 10310 11174 10362
rect 11174 10310 11212 10362
rect 11236 10310 11238 10362
rect 11238 10310 11290 10362
rect 11290 10310 11292 10362
rect 10916 10308 10972 10310
rect 10996 10308 11052 10310
rect 11076 10308 11132 10310
rect 11156 10308 11212 10310
rect 11236 10308 11292 10310
rect 2916 9274 2972 9276
rect 2996 9274 3052 9276
rect 3076 9274 3132 9276
rect 3156 9274 3212 9276
rect 3236 9274 3292 9276
rect 2916 9222 2918 9274
rect 2918 9222 2970 9274
rect 2970 9222 2972 9274
rect 2996 9222 3034 9274
rect 3034 9222 3046 9274
rect 3046 9222 3052 9274
rect 3076 9222 3098 9274
rect 3098 9222 3110 9274
rect 3110 9222 3132 9274
rect 3156 9222 3162 9274
rect 3162 9222 3174 9274
rect 3174 9222 3212 9274
rect 3236 9222 3238 9274
rect 3238 9222 3290 9274
rect 3290 9222 3292 9274
rect 2916 9220 2972 9222
rect 2996 9220 3052 9222
rect 3076 9220 3132 9222
rect 3156 9220 3212 9222
rect 3236 9220 3292 9222
rect 1398 9152 1454 9208
rect 3656 8730 3712 8732
rect 3736 8730 3792 8732
rect 3816 8730 3872 8732
rect 3896 8730 3952 8732
rect 3976 8730 4032 8732
rect 3656 8678 3658 8730
rect 3658 8678 3710 8730
rect 3710 8678 3712 8730
rect 3736 8678 3774 8730
rect 3774 8678 3786 8730
rect 3786 8678 3792 8730
rect 3816 8678 3838 8730
rect 3838 8678 3850 8730
rect 3850 8678 3872 8730
rect 3896 8678 3902 8730
rect 3902 8678 3914 8730
rect 3914 8678 3952 8730
rect 3976 8678 3978 8730
rect 3978 8678 4030 8730
rect 4030 8678 4032 8730
rect 3656 8676 3712 8678
rect 3736 8676 3792 8678
rect 3816 8676 3872 8678
rect 3896 8676 3952 8678
rect 3976 8676 4032 8678
rect 10916 9274 10972 9276
rect 10996 9274 11052 9276
rect 11076 9274 11132 9276
rect 11156 9274 11212 9276
rect 11236 9274 11292 9276
rect 10916 9222 10918 9274
rect 10918 9222 10970 9274
rect 10970 9222 10972 9274
rect 10996 9222 11034 9274
rect 11034 9222 11046 9274
rect 11046 9222 11052 9274
rect 11076 9222 11098 9274
rect 11098 9222 11110 9274
rect 11110 9222 11132 9274
rect 11156 9222 11162 9274
rect 11162 9222 11174 9274
rect 11174 9222 11212 9274
rect 11236 9222 11238 9274
rect 11238 9222 11290 9274
rect 11290 9222 11292 9274
rect 10916 9220 10972 9222
rect 10996 9220 11052 9222
rect 11076 9220 11132 9222
rect 11156 9220 11212 9222
rect 11236 9220 11292 9222
rect 1398 8336 1454 8392
rect 2916 8186 2972 8188
rect 2996 8186 3052 8188
rect 3076 8186 3132 8188
rect 3156 8186 3212 8188
rect 3236 8186 3292 8188
rect 2916 8134 2918 8186
rect 2918 8134 2970 8186
rect 2970 8134 2972 8186
rect 2996 8134 3034 8186
rect 3034 8134 3046 8186
rect 3046 8134 3052 8186
rect 3076 8134 3098 8186
rect 3098 8134 3110 8186
rect 3110 8134 3132 8186
rect 3156 8134 3162 8186
rect 3162 8134 3174 8186
rect 3174 8134 3212 8186
rect 3236 8134 3238 8186
rect 3238 8134 3290 8186
rect 3290 8134 3292 8186
rect 2916 8132 2972 8134
rect 2996 8132 3052 8134
rect 3076 8132 3132 8134
rect 3156 8132 3212 8134
rect 3236 8132 3292 8134
rect 10916 8186 10972 8188
rect 10996 8186 11052 8188
rect 11076 8186 11132 8188
rect 11156 8186 11212 8188
rect 11236 8186 11292 8188
rect 10916 8134 10918 8186
rect 10918 8134 10970 8186
rect 10970 8134 10972 8186
rect 10996 8134 11034 8186
rect 11034 8134 11046 8186
rect 11046 8134 11052 8186
rect 11076 8134 11098 8186
rect 11098 8134 11110 8186
rect 11110 8134 11132 8186
rect 11156 8134 11162 8186
rect 11162 8134 11174 8186
rect 11174 8134 11212 8186
rect 11236 8134 11238 8186
rect 11238 8134 11290 8186
rect 11290 8134 11292 8186
rect 10916 8132 10972 8134
rect 10996 8132 11052 8134
rect 11076 8132 11132 8134
rect 11156 8132 11212 8134
rect 11236 8132 11292 8134
rect 3656 7642 3712 7644
rect 3736 7642 3792 7644
rect 3816 7642 3872 7644
rect 3896 7642 3952 7644
rect 3976 7642 4032 7644
rect 3656 7590 3658 7642
rect 3658 7590 3710 7642
rect 3710 7590 3712 7642
rect 3736 7590 3774 7642
rect 3774 7590 3786 7642
rect 3786 7590 3792 7642
rect 3816 7590 3838 7642
rect 3838 7590 3850 7642
rect 3850 7590 3872 7642
rect 3896 7590 3902 7642
rect 3902 7590 3914 7642
rect 3914 7590 3952 7642
rect 3976 7590 3978 7642
rect 3978 7590 4030 7642
rect 4030 7590 4032 7642
rect 3656 7588 3712 7590
rect 3736 7588 3792 7590
rect 3816 7588 3872 7590
rect 3896 7588 3952 7590
rect 3976 7588 4032 7590
rect 1398 7520 1454 7576
rect 2916 7098 2972 7100
rect 2996 7098 3052 7100
rect 3076 7098 3132 7100
rect 3156 7098 3212 7100
rect 3236 7098 3292 7100
rect 2916 7046 2918 7098
rect 2918 7046 2970 7098
rect 2970 7046 2972 7098
rect 2996 7046 3034 7098
rect 3034 7046 3046 7098
rect 3046 7046 3052 7098
rect 3076 7046 3098 7098
rect 3098 7046 3110 7098
rect 3110 7046 3132 7098
rect 3156 7046 3162 7098
rect 3162 7046 3174 7098
rect 3174 7046 3212 7098
rect 3236 7046 3238 7098
rect 3238 7046 3290 7098
rect 3290 7046 3292 7098
rect 2916 7044 2972 7046
rect 2996 7044 3052 7046
rect 3076 7044 3132 7046
rect 3156 7044 3212 7046
rect 3236 7044 3292 7046
rect 3656 6554 3712 6556
rect 3736 6554 3792 6556
rect 3816 6554 3872 6556
rect 3896 6554 3952 6556
rect 3976 6554 4032 6556
rect 3656 6502 3658 6554
rect 3658 6502 3710 6554
rect 3710 6502 3712 6554
rect 3736 6502 3774 6554
rect 3774 6502 3786 6554
rect 3786 6502 3792 6554
rect 3816 6502 3838 6554
rect 3838 6502 3850 6554
rect 3850 6502 3872 6554
rect 3896 6502 3902 6554
rect 3902 6502 3914 6554
rect 3914 6502 3952 6554
rect 3976 6502 3978 6554
rect 3978 6502 4030 6554
rect 4030 6502 4032 6554
rect 3656 6500 3712 6502
rect 3736 6500 3792 6502
rect 3816 6500 3872 6502
rect 3896 6500 3952 6502
rect 3976 6500 4032 6502
rect 1398 6432 1454 6488
rect 11656 10906 11712 10908
rect 11736 10906 11792 10908
rect 11816 10906 11872 10908
rect 11896 10906 11952 10908
rect 11976 10906 12032 10908
rect 11656 10854 11658 10906
rect 11658 10854 11710 10906
rect 11710 10854 11712 10906
rect 11736 10854 11774 10906
rect 11774 10854 11786 10906
rect 11786 10854 11792 10906
rect 11816 10854 11838 10906
rect 11838 10854 11850 10906
rect 11850 10854 11872 10906
rect 11896 10854 11902 10906
rect 11902 10854 11914 10906
rect 11914 10854 11952 10906
rect 11976 10854 11978 10906
rect 11978 10854 12030 10906
rect 12030 10854 12032 10906
rect 11656 10852 11712 10854
rect 11736 10852 11792 10854
rect 11816 10852 11872 10854
rect 11896 10852 11952 10854
rect 11976 10852 12032 10854
rect 11518 10376 11574 10432
rect 10916 7098 10972 7100
rect 10996 7098 11052 7100
rect 11076 7098 11132 7100
rect 11156 7098 11212 7100
rect 11236 7098 11292 7100
rect 10916 7046 10918 7098
rect 10918 7046 10970 7098
rect 10970 7046 10972 7098
rect 10996 7046 11034 7098
rect 11034 7046 11046 7098
rect 11046 7046 11052 7098
rect 11076 7046 11098 7098
rect 11098 7046 11110 7098
rect 11110 7046 11132 7098
rect 11156 7046 11162 7098
rect 11162 7046 11174 7098
rect 11174 7046 11212 7098
rect 11236 7046 11238 7098
rect 11238 7046 11290 7098
rect 11290 7046 11292 7098
rect 10916 7044 10972 7046
rect 10996 7044 11052 7046
rect 11076 7044 11132 7046
rect 11156 7044 11212 7046
rect 11236 7044 11292 7046
rect 2916 6010 2972 6012
rect 2996 6010 3052 6012
rect 3076 6010 3132 6012
rect 3156 6010 3212 6012
rect 3236 6010 3292 6012
rect 2916 5958 2918 6010
rect 2918 5958 2970 6010
rect 2970 5958 2972 6010
rect 2996 5958 3034 6010
rect 3034 5958 3046 6010
rect 3046 5958 3052 6010
rect 3076 5958 3098 6010
rect 3098 5958 3110 6010
rect 3110 5958 3132 6010
rect 3156 5958 3162 6010
rect 3162 5958 3174 6010
rect 3174 5958 3212 6010
rect 3236 5958 3238 6010
rect 3238 5958 3290 6010
rect 3290 5958 3292 6010
rect 2916 5956 2972 5958
rect 2996 5956 3052 5958
rect 3076 5956 3132 5958
rect 3156 5956 3212 5958
rect 3236 5956 3292 5958
rect 1398 5888 1454 5944
rect 3656 5466 3712 5468
rect 3736 5466 3792 5468
rect 3816 5466 3872 5468
rect 3896 5466 3952 5468
rect 3976 5466 4032 5468
rect 3656 5414 3658 5466
rect 3658 5414 3710 5466
rect 3710 5414 3712 5466
rect 3736 5414 3774 5466
rect 3774 5414 3786 5466
rect 3786 5414 3792 5466
rect 3816 5414 3838 5466
rect 3838 5414 3850 5466
rect 3850 5414 3872 5466
rect 3896 5414 3902 5466
rect 3902 5414 3914 5466
rect 3914 5414 3952 5466
rect 3976 5414 3978 5466
rect 3978 5414 4030 5466
rect 4030 5414 4032 5466
rect 3656 5412 3712 5414
rect 3736 5412 3792 5414
rect 3816 5412 3872 5414
rect 3896 5412 3952 5414
rect 3976 5412 4032 5414
rect 1398 5228 1454 5264
rect 1398 5208 1400 5228
rect 1400 5208 1452 5228
rect 1452 5208 1454 5228
rect 2916 4922 2972 4924
rect 2996 4922 3052 4924
rect 3076 4922 3132 4924
rect 3156 4922 3212 4924
rect 3236 4922 3292 4924
rect 2916 4870 2918 4922
rect 2918 4870 2970 4922
rect 2970 4870 2972 4922
rect 2996 4870 3034 4922
rect 3034 4870 3046 4922
rect 3046 4870 3052 4922
rect 3076 4870 3098 4922
rect 3098 4870 3110 4922
rect 3110 4870 3132 4922
rect 3156 4870 3162 4922
rect 3162 4870 3174 4922
rect 3174 4870 3212 4922
rect 3236 4870 3238 4922
rect 3238 4870 3290 4922
rect 3290 4870 3292 4922
rect 2916 4868 2972 4870
rect 2996 4868 3052 4870
rect 3076 4868 3132 4870
rect 3156 4868 3212 4870
rect 3236 4868 3292 4870
rect 10916 6010 10972 6012
rect 10996 6010 11052 6012
rect 11076 6010 11132 6012
rect 11156 6010 11212 6012
rect 11236 6010 11292 6012
rect 10916 5958 10918 6010
rect 10918 5958 10970 6010
rect 10970 5958 10972 6010
rect 10996 5958 11034 6010
rect 11034 5958 11046 6010
rect 11046 5958 11052 6010
rect 11076 5958 11098 6010
rect 11098 5958 11110 6010
rect 11110 5958 11132 6010
rect 11156 5958 11162 6010
rect 11162 5958 11174 6010
rect 11174 5958 11212 6010
rect 11236 5958 11238 6010
rect 11238 5958 11290 6010
rect 11290 5958 11292 6010
rect 10916 5956 10972 5958
rect 10996 5956 11052 5958
rect 11076 5956 11132 5958
rect 11156 5956 11212 5958
rect 11236 5956 11292 5958
rect 3656 4378 3712 4380
rect 3736 4378 3792 4380
rect 3816 4378 3872 4380
rect 3896 4378 3952 4380
rect 3976 4378 4032 4380
rect 3656 4326 3658 4378
rect 3658 4326 3710 4378
rect 3710 4326 3712 4378
rect 3736 4326 3774 4378
rect 3774 4326 3786 4378
rect 3786 4326 3792 4378
rect 3816 4326 3838 4378
rect 3838 4326 3850 4378
rect 3850 4326 3872 4378
rect 3896 4326 3902 4378
rect 3902 4326 3914 4378
rect 3914 4326 3952 4378
rect 3976 4326 3978 4378
rect 3978 4326 4030 4378
rect 4030 4326 4032 4378
rect 3656 4324 3712 4326
rect 3736 4324 3792 4326
rect 3816 4324 3872 4326
rect 3896 4324 3952 4326
rect 3976 4324 4032 4326
rect 1398 4256 1454 4312
rect 2916 3834 2972 3836
rect 2996 3834 3052 3836
rect 3076 3834 3132 3836
rect 3156 3834 3212 3836
rect 3236 3834 3292 3836
rect 2916 3782 2918 3834
rect 2918 3782 2970 3834
rect 2970 3782 2972 3834
rect 2996 3782 3034 3834
rect 3034 3782 3046 3834
rect 3046 3782 3052 3834
rect 3076 3782 3098 3834
rect 3098 3782 3110 3834
rect 3110 3782 3132 3834
rect 3156 3782 3162 3834
rect 3162 3782 3174 3834
rect 3174 3782 3212 3834
rect 3236 3782 3238 3834
rect 3238 3782 3290 3834
rect 3290 3782 3292 3834
rect 2916 3780 2972 3782
rect 2996 3780 3052 3782
rect 3076 3780 3132 3782
rect 3156 3780 3212 3782
rect 3236 3780 3292 3782
rect 10916 4922 10972 4924
rect 10996 4922 11052 4924
rect 11076 4922 11132 4924
rect 11156 4922 11212 4924
rect 11236 4922 11292 4924
rect 10916 4870 10918 4922
rect 10918 4870 10970 4922
rect 10970 4870 10972 4922
rect 10996 4870 11034 4922
rect 11034 4870 11046 4922
rect 11046 4870 11052 4922
rect 11076 4870 11098 4922
rect 11098 4870 11110 4922
rect 11110 4870 11132 4922
rect 11156 4870 11162 4922
rect 11162 4870 11174 4922
rect 11174 4870 11212 4922
rect 11236 4870 11238 4922
rect 11238 4870 11290 4922
rect 11290 4870 11292 4922
rect 10916 4868 10972 4870
rect 10996 4868 11052 4870
rect 11076 4868 11132 4870
rect 11156 4868 11212 4870
rect 11236 4868 11292 4870
rect 11656 9818 11712 9820
rect 11736 9818 11792 9820
rect 11816 9818 11872 9820
rect 11896 9818 11952 9820
rect 11976 9818 12032 9820
rect 11656 9766 11658 9818
rect 11658 9766 11710 9818
rect 11710 9766 11712 9818
rect 11736 9766 11774 9818
rect 11774 9766 11786 9818
rect 11786 9766 11792 9818
rect 11816 9766 11838 9818
rect 11838 9766 11850 9818
rect 11850 9766 11872 9818
rect 11896 9766 11902 9818
rect 11902 9766 11914 9818
rect 11914 9766 11952 9818
rect 11976 9766 11978 9818
rect 11978 9766 12030 9818
rect 12030 9766 12032 9818
rect 11656 9764 11712 9766
rect 11736 9764 11792 9766
rect 11816 9764 11872 9766
rect 11896 9764 11952 9766
rect 11976 9764 12032 9766
rect 11656 8730 11712 8732
rect 11736 8730 11792 8732
rect 11816 8730 11872 8732
rect 11896 8730 11952 8732
rect 11976 8730 12032 8732
rect 11656 8678 11658 8730
rect 11658 8678 11710 8730
rect 11710 8678 11712 8730
rect 11736 8678 11774 8730
rect 11774 8678 11786 8730
rect 11786 8678 11792 8730
rect 11816 8678 11838 8730
rect 11838 8678 11850 8730
rect 11850 8678 11872 8730
rect 11896 8678 11902 8730
rect 11902 8678 11914 8730
rect 11914 8678 11952 8730
rect 11976 8678 11978 8730
rect 11978 8678 12030 8730
rect 12030 8678 12032 8730
rect 11656 8676 11712 8678
rect 11736 8676 11792 8678
rect 11816 8676 11872 8678
rect 11896 8676 11952 8678
rect 11976 8676 12032 8678
rect 11656 7642 11712 7644
rect 11736 7642 11792 7644
rect 11816 7642 11872 7644
rect 11896 7642 11952 7644
rect 11976 7642 12032 7644
rect 11656 7590 11658 7642
rect 11658 7590 11710 7642
rect 11710 7590 11712 7642
rect 11736 7590 11774 7642
rect 11774 7590 11786 7642
rect 11786 7590 11792 7642
rect 11816 7590 11838 7642
rect 11838 7590 11850 7642
rect 11850 7590 11872 7642
rect 11896 7590 11902 7642
rect 11902 7590 11914 7642
rect 11914 7590 11952 7642
rect 11976 7590 11978 7642
rect 11978 7590 12030 7642
rect 12030 7590 12032 7642
rect 11656 7588 11712 7590
rect 11736 7588 11792 7590
rect 11816 7588 11872 7590
rect 11896 7588 11952 7590
rect 11976 7588 12032 7590
rect 11656 6554 11712 6556
rect 11736 6554 11792 6556
rect 11816 6554 11872 6556
rect 11896 6554 11952 6556
rect 11976 6554 12032 6556
rect 11656 6502 11658 6554
rect 11658 6502 11710 6554
rect 11710 6502 11712 6554
rect 11736 6502 11774 6554
rect 11774 6502 11786 6554
rect 11786 6502 11792 6554
rect 11816 6502 11838 6554
rect 11838 6502 11850 6554
rect 11850 6502 11872 6554
rect 11896 6502 11902 6554
rect 11902 6502 11914 6554
rect 11914 6502 11952 6554
rect 11976 6502 11978 6554
rect 11978 6502 12030 6554
rect 12030 6502 12032 6554
rect 11656 6500 11712 6502
rect 11736 6500 11792 6502
rect 11816 6500 11872 6502
rect 11896 6500 11952 6502
rect 11976 6500 12032 6502
rect 11656 5466 11712 5468
rect 11736 5466 11792 5468
rect 11816 5466 11872 5468
rect 11896 5466 11952 5468
rect 11976 5466 12032 5468
rect 11656 5414 11658 5466
rect 11658 5414 11710 5466
rect 11710 5414 11712 5466
rect 11736 5414 11774 5466
rect 11774 5414 11786 5466
rect 11786 5414 11792 5466
rect 11816 5414 11838 5466
rect 11838 5414 11850 5466
rect 11850 5414 11872 5466
rect 11896 5414 11902 5466
rect 11902 5414 11914 5466
rect 11914 5414 11952 5466
rect 11976 5414 11978 5466
rect 11978 5414 12030 5466
rect 12030 5414 12032 5466
rect 11656 5412 11712 5414
rect 11736 5412 11792 5414
rect 11816 5412 11872 5414
rect 11896 5412 11952 5414
rect 11976 5412 12032 5414
rect 11656 4378 11712 4380
rect 11736 4378 11792 4380
rect 11816 4378 11872 4380
rect 11896 4378 11952 4380
rect 11976 4378 12032 4380
rect 11656 4326 11658 4378
rect 11658 4326 11710 4378
rect 11710 4326 11712 4378
rect 11736 4326 11774 4378
rect 11774 4326 11786 4378
rect 11786 4326 11792 4378
rect 11816 4326 11838 4378
rect 11838 4326 11850 4378
rect 11850 4326 11872 4378
rect 11896 4326 11902 4378
rect 11902 4326 11914 4378
rect 11914 4326 11952 4378
rect 11976 4326 11978 4378
rect 11978 4326 12030 4378
rect 12030 4326 12032 4378
rect 11656 4324 11712 4326
rect 11736 4324 11792 4326
rect 11816 4324 11872 4326
rect 11896 4324 11952 4326
rect 11976 4324 12032 4326
rect 10916 3834 10972 3836
rect 10996 3834 11052 3836
rect 11076 3834 11132 3836
rect 11156 3834 11212 3836
rect 11236 3834 11292 3836
rect 10916 3782 10918 3834
rect 10918 3782 10970 3834
rect 10970 3782 10972 3834
rect 10996 3782 11034 3834
rect 11034 3782 11046 3834
rect 11046 3782 11052 3834
rect 11076 3782 11098 3834
rect 11098 3782 11110 3834
rect 11110 3782 11132 3834
rect 11156 3782 11162 3834
rect 11162 3782 11174 3834
rect 11174 3782 11212 3834
rect 11236 3782 11238 3834
rect 11238 3782 11290 3834
rect 11290 3782 11292 3834
rect 10916 3780 10972 3782
rect 10996 3780 11052 3782
rect 11076 3780 11132 3782
rect 11156 3780 11212 3782
rect 11236 3780 11292 3782
rect 1398 3476 1400 3496
rect 1400 3476 1452 3496
rect 1452 3476 1454 3496
rect 1398 3440 1454 3476
rect 3656 3290 3712 3292
rect 3736 3290 3792 3292
rect 3816 3290 3872 3292
rect 3896 3290 3952 3292
rect 3976 3290 4032 3292
rect 3656 3238 3658 3290
rect 3658 3238 3710 3290
rect 3710 3238 3712 3290
rect 3736 3238 3774 3290
rect 3774 3238 3786 3290
rect 3786 3238 3792 3290
rect 3816 3238 3838 3290
rect 3838 3238 3850 3290
rect 3850 3238 3872 3290
rect 3896 3238 3902 3290
rect 3902 3238 3914 3290
rect 3914 3238 3952 3290
rect 3976 3238 3978 3290
rect 3978 3238 4030 3290
rect 4030 3238 4032 3290
rect 3656 3236 3712 3238
rect 3736 3236 3792 3238
rect 3816 3236 3872 3238
rect 3896 3236 3952 3238
rect 3976 3236 4032 3238
rect 18916 14714 18972 14716
rect 18996 14714 19052 14716
rect 19076 14714 19132 14716
rect 19156 14714 19212 14716
rect 19236 14714 19292 14716
rect 18916 14662 18918 14714
rect 18918 14662 18970 14714
rect 18970 14662 18972 14714
rect 18996 14662 19034 14714
rect 19034 14662 19046 14714
rect 19046 14662 19052 14714
rect 19076 14662 19098 14714
rect 19098 14662 19110 14714
rect 19110 14662 19132 14714
rect 19156 14662 19162 14714
rect 19162 14662 19174 14714
rect 19174 14662 19212 14714
rect 19236 14662 19238 14714
rect 19238 14662 19290 14714
rect 19290 14662 19292 14714
rect 18916 14660 18972 14662
rect 18996 14660 19052 14662
rect 19076 14660 19132 14662
rect 19156 14660 19212 14662
rect 19236 14660 19292 14662
rect 26916 14714 26972 14716
rect 26996 14714 27052 14716
rect 27076 14714 27132 14716
rect 27156 14714 27212 14716
rect 27236 14714 27292 14716
rect 26916 14662 26918 14714
rect 26918 14662 26970 14714
rect 26970 14662 26972 14714
rect 26996 14662 27034 14714
rect 27034 14662 27046 14714
rect 27046 14662 27052 14714
rect 27076 14662 27098 14714
rect 27098 14662 27110 14714
rect 27110 14662 27132 14714
rect 27156 14662 27162 14714
rect 27162 14662 27174 14714
rect 27174 14662 27212 14714
rect 27236 14662 27238 14714
rect 27238 14662 27290 14714
rect 27290 14662 27292 14714
rect 26916 14660 26972 14662
rect 26996 14660 27052 14662
rect 27076 14660 27132 14662
rect 27156 14660 27212 14662
rect 27236 14660 27292 14662
rect 28354 14456 28410 14512
rect 19656 14170 19712 14172
rect 19736 14170 19792 14172
rect 19816 14170 19872 14172
rect 19896 14170 19952 14172
rect 19976 14170 20032 14172
rect 19656 14118 19658 14170
rect 19658 14118 19710 14170
rect 19710 14118 19712 14170
rect 19736 14118 19774 14170
rect 19774 14118 19786 14170
rect 19786 14118 19792 14170
rect 19816 14118 19838 14170
rect 19838 14118 19850 14170
rect 19850 14118 19872 14170
rect 19896 14118 19902 14170
rect 19902 14118 19914 14170
rect 19914 14118 19952 14170
rect 19976 14118 19978 14170
rect 19978 14118 20030 14170
rect 20030 14118 20032 14170
rect 19656 14116 19712 14118
rect 19736 14116 19792 14118
rect 19816 14116 19872 14118
rect 19896 14116 19952 14118
rect 19976 14116 20032 14118
rect 27656 14170 27712 14172
rect 27736 14170 27792 14172
rect 27816 14170 27872 14172
rect 27896 14170 27952 14172
rect 27976 14170 28032 14172
rect 27656 14118 27658 14170
rect 27658 14118 27710 14170
rect 27710 14118 27712 14170
rect 27736 14118 27774 14170
rect 27774 14118 27786 14170
rect 27786 14118 27792 14170
rect 27816 14118 27838 14170
rect 27838 14118 27850 14170
rect 27850 14118 27872 14170
rect 27896 14118 27902 14170
rect 27902 14118 27914 14170
rect 27914 14118 27952 14170
rect 27976 14118 27978 14170
rect 27978 14118 28030 14170
rect 28030 14118 28032 14170
rect 27656 14116 27712 14118
rect 27736 14116 27792 14118
rect 27816 14116 27872 14118
rect 27896 14116 27952 14118
rect 27976 14116 28032 14118
rect 28354 13640 28410 13696
rect 18916 13626 18972 13628
rect 18996 13626 19052 13628
rect 19076 13626 19132 13628
rect 19156 13626 19212 13628
rect 19236 13626 19292 13628
rect 18916 13574 18918 13626
rect 18918 13574 18970 13626
rect 18970 13574 18972 13626
rect 18996 13574 19034 13626
rect 19034 13574 19046 13626
rect 19046 13574 19052 13626
rect 19076 13574 19098 13626
rect 19098 13574 19110 13626
rect 19110 13574 19132 13626
rect 19156 13574 19162 13626
rect 19162 13574 19174 13626
rect 19174 13574 19212 13626
rect 19236 13574 19238 13626
rect 19238 13574 19290 13626
rect 19290 13574 19292 13626
rect 18916 13572 18972 13574
rect 18996 13572 19052 13574
rect 19076 13572 19132 13574
rect 19156 13572 19212 13574
rect 19236 13572 19292 13574
rect 26916 13626 26972 13628
rect 26996 13626 27052 13628
rect 27076 13626 27132 13628
rect 27156 13626 27212 13628
rect 27236 13626 27292 13628
rect 26916 13574 26918 13626
rect 26918 13574 26970 13626
rect 26970 13574 26972 13626
rect 26996 13574 27034 13626
rect 27034 13574 27046 13626
rect 27046 13574 27052 13626
rect 27076 13574 27098 13626
rect 27098 13574 27110 13626
rect 27110 13574 27132 13626
rect 27156 13574 27162 13626
rect 27162 13574 27174 13626
rect 27174 13574 27212 13626
rect 27236 13574 27238 13626
rect 27238 13574 27290 13626
rect 27290 13574 27292 13626
rect 26916 13572 26972 13574
rect 26996 13572 27052 13574
rect 27076 13572 27132 13574
rect 27156 13572 27212 13574
rect 27236 13572 27292 13574
rect 19656 13082 19712 13084
rect 19736 13082 19792 13084
rect 19816 13082 19872 13084
rect 19896 13082 19952 13084
rect 19976 13082 20032 13084
rect 19656 13030 19658 13082
rect 19658 13030 19710 13082
rect 19710 13030 19712 13082
rect 19736 13030 19774 13082
rect 19774 13030 19786 13082
rect 19786 13030 19792 13082
rect 19816 13030 19838 13082
rect 19838 13030 19850 13082
rect 19850 13030 19872 13082
rect 19896 13030 19902 13082
rect 19902 13030 19914 13082
rect 19914 13030 19952 13082
rect 19976 13030 19978 13082
rect 19978 13030 20030 13082
rect 20030 13030 20032 13082
rect 19656 13028 19712 13030
rect 19736 13028 19792 13030
rect 19816 13028 19872 13030
rect 19896 13028 19952 13030
rect 19976 13028 20032 13030
rect 27656 13082 27712 13084
rect 27736 13082 27792 13084
rect 27816 13082 27872 13084
rect 27896 13082 27952 13084
rect 27976 13082 28032 13084
rect 27656 13030 27658 13082
rect 27658 13030 27710 13082
rect 27710 13030 27712 13082
rect 27736 13030 27774 13082
rect 27774 13030 27786 13082
rect 27786 13030 27792 13082
rect 27816 13030 27838 13082
rect 27838 13030 27850 13082
rect 27850 13030 27872 13082
rect 27896 13030 27902 13082
rect 27902 13030 27914 13082
rect 27914 13030 27952 13082
rect 27976 13030 27978 13082
rect 27978 13030 28030 13082
rect 28030 13030 28032 13082
rect 27656 13028 27712 13030
rect 27736 13028 27792 13030
rect 27816 13028 27872 13030
rect 27896 13028 27952 13030
rect 27976 13028 28032 13030
rect 28354 12824 28410 12880
rect 18916 12538 18972 12540
rect 18996 12538 19052 12540
rect 19076 12538 19132 12540
rect 19156 12538 19212 12540
rect 19236 12538 19292 12540
rect 18916 12486 18918 12538
rect 18918 12486 18970 12538
rect 18970 12486 18972 12538
rect 18996 12486 19034 12538
rect 19034 12486 19046 12538
rect 19046 12486 19052 12538
rect 19076 12486 19098 12538
rect 19098 12486 19110 12538
rect 19110 12486 19132 12538
rect 19156 12486 19162 12538
rect 19162 12486 19174 12538
rect 19174 12486 19212 12538
rect 19236 12486 19238 12538
rect 19238 12486 19290 12538
rect 19290 12486 19292 12538
rect 18916 12484 18972 12486
rect 18996 12484 19052 12486
rect 19076 12484 19132 12486
rect 19156 12484 19212 12486
rect 19236 12484 19292 12486
rect 26916 12538 26972 12540
rect 26996 12538 27052 12540
rect 27076 12538 27132 12540
rect 27156 12538 27212 12540
rect 27236 12538 27292 12540
rect 26916 12486 26918 12538
rect 26918 12486 26970 12538
rect 26970 12486 26972 12538
rect 26996 12486 27034 12538
rect 27034 12486 27046 12538
rect 27046 12486 27052 12538
rect 27076 12486 27098 12538
rect 27098 12486 27110 12538
rect 27110 12486 27132 12538
rect 27156 12486 27162 12538
rect 27162 12486 27174 12538
rect 27174 12486 27212 12538
rect 27236 12486 27238 12538
rect 27238 12486 27290 12538
rect 27290 12486 27292 12538
rect 26916 12484 26972 12486
rect 26996 12484 27052 12486
rect 27076 12484 27132 12486
rect 27156 12484 27212 12486
rect 27236 12484 27292 12486
rect 28354 12008 28410 12064
rect 19656 11994 19712 11996
rect 19736 11994 19792 11996
rect 19816 11994 19872 11996
rect 19896 11994 19952 11996
rect 19976 11994 20032 11996
rect 19656 11942 19658 11994
rect 19658 11942 19710 11994
rect 19710 11942 19712 11994
rect 19736 11942 19774 11994
rect 19774 11942 19786 11994
rect 19786 11942 19792 11994
rect 19816 11942 19838 11994
rect 19838 11942 19850 11994
rect 19850 11942 19872 11994
rect 19896 11942 19902 11994
rect 19902 11942 19914 11994
rect 19914 11942 19952 11994
rect 19976 11942 19978 11994
rect 19978 11942 20030 11994
rect 20030 11942 20032 11994
rect 19656 11940 19712 11942
rect 19736 11940 19792 11942
rect 19816 11940 19872 11942
rect 19896 11940 19952 11942
rect 19976 11940 20032 11942
rect 27656 11994 27712 11996
rect 27736 11994 27792 11996
rect 27816 11994 27872 11996
rect 27896 11994 27952 11996
rect 27976 11994 28032 11996
rect 27656 11942 27658 11994
rect 27658 11942 27710 11994
rect 27710 11942 27712 11994
rect 27736 11942 27774 11994
rect 27774 11942 27786 11994
rect 27786 11942 27792 11994
rect 27816 11942 27838 11994
rect 27838 11942 27850 11994
rect 27850 11942 27872 11994
rect 27896 11942 27902 11994
rect 27902 11942 27914 11994
rect 27914 11942 27952 11994
rect 27976 11942 27978 11994
rect 27978 11942 28030 11994
rect 28030 11942 28032 11994
rect 27656 11940 27712 11942
rect 27736 11940 27792 11942
rect 27816 11940 27872 11942
rect 27896 11940 27952 11942
rect 27976 11940 28032 11942
rect 18916 11450 18972 11452
rect 18996 11450 19052 11452
rect 19076 11450 19132 11452
rect 19156 11450 19212 11452
rect 19236 11450 19292 11452
rect 18916 11398 18918 11450
rect 18918 11398 18970 11450
rect 18970 11398 18972 11450
rect 18996 11398 19034 11450
rect 19034 11398 19046 11450
rect 19046 11398 19052 11450
rect 19076 11398 19098 11450
rect 19098 11398 19110 11450
rect 19110 11398 19132 11450
rect 19156 11398 19162 11450
rect 19162 11398 19174 11450
rect 19174 11398 19212 11450
rect 19236 11398 19238 11450
rect 19238 11398 19290 11450
rect 19290 11398 19292 11450
rect 18916 11396 18972 11398
rect 18996 11396 19052 11398
rect 19076 11396 19132 11398
rect 19156 11396 19212 11398
rect 19236 11396 19292 11398
rect 26916 11450 26972 11452
rect 26996 11450 27052 11452
rect 27076 11450 27132 11452
rect 27156 11450 27212 11452
rect 27236 11450 27292 11452
rect 26916 11398 26918 11450
rect 26918 11398 26970 11450
rect 26970 11398 26972 11450
rect 26996 11398 27034 11450
rect 27034 11398 27046 11450
rect 27046 11398 27052 11450
rect 27076 11398 27098 11450
rect 27098 11398 27110 11450
rect 27110 11398 27132 11450
rect 27156 11398 27162 11450
rect 27162 11398 27174 11450
rect 27174 11398 27212 11450
rect 27236 11398 27238 11450
rect 27238 11398 27290 11450
rect 27290 11398 27292 11450
rect 26916 11396 26972 11398
rect 26996 11396 27052 11398
rect 27076 11396 27132 11398
rect 27156 11396 27212 11398
rect 27236 11396 27292 11398
rect 28354 11192 28410 11248
rect 19656 10906 19712 10908
rect 19736 10906 19792 10908
rect 19816 10906 19872 10908
rect 19896 10906 19952 10908
rect 19976 10906 20032 10908
rect 19656 10854 19658 10906
rect 19658 10854 19710 10906
rect 19710 10854 19712 10906
rect 19736 10854 19774 10906
rect 19774 10854 19786 10906
rect 19786 10854 19792 10906
rect 19816 10854 19838 10906
rect 19838 10854 19850 10906
rect 19850 10854 19872 10906
rect 19896 10854 19902 10906
rect 19902 10854 19914 10906
rect 19914 10854 19952 10906
rect 19976 10854 19978 10906
rect 19978 10854 20030 10906
rect 20030 10854 20032 10906
rect 19656 10852 19712 10854
rect 19736 10852 19792 10854
rect 19816 10852 19872 10854
rect 19896 10852 19952 10854
rect 19976 10852 20032 10854
rect 27656 10906 27712 10908
rect 27736 10906 27792 10908
rect 27816 10906 27872 10908
rect 27896 10906 27952 10908
rect 27976 10906 28032 10908
rect 27656 10854 27658 10906
rect 27658 10854 27710 10906
rect 27710 10854 27712 10906
rect 27736 10854 27774 10906
rect 27774 10854 27786 10906
rect 27786 10854 27792 10906
rect 27816 10854 27838 10906
rect 27838 10854 27850 10906
rect 27850 10854 27872 10906
rect 27896 10854 27902 10906
rect 27902 10854 27914 10906
rect 27914 10854 27952 10906
rect 27976 10854 27978 10906
rect 27978 10854 28030 10906
rect 28030 10854 28032 10906
rect 27656 10852 27712 10854
rect 27736 10852 27792 10854
rect 27816 10852 27872 10854
rect 27896 10852 27952 10854
rect 27976 10852 28032 10854
rect 28354 10376 28410 10432
rect 18916 10362 18972 10364
rect 18996 10362 19052 10364
rect 19076 10362 19132 10364
rect 19156 10362 19212 10364
rect 19236 10362 19292 10364
rect 18916 10310 18918 10362
rect 18918 10310 18970 10362
rect 18970 10310 18972 10362
rect 18996 10310 19034 10362
rect 19034 10310 19046 10362
rect 19046 10310 19052 10362
rect 19076 10310 19098 10362
rect 19098 10310 19110 10362
rect 19110 10310 19132 10362
rect 19156 10310 19162 10362
rect 19162 10310 19174 10362
rect 19174 10310 19212 10362
rect 19236 10310 19238 10362
rect 19238 10310 19290 10362
rect 19290 10310 19292 10362
rect 18916 10308 18972 10310
rect 18996 10308 19052 10310
rect 19076 10308 19132 10310
rect 19156 10308 19212 10310
rect 19236 10308 19292 10310
rect 26916 10362 26972 10364
rect 26996 10362 27052 10364
rect 27076 10362 27132 10364
rect 27156 10362 27212 10364
rect 27236 10362 27292 10364
rect 26916 10310 26918 10362
rect 26918 10310 26970 10362
rect 26970 10310 26972 10362
rect 26996 10310 27034 10362
rect 27034 10310 27046 10362
rect 27046 10310 27052 10362
rect 27076 10310 27098 10362
rect 27098 10310 27110 10362
rect 27110 10310 27132 10362
rect 27156 10310 27162 10362
rect 27162 10310 27174 10362
rect 27174 10310 27212 10362
rect 27236 10310 27238 10362
rect 27238 10310 27290 10362
rect 27290 10310 27292 10362
rect 26916 10308 26972 10310
rect 26996 10308 27052 10310
rect 27076 10308 27132 10310
rect 27156 10308 27212 10310
rect 27236 10308 27292 10310
rect 19656 9818 19712 9820
rect 19736 9818 19792 9820
rect 19816 9818 19872 9820
rect 19896 9818 19952 9820
rect 19976 9818 20032 9820
rect 19656 9766 19658 9818
rect 19658 9766 19710 9818
rect 19710 9766 19712 9818
rect 19736 9766 19774 9818
rect 19774 9766 19786 9818
rect 19786 9766 19792 9818
rect 19816 9766 19838 9818
rect 19838 9766 19850 9818
rect 19850 9766 19872 9818
rect 19896 9766 19902 9818
rect 19902 9766 19914 9818
rect 19914 9766 19952 9818
rect 19976 9766 19978 9818
rect 19978 9766 20030 9818
rect 20030 9766 20032 9818
rect 19656 9764 19712 9766
rect 19736 9764 19792 9766
rect 19816 9764 19872 9766
rect 19896 9764 19952 9766
rect 19976 9764 20032 9766
rect 27656 9818 27712 9820
rect 27736 9818 27792 9820
rect 27816 9818 27872 9820
rect 27896 9818 27952 9820
rect 27976 9818 28032 9820
rect 27656 9766 27658 9818
rect 27658 9766 27710 9818
rect 27710 9766 27712 9818
rect 27736 9766 27774 9818
rect 27774 9766 27786 9818
rect 27786 9766 27792 9818
rect 27816 9766 27838 9818
rect 27838 9766 27850 9818
rect 27850 9766 27872 9818
rect 27896 9766 27902 9818
rect 27902 9766 27914 9818
rect 27914 9766 27952 9818
rect 27976 9766 27978 9818
rect 27978 9766 28030 9818
rect 28030 9766 28032 9818
rect 27656 9764 27712 9766
rect 27736 9764 27792 9766
rect 27816 9764 27872 9766
rect 27896 9764 27952 9766
rect 27976 9764 28032 9766
rect 28354 9560 28410 9616
rect 18916 9274 18972 9276
rect 18996 9274 19052 9276
rect 19076 9274 19132 9276
rect 19156 9274 19212 9276
rect 19236 9274 19292 9276
rect 18916 9222 18918 9274
rect 18918 9222 18970 9274
rect 18970 9222 18972 9274
rect 18996 9222 19034 9274
rect 19034 9222 19046 9274
rect 19046 9222 19052 9274
rect 19076 9222 19098 9274
rect 19098 9222 19110 9274
rect 19110 9222 19132 9274
rect 19156 9222 19162 9274
rect 19162 9222 19174 9274
rect 19174 9222 19212 9274
rect 19236 9222 19238 9274
rect 19238 9222 19290 9274
rect 19290 9222 19292 9274
rect 18916 9220 18972 9222
rect 18996 9220 19052 9222
rect 19076 9220 19132 9222
rect 19156 9220 19212 9222
rect 19236 9220 19292 9222
rect 26916 9274 26972 9276
rect 26996 9274 27052 9276
rect 27076 9274 27132 9276
rect 27156 9274 27212 9276
rect 27236 9274 27292 9276
rect 26916 9222 26918 9274
rect 26918 9222 26970 9274
rect 26970 9222 26972 9274
rect 26996 9222 27034 9274
rect 27034 9222 27046 9274
rect 27046 9222 27052 9274
rect 27076 9222 27098 9274
rect 27098 9222 27110 9274
rect 27110 9222 27132 9274
rect 27156 9222 27162 9274
rect 27162 9222 27174 9274
rect 27174 9222 27212 9274
rect 27236 9222 27238 9274
rect 27238 9222 27290 9274
rect 27290 9222 27292 9274
rect 26916 9220 26972 9222
rect 26996 9220 27052 9222
rect 27076 9220 27132 9222
rect 27156 9220 27212 9222
rect 27236 9220 27292 9222
rect 28354 8744 28410 8800
rect 19656 8730 19712 8732
rect 19736 8730 19792 8732
rect 19816 8730 19872 8732
rect 19896 8730 19952 8732
rect 19976 8730 20032 8732
rect 19656 8678 19658 8730
rect 19658 8678 19710 8730
rect 19710 8678 19712 8730
rect 19736 8678 19774 8730
rect 19774 8678 19786 8730
rect 19786 8678 19792 8730
rect 19816 8678 19838 8730
rect 19838 8678 19850 8730
rect 19850 8678 19872 8730
rect 19896 8678 19902 8730
rect 19902 8678 19914 8730
rect 19914 8678 19952 8730
rect 19976 8678 19978 8730
rect 19978 8678 20030 8730
rect 20030 8678 20032 8730
rect 19656 8676 19712 8678
rect 19736 8676 19792 8678
rect 19816 8676 19872 8678
rect 19896 8676 19952 8678
rect 19976 8676 20032 8678
rect 27656 8730 27712 8732
rect 27736 8730 27792 8732
rect 27816 8730 27872 8732
rect 27896 8730 27952 8732
rect 27976 8730 28032 8732
rect 27656 8678 27658 8730
rect 27658 8678 27710 8730
rect 27710 8678 27712 8730
rect 27736 8678 27774 8730
rect 27774 8678 27786 8730
rect 27786 8678 27792 8730
rect 27816 8678 27838 8730
rect 27838 8678 27850 8730
rect 27850 8678 27872 8730
rect 27896 8678 27902 8730
rect 27902 8678 27914 8730
rect 27914 8678 27952 8730
rect 27976 8678 27978 8730
rect 27978 8678 28030 8730
rect 28030 8678 28032 8730
rect 27656 8676 27712 8678
rect 27736 8676 27792 8678
rect 27816 8676 27872 8678
rect 27896 8676 27952 8678
rect 27976 8676 28032 8678
rect 18916 8186 18972 8188
rect 18996 8186 19052 8188
rect 19076 8186 19132 8188
rect 19156 8186 19212 8188
rect 19236 8186 19292 8188
rect 18916 8134 18918 8186
rect 18918 8134 18970 8186
rect 18970 8134 18972 8186
rect 18996 8134 19034 8186
rect 19034 8134 19046 8186
rect 19046 8134 19052 8186
rect 19076 8134 19098 8186
rect 19098 8134 19110 8186
rect 19110 8134 19132 8186
rect 19156 8134 19162 8186
rect 19162 8134 19174 8186
rect 19174 8134 19212 8186
rect 19236 8134 19238 8186
rect 19238 8134 19290 8186
rect 19290 8134 19292 8186
rect 18916 8132 18972 8134
rect 18996 8132 19052 8134
rect 19076 8132 19132 8134
rect 19156 8132 19212 8134
rect 19236 8132 19292 8134
rect 26916 8186 26972 8188
rect 26996 8186 27052 8188
rect 27076 8186 27132 8188
rect 27156 8186 27212 8188
rect 27236 8186 27292 8188
rect 26916 8134 26918 8186
rect 26918 8134 26970 8186
rect 26970 8134 26972 8186
rect 26996 8134 27034 8186
rect 27034 8134 27046 8186
rect 27046 8134 27052 8186
rect 27076 8134 27098 8186
rect 27098 8134 27110 8186
rect 27110 8134 27132 8186
rect 27156 8134 27162 8186
rect 27162 8134 27174 8186
rect 27174 8134 27212 8186
rect 27236 8134 27238 8186
rect 27238 8134 27290 8186
rect 27290 8134 27292 8186
rect 26916 8132 26972 8134
rect 26996 8132 27052 8134
rect 27076 8132 27132 8134
rect 27156 8132 27212 8134
rect 27236 8132 27292 8134
rect 28354 7928 28410 7984
rect 19656 7642 19712 7644
rect 19736 7642 19792 7644
rect 19816 7642 19872 7644
rect 19896 7642 19952 7644
rect 19976 7642 20032 7644
rect 19656 7590 19658 7642
rect 19658 7590 19710 7642
rect 19710 7590 19712 7642
rect 19736 7590 19774 7642
rect 19774 7590 19786 7642
rect 19786 7590 19792 7642
rect 19816 7590 19838 7642
rect 19838 7590 19850 7642
rect 19850 7590 19872 7642
rect 19896 7590 19902 7642
rect 19902 7590 19914 7642
rect 19914 7590 19952 7642
rect 19976 7590 19978 7642
rect 19978 7590 20030 7642
rect 20030 7590 20032 7642
rect 19656 7588 19712 7590
rect 19736 7588 19792 7590
rect 19816 7588 19872 7590
rect 19896 7588 19952 7590
rect 19976 7588 20032 7590
rect 27656 7642 27712 7644
rect 27736 7642 27792 7644
rect 27816 7642 27872 7644
rect 27896 7642 27952 7644
rect 27976 7642 28032 7644
rect 27656 7590 27658 7642
rect 27658 7590 27710 7642
rect 27710 7590 27712 7642
rect 27736 7590 27774 7642
rect 27774 7590 27786 7642
rect 27786 7590 27792 7642
rect 27816 7590 27838 7642
rect 27838 7590 27850 7642
rect 27850 7590 27872 7642
rect 27896 7590 27902 7642
rect 27902 7590 27914 7642
rect 27914 7590 27952 7642
rect 27976 7590 27978 7642
rect 27978 7590 28030 7642
rect 28030 7590 28032 7642
rect 27656 7588 27712 7590
rect 27736 7588 27792 7590
rect 27816 7588 27872 7590
rect 27896 7588 27952 7590
rect 27976 7588 28032 7590
rect 28354 7112 28410 7168
rect 18916 7098 18972 7100
rect 18996 7098 19052 7100
rect 19076 7098 19132 7100
rect 19156 7098 19212 7100
rect 19236 7098 19292 7100
rect 18916 7046 18918 7098
rect 18918 7046 18970 7098
rect 18970 7046 18972 7098
rect 18996 7046 19034 7098
rect 19034 7046 19046 7098
rect 19046 7046 19052 7098
rect 19076 7046 19098 7098
rect 19098 7046 19110 7098
rect 19110 7046 19132 7098
rect 19156 7046 19162 7098
rect 19162 7046 19174 7098
rect 19174 7046 19212 7098
rect 19236 7046 19238 7098
rect 19238 7046 19290 7098
rect 19290 7046 19292 7098
rect 18916 7044 18972 7046
rect 18996 7044 19052 7046
rect 19076 7044 19132 7046
rect 19156 7044 19212 7046
rect 19236 7044 19292 7046
rect 26916 7098 26972 7100
rect 26996 7098 27052 7100
rect 27076 7098 27132 7100
rect 27156 7098 27212 7100
rect 27236 7098 27292 7100
rect 26916 7046 26918 7098
rect 26918 7046 26970 7098
rect 26970 7046 26972 7098
rect 26996 7046 27034 7098
rect 27034 7046 27046 7098
rect 27046 7046 27052 7098
rect 27076 7046 27098 7098
rect 27098 7046 27110 7098
rect 27110 7046 27132 7098
rect 27156 7046 27162 7098
rect 27162 7046 27174 7098
rect 27174 7046 27212 7098
rect 27236 7046 27238 7098
rect 27238 7046 27290 7098
rect 27290 7046 27292 7098
rect 26916 7044 26972 7046
rect 26996 7044 27052 7046
rect 27076 7044 27132 7046
rect 27156 7044 27212 7046
rect 27236 7044 27292 7046
rect 19656 6554 19712 6556
rect 19736 6554 19792 6556
rect 19816 6554 19872 6556
rect 19896 6554 19952 6556
rect 19976 6554 20032 6556
rect 19656 6502 19658 6554
rect 19658 6502 19710 6554
rect 19710 6502 19712 6554
rect 19736 6502 19774 6554
rect 19774 6502 19786 6554
rect 19786 6502 19792 6554
rect 19816 6502 19838 6554
rect 19838 6502 19850 6554
rect 19850 6502 19872 6554
rect 19896 6502 19902 6554
rect 19902 6502 19914 6554
rect 19914 6502 19952 6554
rect 19976 6502 19978 6554
rect 19978 6502 20030 6554
rect 20030 6502 20032 6554
rect 19656 6500 19712 6502
rect 19736 6500 19792 6502
rect 19816 6500 19872 6502
rect 19896 6500 19952 6502
rect 19976 6500 20032 6502
rect 27656 6554 27712 6556
rect 27736 6554 27792 6556
rect 27816 6554 27872 6556
rect 27896 6554 27952 6556
rect 27976 6554 28032 6556
rect 27656 6502 27658 6554
rect 27658 6502 27710 6554
rect 27710 6502 27712 6554
rect 27736 6502 27774 6554
rect 27774 6502 27786 6554
rect 27786 6502 27792 6554
rect 27816 6502 27838 6554
rect 27838 6502 27850 6554
rect 27850 6502 27872 6554
rect 27896 6502 27902 6554
rect 27902 6502 27914 6554
rect 27914 6502 27952 6554
rect 27976 6502 27978 6554
rect 27978 6502 28030 6554
rect 28030 6502 28032 6554
rect 27656 6500 27712 6502
rect 27736 6500 27792 6502
rect 27816 6500 27872 6502
rect 27896 6500 27952 6502
rect 27976 6500 28032 6502
rect 28354 6296 28410 6352
rect 18916 6010 18972 6012
rect 18996 6010 19052 6012
rect 19076 6010 19132 6012
rect 19156 6010 19212 6012
rect 19236 6010 19292 6012
rect 18916 5958 18918 6010
rect 18918 5958 18970 6010
rect 18970 5958 18972 6010
rect 18996 5958 19034 6010
rect 19034 5958 19046 6010
rect 19046 5958 19052 6010
rect 19076 5958 19098 6010
rect 19098 5958 19110 6010
rect 19110 5958 19132 6010
rect 19156 5958 19162 6010
rect 19162 5958 19174 6010
rect 19174 5958 19212 6010
rect 19236 5958 19238 6010
rect 19238 5958 19290 6010
rect 19290 5958 19292 6010
rect 18916 5956 18972 5958
rect 18996 5956 19052 5958
rect 19076 5956 19132 5958
rect 19156 5956 19212 5958
rect 19236 5956 19292 5958
rect 26916 6010 26972 6012
rect 26996 6010 27052 6012
rect 27076 6010 27132 6012
rect 27156 6010 27212 6012
rect 27236 6010 27292 6012
rect 26916 5958 26918 6010
rect 26918 5958 26970 6010
rect 26970 5958 26972 6010
rect 26996 5958 27034 6010
rect 27034 5958 27046 6010
rect 27046 5958 27052 6010
rect 27076 5958 27098 6010
rect 27098 5958 27110 6010
rect 27110 5958 27132 6010
rect 27156 5958 27162 6010
rect 27162 5958 27174 6010
rect 27174 5958 27212 6010
rect 27236 5958 27238 6010
rect 27238 5958 27290 6010
rect 27290 5958 27292 6010
rect 26916 5956 26972 5958
rect 26996 5956 27052 5958
rect 27076 5956 27132 5958
rect 27156 5956 27212 5958
rect 27236 5956 27292 5958
rect 28354 5480 28410 5536
rect 19656 5466 19712 5468
rect 19736 5466 19792 5468
rect 19816 5466 19872 5468
rect 19896 5466 19952 5468
rect 19976 5466 20032 5468
rect 19656 5414 19658 5466
rect 19658 5414 19710 5466
rect 19710 5414 19712 5466
rect 19736 5414 19774 5466
rect 19774 5414 19786 5466
rect 19786 5414 19792 5466
rect 19816 5414 19838 5466
rect 19838 5414 19850 5466
rect 19850 5414 19872 5466
rect 19896 5414 19902 5466
rect 19902 5414 19914 5466
rect 19914 5414 19952 5466
rect 19976 5414 19978 5466
rect 19978 5414 20030 5466
rect 20030 5414 20032 5466
rect 19656 5412 19712 5414
rect 19736 5412 19792 5414
rect 19816 5412 19872 5414
rect 19896 5412 19952 5414
rect 19976 5412 20032 5414
rect 27656 5466 27712 5468
rect 27736 5466 27792 5468
rect 27816 5466 27872 5468
rect 27896 5466 27952 5468
rect 27976 5466 28032 5468
rect 27656 5414 27658 5466
rect 27658 5414 27710 5466
rect 27710 5414 27712 5466
rect 27736 5414 27774 5466
rect 27774 5414 27786 5466
rect 27786 5414 27792 5466
rect 27816 5414 27838 5466
rect 27838 5414 27850 5466
rect 27850 5414 27872 5466
rect 27896 5414 27902 5466
rect 27902 5414 27914 5466
rect 27914 5414 27952 5466
rect 27976 5414 27978 5466
rect 27978 5414 28030 5466
rect 28030 5414 28032 5466
rect 27656 5412 27712 5414
rect 27736 5412 27792 5414
rect 27816 5412 27872 5414
rect 27896 5412 27952 5414
rect 27976 5412 28032 5414
rect 18916 4922 18972 4924
rect 18996 4922 19052 4924
rect 19076 4922 19132 4924
rect 19156 4922 19212 4924
rect 19236 4922 19292 4924
rect 18916 4870 18918 4922
rect 18918 4870 18970 4922
rect 18970 4870 18972 4922
rect 18996 4870 19034 4922
rect 19034 4870 19046 4922
rect 19046 4870 19052 4922
rect 19076 4870 19098 4922
rect 19098 4870 19110 4922
rect 19110 4870 19132 4922
rect 19156 4870 19162 4922
rect 19162 4870 19174 4922
rect 19174 4870 19212 4922
rect 19236 4870 19238 4922
rect 19238 4870 19290 4922
rect 19290 4870 19292 4922
rect 18916 4868 18972 4870
rect 18996 4868 19052 4870
rect 19076 4868 19132 4870
rect 19156 4868 19212 4870
rect 19236 4868 19292 4870
rect 26916 4922 26972 4924
rect 26996 4922 27052 4924
rect 27076 4922 27132 4924
rect 27156 4922 27212 4924
rect 27236 4922 27292 4924
rect 26916 4870 26918 4922
rect 26918 4870 26970 4922
rect 26970 4870 26972 4922
rect 26996 4870 27034 4922
rect 27034 4870 27046 4922
rect 27046 4870 27052 4922
rect 27076 4870 27098 4922
rect 27098 4870 27110 4922
rect 27110 4870 27132 4922
rect 27156 4870 27162 4922
rect 27162 4870 27174 4922
rect 27174 4870 27212 4922
rect 27236 4870 27238 4922
rect 27238 4870 27290 4922
rect 27290 4870 27292 4922
rect 26916 4868 26972 4870
rect 26996 4868 27052 4870
rect 27076 4868 27132 4870
rect 27156 4868 27212 4870
rect 27236 4868 27292 4870
rect 19656 4378 19712 4380
rect 19736 4378 19792 4380
rect 19816 4378 19872 4380
rect 19896 4378 19952 4380
rect 19976 4378 20032 4380
rect 19656 4326 19658 4378
rect 19658 4326 19710 4378
rect 19710 4326 19712 4378
rect 19736 4326 19774 4378
rect 19774 4326 19786 4378
rect 19786 4326 19792 4378
rect 19816 4326 19838 4378
rect 19838 4326 19850 4378
rect 19850 4326 19872 4378
rect 19896 4326 19902 4378
rect 19902 4326 19914 4378
rect 19914 4326 19952 4378
rect 19976 4326 19978 4378
rect 19978 4326 20030 4378
rect 20030 4326 20032 4378
rect 19656 4324 19712 4326
rect 19736 4324 19792 4326
rect 19816 4324 19872 4326
rect 19896 4324 19952 4326
rect 19976 4324 20032 4326
rect 27656 4378 27712 4380
rect 27736 4378 27792 4380
rect 27816 4378 27872 4380
rect 27896 4378 27952 4380
rect 27976 4378 28032 4380
rect 27656 4326 27658 4378
rect 27658 4326 27710 4378
rect 27710 4326 27712 4378
rect 27736 4326 27774 4378
rect 27774 4326 27786 4378
rect 27786 4326 27792 4378
rect 27816 4326 27838 4378
rect 27838 4326 27850 4378
rect 27850 4326 27872 4378
rect 27896 4326 27902 4378
rect 27902 4326 27914 4378
rect 27914 4326 27952 4378
rect 27976 4326 27978 4378
rect 27978 4326 28030 4378
rect 28030 4326 28032 4378
rect 27656 4324 27712 4326
rect 27736 4324 27792 4326
rect 27816 4324 27872 4326
rect 27896 4324 27952 4326
rect 27976 4324 28032 4326
rect 28354 4664 28410 4720
rect 28354 3848 28410 3904
rect 18916 3834 18972 3836
rect 18996 3834 19052 3836
rect 19076 3834 19132 3836
rect 19156 3834 19212 3836
rect 19236 3834 19292 3836
rect 18916 3782 18918 3834
rect 18918 3782 18970 3834
rect 18970 3782 18972 3834
rect 18996 3782 19034 3834
rect 19034 3782 19046 3834
rect 19046 3782 19052 3834
rect 19076 3782 19098 3834
rect 19098 3782 19110 3834
rect 19110 3782 19132 3834
rect 19156 3782 19162 3834
rect 19162 3782 19174 3834
rect 19174 3782 19212 3834
rect 19236 3782 19238 3834
rect 19238 3782 19290 3834
rect 19290 3782 19292 3834
rect 18916 3780 18972 3782
rect 18996 3780 19052 3782
rect 19076 3780 19132 3782
rect 19156 3780 19212 3782
rect 19236 3780 19292 3782
rect 26916 3834 26972 3836
rect 26996 3834 27052 3836
rect 27076 3834 27132 3836
rect 27156 3834 27212 3836
rect 27236 3834 27292 3836
rect 26916 3782 26918 3834
rect 26918 3782 26970 3834
rect 26970 3782 26972 3834
rect 26996 3782 27034 3834
rect 27034 3782 27046 3834
rect 27046 3782 27052 3834
rect 27076 3782 27098 3834
rect 27098 3782 27110 3834
rect 27110 3782 27132 3834
rect 27156 3782 27162 3834
rect 27162 3782 27174 3834
rect 27174 3782 27212 3834
rect 27236 3782 27238 3834
rect 27238 3782 27290 3834
rect 27290 3782 27292 3834
rect 26916 3780 26972 3782
rect 26996 3780 27052 3782
rect 27076 3780 27132 3782
rect 27156 3780 27212 3782
rect 27236 3780 27292 3782
rect 11656 3290 11712 3292
rect 11736 3290 11792 3292
rect 11816 3290 11872 3292
rect 11896 3290 11952 3292
rect 11976 3290 12032 3292
rect 11656 3238 11658 3290
rect 11658 3238 11710 3290
rect 11710 3238 11712 3290
rect 11736 3238 11774 3290
rect 11774 3238 11786 3290
rect 11786 3238 11792 3290
rect 11816 3238 11838 3290
rect 11838 3238 11850 3290
rect 11850 3238 11872 3290
rect 11896 3238 11902 3290
rect 11902 3238 11914 3290
rect 11914 3238 11952 3290
rect 11976 3238 11978 3290
rect 11978 3238 12030 3290
rect 12030 3238 12032 3290
rect 11656 3236 11712 3238
rect 11736 3236 11792 3238
rect 11816 3236 11872 3238
rect 11896 3236 11952 3238
rect 11976 3236 12032 3238
rect 2916 2746 2972 2748
rect 2996 2746 3052 2748
rect 3076 2746 3132 2748
rect 3156 2746 3212 2748
rect 3236 2746 3292 2748
rect 2916 2694 2918 2746
rect 2918 2694 2970 2746
rect 2970 2694 2972 2746
rect 2996 2694 3034 2746
rect 3034 2694 3046 2746
rect 3046 2694 3052 2746
rect 3076 2694 3098 2746
rect 3098 2694 3110 2746
rect 3110 2694 3132 2746
rect 3156 2694 3162 2746
rect 3162 2694 3174 2746
rect 3174 2694 3212 2746
rect 3236 2694 3238 2746
rect 3238 2694 3290 2746
rect 3290 2694 3292 2746
rect 2916 2692 2972 2694
rect 2996 2692 3052 2694
rect 3076 2692 3132 2694
rect 3156 2692 3212 2694
rect 3236 2692 3292 2694
rect 10916 2746 10972 2748
rect 10996 2746 11052 2748
rect 11076 2746 11132 2748
rect 11156 2746 11212 2748
rect 11236 2746 11292 2748
rect 10916 2694 10918 2746
rect 10918 2694 10970 2746
rect 10970 2694 10972 2746
rect 10996 2694 11034 2746
rect 11034 2694 11046 2746
rect 11046 2694 11052 2746
rect 11076 2694 11098 2746
rect 11098 2694 11110 2746
rect 11110 2694 11132 2746
rect 11156 2694 11162 2746
rect 11162 2694 11174 2746
rect 11174 2694 11212 2746
rect 11236 2694 11238 2746
rect 11238 2694 11290 2746
rect 11290 2694 11292 2746
rect 10916 2692 10972 2694
rect 10996 2692 11052 2694
rect 11076 2692 11132 2694
rect 11156 2692 11212 2694
rect 11236 2692 11292 2694
rect 846 2624 902 2680
rect 19656 3290 19712 3292
rect 19736 3290 19792 3292
rect 19816 3290 19872 3292
rect 19896 3290 19952 3292
rect 19976 3290 20032 3292
rect 19656 3238 19658 3290
rect 19658 3238 19710 3290
rect 19710 3238 19712 3290
rect 19736 3238 19774 3290
rect 19774 3238 19786 3290
rect 19786 3238 19792 3290
rect 19816 3238 19838 3290
rect 19838 3238 19850 3290
rect 19850 3238 19872 3290
rect 19896 3238 19902 3290
rect 19902 3238 19914 3290
rect 19914 3238 19952 3290
rect 19976 3238 19978 3290
rect 19978 3238 20030 3290
rect 20030 3238 20032 3290
rect 19656 3236 19712 3238
rect 19736 3236 19792 3238
rect 19816 3236 19872 3238
rect 19896 3236 19952 3238
rect 19976 3236 20032 3238
rect 27656 3290 27712 3292
rect 27736 3290 27792 3292
rect 27816 3290 27872 3292
rect 27896 3290 27952 3292
rect 27976 3290 28032 3292
rect 27656 3238 27658 3290
rect 27658 3238 27710 3290
rect 27710 3238 27712 3290
rect 27736 3238 27774 3290
rect 27774 3238 27786 3290
rect 27786 3238 27792 3290
rect 27816 3238 27838 3290
rect 27838 3238 27850 3290
rect 27850 3238 27872 3290
rect 27896 3238 27902 3290
rect 27902 3238 27914 3290
rect 27914 3238 27952 3290
rect 27976 3238 27978 3290
rect 27978 3238 28030 3290
rect 28030 3238 28032 3290
rect 27656 3236 27712 3238
rect 27736 3236 27792 3238
rect 27816 3236 27872 3238
rect 27896 3236 27952 3238
rect 27976 3236 28032 3238
rect 28354 3032 28410 3088
rect 18916 2746 18972 2748
rect 18996 2746 19052 2748
rect 19076 2746 19132 2748
rect 19156 2746 19212 2748
rect 19236 2746 19292 2748
rect 18916 2694 18918 2746
rect 18918 2694 18970 2746
rect 18970 2694 18972 2746
rect 18996 2694 19034 2746
rect 19034 2694 19046 2746
rect 19046 2694 19052 2746
rect 19076 2694 19098 2746
rect 19098 2694 19110 2746
rect 19110 2694 19132 2746
rect 19156 2694 19162 2746
rect 19162 2694 19174 2746
rect 19174 2694 19212 2746
rect 19236 2694 19238 2746
rect 19238 2694 19290 2746
rect 19290 2694 19292 2746
rect 18916 2692 18972 2694
rect 18996 2692 19052 2694
rect 19076 2692 19132 2694
rect 19156 2692 19212 2694
rect 19236 2692 19292 2694
rect 26916 2746 26972 2748
rect 26996 2746 27052 2748
rect 27076 2746 27132 2748
rect 27156 2746 27212 2748
rect 27236 2746 27292 2748
rect 26916 2694 26918 2746
rect 26918 2694 26970 2746
rect 26970 2694 26972 2746
rect 26996 2694 27034 2746
rect 27034 2694 27046 2746
rect 27046 2694 27052 2746
rect 27076 2694 27098 2746
rect 27098 2694 27110 2746
rect 27110 2694 27132 2746
rect 27156 2694 27162 2746
rect 27162 2694 27174 2746
rect 27174 2694 27212 2746
rect 27236 2694 27238 2746
rect 27238 2694 27290 2746
rect 27290 2694 27292 2746
rect 26916 2692 26972 2694
rect 26996 2692 27052 2694
rect 27076 2692 27132 2694
rect 27156 2692 27212 2694
rect 27236 2692 27292 2694
rect 28354 2216 28410 2272
rect 3656 2202 3712 2204
rect 3736 2202 3792 2204
rect 3816 2202 3872 2204
rect 3896 2202 3952 2204
rect 3976 2202 4032 2204
rect 3656 2150 3658 2202
rect 3658 2150 3710 2202
rect 3710 2150 3712 2202
rect 3736 2150 3774 2202
rect 3774 2150 3786 2202
rect 3786 2150 3792 2202
rect 3816 2150 3838 2202
rect 3838 2150 3850 2202
rect 3850 2150 3872 2202
rect 3896 2150 3902 2202
rect 3902 2150 3914 2202
rect 3914 2150 3952 2202
rect 3976 2150 3978 2202
rect 3978 2150 4030 2202
rect 4030 2150 4032 2202
rect 3656 2148 3712 2150
rect 3736 2148 3792 2150
rect 3816 2148 3872 2150
rect 3896 2148 3952 2150
rect 3976 2148 4032 2150
rect 11656 2202 11712 2204
rect 11736 2202 11792 2204
rect 11816 2202 11872 2204
rect 11896 2202 11952 2204
rect 11976 2202 12032 2204
rect 11656 2150 11658 2202
rect 11658 2150 11710 2202
rect 11710 2150 11712 2202
rect 11736 2150 11774 2202
rect 11774 2150 11786 2202
rect 11786 2150 11792 2202
rect 11816 2150 11838 2202
rect 11838 2150 11850 2202
rect 11850 2150 11872 2202
rect 11896 2150 11902 2202
rect 11902 2150 11914 2202
rect 11914 2150 11952 2202
rect 11976 2150 11978 2202
rect 11978 2150 12030 2202
rect 12030 2150 12032 2202
rect 11656 2148 11712 2150
rect 11736 2148 11792 2150
rect 11816 2148 11872 2150
rect 11896 2148 11952 2150
rect 11976 2148 12032 2150
rect 19656 2202 19712 2204
rect 19736 2202 19792 2204
rect 19816 2202 19872 2204
rect 19896 2202 19952 2204
rect 19976 2202 20032 2204
rect 19656 2150 19658 2202
rect 19658 2150 19710 2202
rect 19710 2150 19712 2202
rect 19736 2150 19774 2202
rect 19774 2150 19786 2202
rect 19786 2150 19792 2202
rect 19816 2150 19838 2202
rect 19838 2150 19850 2202
rect 19850 2150 19872 2202
rect 19896 2150 19902 2202
rect 19902 2150 19914 2202
rect 19914 2150 19952 2202
rect 19976 2150 19978 2202
rect 19978 2150 20030 2202
rect 20030 2150 20032 2202
rect 19656 2148 19712 2150
rect 19736 2148 19792 2150
rect 19816 2148 19872 2150
rect 19896 2148 19952 2150
rect 19976 2148 20032 2150
rect 27656 2202 27712 2204
rect 27736 2202 27792 2204
rect 27816 2202 27872 2204
rect 27896 2202 27952 2204
rect 27976 2202 28032 2204
rect 27656 2150 27658 2202
rect 27658 2150 27710 2202
rect 27710 2150 27712 2202
rect 27736 2150 27774 2202
rect 27774 2150 27786 2202
rect 27786 2150 27792 2202
rect 27816 2150 27838 2202
rect 27838 2150 27850 2202
rect 27850 2150 27872 2202
rect 27896 2150 27902 2202
rect 27902 2150 27914 2202
rect 27914 2150 27952 2202
rect 27976 2150 27978 2202
rect 27978 2150 28030 2202
rect 28030 2150 28032 2202
rect 27656 2148 27712 2150
rect 27736 2148 27792 2150
rect 27816 2148 27872 2150
rect 27896 2148 27952 2150
rect 27976 2148 28032 2150
rect 846 1808 902 1864
rect 110 1128 166 1184
<< metal3 >>
rect 0 28658 800 28688
rect 1025 28658 1091 28661
rect 0 28656 1091 28658
rect 0 28600 1030 28656
rect 1086 28600 1091 28656
rect 0 28598 1091 28600
rect 0 28568 800 28598
rect 1025 28595 1091 28598
rect 0 27842 800 27872
rect 933 27842 999 27845
rect 0 27840 999 27842
rect 0 27784 938 27840
rect 994 27784 999 27840
rect 0 27782 999 27784
rect 0 27752 800 27782
rect 933 27779 999 27782
rect 2906 27776 3302 27777
rect 2906 27712 2912 27776
rect 2976 27712 2992 27776
rect 3056 27712 3072 27776
rect 3136 27712 3152 27776
rect 3216 27712 3232 27776
rect 3296 27712 3302 27776
rect 2906 27711 3302 27712
rect 10906 27776 11302 27777
rect 10906 27712 10912 27776
rect 10976 27712 10992 27776
rect 11056 27712 11072 27776
rect 11136 27712 11152 27776
rect 11216 27712 11232 27776
rect 11296 27712 11302 27776
rect 10906 27711 11302 27712
rect 18906 27776 19302 27777
rect 18906 27712 18912 27776
rect 18976 27712 18992 27776
rect 19056 27712 19072 27776
rect 19136 27712 19152 27776
rect 19216 27712 19232 27776
rect 19296 27712 19302 27776
rect 18906 27711 19302 27712
rect 26906 27776 27302 27777
rect 26906 27712 26912 27776
rect 26976 27712 26992 27776
rect 27056 27712 27072 27776
rect 27136 27712 27152 27776
rect 27216 27712 27232 27776
rect 27296 27712 27302 27776
rect 26906 27711 27302 27712
rect 28349 27570 28415 27573
rect 29200 27570 30000 27600
rect 28349 27568 30000 27570
rect 28349 27512 28354 27568
rect 28410 27512 30000 27568
rect 28349 27510 30000 27512
rect 28349 27507 28415 27510
rect 29200 27480 30000 27510
rect 3646 27232 4042 27233
rect 3646 27168 3652 27232
rect 3716 27168 3732 27232
rect 3796 27168 3812 27232
rect 3876 27168 3892 27232
rect 3956 27168 3972 27232
rect 4036 27168 4042 27232
rect 3646 27167 4042 27168
rect 11646 27232 12042 27233
rect 11646 27168 11652 27232
rect 11716 27168 11732 27232
rect 11796 27168 11812 27232
rect 11876 27168 11892 27232
rect 11956 27168 11972 27232
rect 12036 27168 12042 27232
rect 11646 27167 12042 27168
rect 19646 27232 20042 27233
rect 19646 27168 19652 27232
rect 19716 27168 19732 27232
rect 19796 27168 19812 27232
rect 19876 27168 19892 27232
rect 19956 27168 19972 27232
rect 20036 27168 20042 27232
rect 19646 27167 20042 27168
rect 27646 27232 28042 27233
rect 27646 27168 27652 27232
rect 27716 27168 27732 27232
rect 27796 27168 27812 27232
rect 27876 27168 27892 27232
rect 27956 27168 27972 27232
rect 28036 27168 28042 27232
rect 27646 27167 28042 27168
rect 841 27162 907 27165
rect 798 27160 907 27162
rect 798 27104 846 27160
rect 902 27104 907 27160
rect 798 27099 907 27104
rect 798 27056 858 27099
rect 0 26966 858 27056
rect 0 26936 800 26966
rect 28349 26754 28415 26757
rect 29200 26754 30000 26784
rect 28349 26752 30000 26754
rect 28349 26696 28354 26752
rect 28410 26696 30000 26752
rect 28349 26694 30000 26696
rect 28349 26691 28415 26694
rect 2906 26688 3302 26689
rect 2906 26624 2912 26688
rect 2976 26624 2992 26688
rect 3056 26624 3072 26688
rect 3136 26624 3152 26688
rect 3216 26624 3232 26688
rect 3296 26624 3302 26688
rect 2906 26623 3302 26624
rect 10906 26688 11302 26689
rect 10906 26624 10912 26688
rect 10976 26624 10992 26688
rect 11056 26624 11072 26688
rect 11136 26624 11152 26688
rect 11216 26624 11232 26688
rect 11296 26624 11302 26688
rect 10906 26623 11302 26624
rect 18906 26688 19302 26689
rect 18906 26624 18912 26688
rect 18976 26624 18992 26688
rect 19056 26624 19072 26688
rect 19136 26624 19152 26688
rect 19216 26624 19232 26688
rect 19296 26624 19302 26688
rect 18906 26623 19302 26624
rect 26906 26688 27302 26689
rect 26906 26624 26912 26688
rect 26976 26624 26992 26688
rect 27056 26624 27072 26688
rect 27136 26624 27152 26688
rect 27216 26624 27232 26688
rect 27296 26624 27302 26688
rect 29200 26664 30000 26694
rect 26906 26623 27302 26624
rect 0 26210 800 26240
rect 0 26120 858 26210
rect 798 26077 858 26120
rect 3646 26144 4042 26145
rect 3646 26080 3652 26144
rect 3716 26080 3732 26144
rect 3796 26080 3812 26144
rect 3876 26080 3892 26144
rect 3956 26080 3972 26144
rect 4036 26080 4042 26144
rect 3646 26079 4042 26080
rect 11646 26144 12042 26145
rect 11646 26080 11652 26144
rect 11716 26080 11732 26144
rect 11796 26080 11812 26144
rect 11876 26080 11892 26144
rect 11956 26080 11972 26144
rect 12036 26080 12042 26144
rect 11646 26079 12042 26080
rect 19646 26144 20042 26145
rect 19646 26080 19652 26144
rect 19716 26080 19732 26144
rect 19796 26080 19812 26144
rect 19876 26080 19892 26144
rect 19956 26080 19972 26144
rect 20036 26080 20042 26144
rect 19646 26079 20042 26080
rect 27646 26144 28042 26145
rect 27646 26080 27652 26144
rect 27716 26080 27732 26144
rect 27796 26080 27812 26144
rect 27876 26080 27892 26144
rect 27956 26080 27972 26144
rect 28036 26080 28042 26144
rect 27646 26079 28042 26080
rect 798 26072 907 26077
rect 798 26016 846 26072
rect 902 26016 907 26072
rect 798 26014 907 26016
rect 841 26011 907 26014
rect 28349 25938 28415 25941
rect 29200 25938 30000 25968
rect 28349 25936 30000 25938
rect 28349 25880 28354 25936
rect 28410 25880 30000 25936
rect 28349 25878 30000 25880
rect 28349 25875 28415 25878
rect 29200 25848 30000 25878
rect 2906 25600 3302 25601
rect 2906 25536 2912 25600
rect 2976 25536 2992 25600
rect 3056 25536 3072 25600
rect 3136 25536 3152 25600
rect 3216 25536 3232 25600
rect 3296 25536 3302 25600
rect 2906 25535 3302 25536
rect 10906 25600 11302 25601
rect 10906 25536 10912 25600
rect 10976 25536 10992 25600
rect 11056 25536 11072 25600
rect 11136 25536 11152 25600
rect 11216 25536 11232 25600
rect 11296 25536 11302 25600
rect 10906 25535 11302 25536
rect 18906 25600 19302 25601
rect 18906 25536 18912 25600
rect 18976 25536 18992 25600
rect 19056 25536 19072 25600
rect 19136 25536 19152 25600
rect 19216 25536 19232 25600
rect 19296 25536 19302 25600
rect 18906 25535 19302 25536
rect 26906 25600 27302 25601
rect 26906 25536 26912 25600
rect 26976 25536 26992 25600
rect 27056 25536 27072 25600
rect 27136 25536 27152 25600
rect 27216 25536 27232 25600
rect 27296 25536 27302 25600
rect 26906 25535 27302 25536
rect 841 25530 907 25533
rect 798 25528 907 25530
rect 798 25472 846 25528
rect 902 25472 907 25528
rect 798 25467 907 25472
rect 798 25424 858 25467
rect 0 25334 858 25424
rect 0 25304 800 25334
rect 28349 25122 28415 25125
rect 29200 25122 30000 25152
rect 28349 25120 30000 25122
rect 28349 25064 28354 25120
rect 28410 25064 30000 25120
rect 28349 25062 30000 25064
rect 28349 25059 28415 25062
rect 3646 25056 4042 25057
rect 3646 24992 3652 25056
rect 3716 24992 3732 25056
rect 3796 24992 3812 25056
rect 3876 24992 3892 25056
rect 3956 24992 3972 25056
rect 4036 24992 4042 25056
rect 3646 24991 4042 24992
rect 11646 25056 12042 25057
rect 11646 24992 11652 25056
rect 11716 24992 11732 25056
rect 11796 24992 11812 25056
rect 11876 24992 11892 25056
rect 11956 24992 11972 25056
rect 12036 24992 12042 25056
rect 11646 24991 12042 24992
rect 19646 25056 20042 25057
rect 19646 24992 19652 25056
rect 19716 24992 19732 25056
rect 19796 24992 19812 25056
rect 19876 24992 19892 25056
rect 19956 24992 19972 25056
rect 20036 24992 20042 25056
rect 19646 24991 20042 24992
rect 27646 25056 28042 25057
rect 27646 24992 27652 25056
rect 27716 24992 27732 25056
rect 27796 24992 27812 25056
rect 27876 24992 27892 25056
rect 27956 24992 27972 25056
rect 28036 24992 28042 25056
rect 29200 25032 30000 25062
rect 27646 24991 28042 24992
rect 841 24714 907 24717
rect 798 24712 907 24714
rect 798 24656 846 24712
rect 902 24656 907 24712
rect 798 24651 907 24656
rect 798 24608 858 24651
rect 0 24518 858 24608
rect 0 24488 800 24518
rect 2906 24512 3302 24513
rect 2906 24448 2912 24512
rect 2976 24448 2992 24512
rect 3056 24448 3072 24512
rect 3136 24448 3152 24512
rect 3216 24448 3232 24512
rect 3296 24448 3302 24512
rect 2906 24447 3302 24448
rect 10906 24512 11302 24513
rect 10906 24448 10912 24512
rect 10976 24448 10992 24512
rect 11056 24448 11072 24512
rect 11136 24448 11152 24512
rect 11216 24448 11232 24512
rect 11296 24448 11302 24512
rect 10906 24447 11302 24448
rect 18906 24512 19302 24513
rect 18906 24448 18912 24512
rect 18976 24448 18992 24512
rect 19056 24448 19072 24512
rect 19136 24448 19152 24512
rect 19216 24448 19232 24512
rect 19296 24448 19302 24512
rect 18906 24447 19302 24448
rect 26906 24512 27302 24513
rect 26906 24448 26912 24512
rect 26976 24448 26992 24512
rect 27056 24448 27072 24512
rect 27136 24448 27152 24512
rect 27216 24448 27232 24512
rect 27296 24448 27302 24512
rect 26906 24447 27302 24448
rect 28349 24306 28415 24309
rect 29200 24306 30000 24336
rect 28349 24304 30000 24306
rect 28349 24248 28354 24304
rect 28410 24248 30000 24304
rect 28349 24246 30000 24248
rect 28349 24243 28415 24246
rect 29200 24216 30000 24246
rect 3646 23968 4042 23969
rect 3646 23904 3652 23968
rect 3716 23904 3732 23968
rect 3796 23904 3812 23968
rect 3876 23904 3892 23968
rect 3956 23904 3972 23968
rect 4036 23904 4042 23968
rect 3646 23903 4042 23904
rect 11646 23968 12042 23969
rect 11646 23904 11652 23968
rect 11716 23904 11732 23968
rect 11796 23904 11812 23968
rect 11876 23904 11892 23968
rect 11956 23904 11972 23968
rect 12036 23904 12042 23968
rect 11646 23903 12042 23904
rect 19646 23968 20042 23969
rect 19646 23904 19652 23968
rect 19716 23904 19732 23968
rect 19796 23904 19812 23968
rect 19876 23904 19892 23968
rect 19956 23904 19972 23968
rect 20036 23904 20042 23968
rect 19646 23903 20042 23904
rect 27646 23968 28042 23969
rect 27646 23904 27652 23968
rect 27716 23904 27732 23968
rect 27796 23904 27812 23968
rect 27876 23904 27892 23968
rect 27956 23904 27972 23968
rect 28036 23904 28042 23968
rect 27646 23903 28042 23904
rect 841 23898 907 23901
rect 798 23896 907 23898
rect 798 23840 846 23896
rect 902 23840 907 23896
rect 798 23835 907 23840
rect 798 23792 858 23835
rect 0 23702 858 23792
rect 0 23672 800 23702
rect 28349 23490 28415 23493
rect 29200 23490 30000 23520
rect 28349 23488 30000 23490
rect 28349 23432 28354 23488
rect 28410 23432 30000 23488
rect 28349 23430 30000 23432
rect 28349 23427 28415 23430
rect 2906 23424 3302 23425
rect 2906 23360 2912 23424
rect 2976 23360 2992 23424
rect 3056 23360 3072 23424
rect 3136 23360 3152 23424
rect 3216 23360 3232 23424
rect 3296 23360 3302 23424
rect 2906 23359 3302 23360
rect 10906 23424 11302 23425
rect 10906 23360 10912 23424
rect 10976 23360 10992 23424
rect 11056 23360 11072 23424
rect 11136 23360 11152 23424
rect 11216 23360 11232 23424
rect 11296 23360 11302 23424
rect 10906 23359 11302 23360
rect 18906 23424 19302 23425
rect 18906 23360 18912 23424
rect 18976 23360 18992 23424
rect 19056 23360 19072 23424
rect 19136 23360 19152 23424
rect 19216 23360 19232 23424
rect 19296 23360 19302 23424
rect 18906 23359 19302 23360
rect 26906 23424 27302 23425
rect 26906 23360 26912 23424
rect 26976 23360 26992 23424
rect 27056 23360 27072 23424
rect 27136 23360 27152 23424
rect 27216 23360 27232 23424
rect 27296 23360 27302 23424
rect 29200 23400 30000 23430
rect 26906 23359 27302 23360
rect 841 23082 907 23085
rect 798 23080 907 23082
rect 798 23024 846 23080
rect 902 23024 907 23080
rect 798 23019 907 23024
rect 798 22976 858 23019
rect 0 22886 858 22976
rect 0 22856 800 22886
rect 3646 22880 4042 22881
rect 3646 22816 3652 22880
rect 3716 22816 3732 22880
rect 3796 22816 3812 22880
rect 3876 22816 3892 22880
rect 3956 22816 3972 22880
rect 4036 22816 4042 22880
rect 3646 22815 4042 22816
rect 11646 22880 12042 22881
rect 11646 22816 11652 22880
rect 11716 22816 11732 22880
rect 11796 22816 11812 22880
rect 11876 22816 11892 22880
rect 11956 22816 11972 22880
rect 12036 22816 12042 22880
rect 11646 22815 12042 22816
rect 19646 22880 20042 22881
rect 19646 22816 19652 22880
rect 19716 22816 19732 22880
rect 19796 22816 19812 22880
rect 19876 22816 19892 22880
rect 19956 22816 19972 22880
rect 20036 22816 20042 22880
rect 19646 22815 20042 22816
rect 27646 22880 28042 22881
rect 27646 22816 27652 22880
rect 27716 22816 27732 22880
rect 27796 22816 27812 22880
rect 27876 22816 27892 22880
rect 27956 22816 27972 22880
rect 28036 22816 28042 22880
rect 27646 22815 28042 22816
rect 28349 22674 28415 22677
rect 29200 22674 30000 22704
rect 28349 22672 30000 22674
rect 28349 22616 28354 22672
rect 28410 22616 30000 22672
rect 28349 22614 30000 22616
rect 28349 22611 28415 22614
rect 29200 22584 30000 22614
rect 2906 22336 3302 22337
rect 2906 22272 2912 22336
rect 2976 22272 2992 22336
rect 3056 22272 3072 22336
rect 3136 22272 3152 22336
rect 3216 22272 3232 22336
rect 3296 22272 3302 22336
rect 2906 22271 3302 22272
rect 10906 22336 11302 22337
rect 10906 22272 10912 22336
rect 10976 22272 10992 22336
rect 11056 22272 11072 22336
rect 11136 22272 11152 22336
rect 11216 22272 11232 22336
rect 11296 22272 11302 22336
rect 10906 22271 11302 22272
rect 18906 22336 19302 22337
rect 18906 22272 18912 22336
rect 18976 22272 18992 22336
rect 19056 22272 19072 22336
rect 19136 22272 19152 22336
rect 19216 22272 19232 22336
rect 19296 22272 19302 22336
rect 18906 22271 19302 22272
rect 26906 22336 27302 22337
rect 26906 22272 26912 22336
rect 26976 22272 26992 22336
rect 27056 22272 27072 22336
rect 27136 22272 27152 22336
rect 27216 22272 27232 22336
rect 27296 22272 27302 22336
rect 26906 22271 27302 22272
rect 841 22266 907 22269
rect 798 22264 907 22266
rect 798 22208 846 22264
rect 902 22208 907 22264
rect 798 22203 907 22208
rect 798 22160 858 22203
rect 0 22070 858 22160
rect 0 22040 800 22070
rect 28349 21858 28415 21861
rect 29200 21858 30000 21888
rect 28349 21856 30000 21858
rect 28349 21800 28354 21856
rect 28410 21800 30000 21856
rect 28349 21798 30000 21800
rect 28349 21795 28415 21798
rect 3646 21792 4042 21793
rect 3646 21728 3652 21792
rect 3716 21728 3732 21792
rect 3796 21728 3812 21792
rect 3876 21728 3892 21792
rect 3956 21728 3972 21792
rect 4036 21728 4042 21792
rect 3646 21727 4042 21728
rect 11646 21792 12042 21793
rect 11646 21728 11652 21792
rect 11716 21728 11732 21792
rect 11796 21728 11812 21792
rect 11876 21728 11892 21792
rect 11956 21728 11972 21792
rect 12036 21728 12042 21792
rect 11646 21727 12042 21728
rect 19646 21792 20042 21793
rect 19646 21728 19652 21792
rect 19716 21728 19732 21792
rect 19796 21728 19812 21792
rect 19876 21728 19892 21792
rect 19956 21728 19972 21792
rect 20036 21728 20042 21792
rect 19646 21727 20042 21728
rect 27646 21792 28042 21793
rect 27646 21728 27652 21792
rect 27716 21728 27732 21792
rect 27796 21728 27812 21792
rect 27876 21728 27892 21792
rect 27956 21728 27972 21792
rect 28036 21728 28042 21792
rect 29200 21768 30000 21798
rect 27646 21727 28042 21728
rect 1393 21450 1459 21453
rect 798 21448 1459 21450
rect 798 21392 1398 21448
rect 1454 21392 1459 21448
rect 798 21390 1459 21392
rect 798 21344 858 21390
rect 1393 21387 1459 21390
rect 0 21254 858 21344
rect 0 21224 800 21254
rect 2906 21248 3302 21249
rect 2906 21184 2912 21248
rect 2976 21184 2992 21248
rect 3056 21184 3072 21248
rect 3136 21184 3152 21248
rect 3216 21184 3232 21248
rect 3296 21184 3302 21248
rect 2906 21183 3302 21184
rect 10906 21248 11302 21249
rect 10906 21184 10912 21248
rect 10976 21184 10992 21248
rect 11056 21184 11072 21248
rect 11136 21184 11152 21248
rect 11216 21184 11232 21248
rect 11296 21184 11302 21248
rect 10906 21183 11302 21184
rect 18906 21248 19302 21249
rect 18906 21184 18912 21248
rect 18976 21184 18992 21248
rect 19056 21184 19072 21248
rect 19136 21184 19152 21248
rect 19216 21184 19232 21248
rect 19296 21184 19302 21248
rect 18906 21183 19302 21184
rect 26906 21248 27302 21249
rect 26906 21184 26912 21248
rect 26976 21184 26992 21248
rect 27056 21184 27072 21248
rect 27136 21184 27152 21248
rect 27216 21184 27232 21248
rect 27296 21184 27302 21248
rect 26906 21183 27302 21184
rect 28349 21042 28415 21045
rect 29200 21042 30000 21072
rect 28349 21040 30000 21042
rect 28349 20984 28354 21040
rect 28410 20984 30000 21040
rect 28349 20982 30000 20984
rect 28349 20979 28415 20982
rect 29200 20952 30000 20982
rect 3646 20704 4042 20705
rect 3646 20640 3652 20704
rect 3716 20640 3732 20704
rect 3796 20640 3812 20704
rect 3876 20640 3892 20704
rect 3956 20640 3972 20704
rect 4036 20640 4042 20704
rect 3646 20639 4042 20640
rect 11646 20704 12042 20705
rect 11646 20640 11652 20704
rect 11716 20640 11732 20704
rect 11796 20640 11812 20704
rect 11876 20640 11892 20704
rect 11956 20640 11972 20704
rect 12036 20640 12042 20704
rect 11646 20639 12042 20640
rect 19646 20704 20042 20705
rect 19646 20640 19652 20704
rect 19716 20640 19732 20704
rect 19796 20640 19812 20704
rect 19876 20640 19892 20704
rect 19956 20640 19972 20704
rect 20036 20640 20042 20704
rect 19646 20639 20042 20640
rect 27646 20704 28042 20705
rect 27646 20640 27652 20704
rect 27716 20640 27732 20704
rect 27796 20640 27812 20704
rect 27876 20640 27892 20704
rect 27956 20640 27972 20704
rect 28036 20640 28042 20704
rect 27646 20639 28042 20640
rect 1393 20634 1459 20637
rect 798 20632 1459 20634
rect 798 20576 1398 20632
rect 1454 20576 1459 20632
rect 798 20574 1459 20576
rect 798 20528 858 20574
rect 1393 20571 1459 20574
rect 0 20438 858 20528
rect 0 20408 800 20438
rect 28349 20226 28415 20229
rect 29200 20226 30000 20256
rect 28349 20224 30000 20226
rect 28349 20168 28354 20224
rect 28410 20168 30000 20224
rect 28349 20166 30000 20168
rect 28349 20163 28415 20166
rect 2906 20160 3302 20161
rect 2906 20096 2912 20160
rect 2976 20096 2992 20160
rect 3056 20096 3072 20160
rect 3136 20096 3152 20160
rect 3216 20096 3232 20160
rect 3296 20096 3302 20160
rect 2906 20095 3302 20096
rect 10906 20160 11302 20161
rect 10906 20096 10912 20160
rect 10976 20096 10992 20160
rect 11056 20096 11072 20160
rect 11136 20096 11152 20160
rect 11216 20096 11232 20160
rect 11296 20096 11302 20160
rect 10906 20095 11302 20096
rect 18906 20160 19302 20161
rect 18906 20096 18912 20160
rect 18976 20096 18992 20160
rect 19056 20096 19072 20160
rect 19136 20096 19152 20160
rect 19216 20096 19232 20160
rect 19296 20096 19302 20160
rect 18906 20095 19302 20096
rect 26906 20160 27302 20161
rect 26906 20096 26912 20160
rect 26976 20096 26992 20160
rect 27056 20096 27072 20160
rect 27136 20096 27152 20160
rect 27216 20096 27232 20160
rect 27296 20096 27302 20160
rect 29200 20136 30000 20166
rect 26906 20095 27302 20096
rect 1393 19818 1459 19821
rect 798 19816 1459 19818
rect 798 19760 1398 19816
rect 1454 19760 1459 19816
rect 798 19758 1459 19760
rect 798 19712 858 19758
rect 1393 19755 1459 19758
rect 0 19622 858 19712
rect 0 19592 800 19622
rect 3646 19616 4042 19617
rect 3646 19552 3652 19616
rect 3716 19552 3732 19616
rect 3796 19552 3812 19616
rect 3876 19552 3892 19616
rect 3956 19552 3972 19616
rect 4036 19552 4042 19616
rect 3646 19551 4042 19552
rect 11646 19616 12042 19617
rect 11646 19552 11652 19616
rect 11716 19552 11732 19616
rect 11796 19552 11812 19616
rect 11876 19552 11892 19616
rect 11956 19552 11972 19616
rect 12036 19552 12042 19616
rect 11646 19551 12042 19552
rect 19646 19616 20042 19617
rect 19646 19552 19652 19616
rect 19716 19552 19732 19616
rect 19796 19552 19812 19616
rect 19876 19552 19892 19616
rect 19956 19552 19972 19616
rect 20036 19552 20042 19616
rect 19646 19551 20042 19552
rect 27646 19616 28042 19617
rect 27646 19552 27652 19616
rect 27716 19552 27732 19616
rect 27796 19552 27812 19616
rect 27876 19552 27892 19616
rect 27956 19552 27972 19616
rect 28036 19552 28042 19616
rect 27646 19551 28042 19552
rect 28349 19410 28415 19413
rect 29200 19410 30000 19440
rect 28349 19408 30000 19410
rect 28349 19352 28354 19408
rect 28410 19352 30000 19408
rect 28349 19350 30000 19352
rect 28349 19347 28415 19350
rect 29200 19320 30000 19350
rect 2906 19072 3302 19073
rect 2906 19008 2912 19072
rect 2976 19008 2992 19072
rect 3056 19008 3072 19072
rect 3136 19008 3152 19072
rect 3216 19008 3232 19072
rect 3296 19008 3302 19072
rect 2906 19007 3302 19008
rect 10906 19072 11302 19073
rect 10906 19008 10912 19072
rect 10976 19008 10992 19072
rect 11056 19008 11072 19072
rect 11136 19008 11152 19072
rect 11216 19008 11232 19072
rect 11296 19008 11302 19072
rect 10906 19007 11302 19008
rect 18906 19072 19302 19073
rect 18906 19008 18912 19072
rect 18976 19008 18992 19072
rect 19056 19008 19072 19072
rect 19136 19008 19152 19072
rect 19216 19008 19232 19072
rect 19296 19008 19302 19072
rect 18906 19007 19302 19008
rect 26906 19072 27302 19073
rect 26906 19008 26912 19072
rect 26976 19008 26992 19072
rect 27056 19008 27072 19072
rect 27136 19008 27152 19072
rect 27216 19008 27232 19072
rect 27296 19008 27302 19072
rect 26906 19007 27302 19008
rect 841 19002 907 19005
rect 798 19000 907 19002
rect 798 18944 846 19000
rect 902 18944 907 19000
rect 798 18939 907 18944
rect 798 18896 858 18939
rect 0 18806 858 18896
rect 0 18776 800 18806
rect 28349 18594 28415 18597
rect 29200 18594 30000 18624
rect 28349 18592 30000 18594
rect 28349 18536 28354 18592
rect 28410 18536 30000 18592
rect 28349 18534 30000 18536
rect 28349 18531 28415 18534
rect 3646 18528 4042 18529
rect 3646 18464 3652 18528
rect 3716 18464 3732 18528
rect 3796 18464 3812 18528
rect 3876 18464 3892 18528
rect 3956 18464 3972 18528
rect 4036 18464 4042 18528
rect 3646 18463 4042 18464
rect 11646 18528 12042 18529
rect 11646 18464 11652 18528
rect 11716 18464 11732 18528
rect 11796 18464 11812 18528
rect 11876 18464 11892 18528
rect 11956 18464 11972 18528
rect 12036 18464 12042 18528
rect 11646 18463 12042 18464
rect 19646 18528 20042 18529
rect 19646 18464 19652 18528
rect 19716 18464 19732 18528
rect 19796 18464 19812 18528
rect 19876 18464 19892 18528
rect 19956 18464 19972 18528
rect 20036 18464 20042 18528
rect 19646 18463 20042 18464
rect 27646 18528 28042 18529
rect 27646 18464 27652 18528
rect 27716 18464 27732 18528
rect 27796 18464 27812 18528
rect 27876 18464 27892 18528
rect 27956 18464 27972 18528
rect 28036 18464 28042 18528
rect 29200 18504 30000 18534
rect 27646 18463 28042 18464
rect 0 18050 800 18080
rect 1393 18050 1459 18053
rect 0 18048 1459 18050
rect 0 17992 1398 18048
rect 1454 17992 1459 18048
rect 0 17990 1459 17992
rect 0 17960 800 17990
rect 1393 17987 1459 17990
rect 2906 17984 3302 17985
rect 2906 17920 2912 17984
rect 2976 17920 2992 17984
rect 3056 17920 3072 17984
rect 3136 17920 3152 17984
rect 3216 17920 3232 17984
rect 3296 17920 3302 17984
rect 2906 17919 3302 17920
rect 10906 17984 11302 17985
rect 10906 17920 10912 17984
rect 10976 17920 10992 17984
rect 11056 17920 11072 17984
rect 11136 17920 11152 17984
rect 11216 17920 11232 17984
rect 11296 17920 11302 17984
rect 10906 17919 11302 17920
rect 18906 17984 19302 17985
rect 18906 17920 18912 17984
rect 18976 17920 18992 17984
rect 19056 17920 19072 17984
rect 19136 17920 19152 17984
rect 19216 17920 19232 17984
rect 19296 17920 19302 17984
rect 18906 17919 19302 17920
rect 26906 17984 27302 17985
rect 26906 17920 26912 17984
rect 26976 17920 26992 17984
rect 27056 17920 27072 17984
rect 27136 17920 27152 17984
rect 27216 17920 27232 17984
rect 27296 17920 27302 17984
rect 26906 17919 27302 17920
rect 28349 17778 28415 17781
rect 29200 17778 30000 17808
rect 28349 17776 30000 17778
rect 28349 17720 28354 17776
rect 28410 17720 30000 17776
rect 28349 17718 30000 17720
rect 28349 17715 28415 17718
rect 29200 17688 30000 17718
rect 3646 17440 4042 17441
rect 3646 17376 3652 17440
rect 3716 17376 3732 17440
rect 3796 17376 3812 17440
rect 3876 17376 3892 17440
rect 3956 17376 3972 17440
rect 4036 17376 4042 17440
rect 3646 17375 4042 17376
rect 11646 17440 12042 17441
rect 11646 17376 11652 17440
rect 11716 17376 11732 17440
rect 11796 17376 11812 17440
rect 11876 17376 11892 17440
rect 11956 17376 11972 17440
rect 12036 17376 12042 17440
rect 11646 17375 12042 17376
rect 19646 17440 20042 17441
rect 19646 17376 19652 17440
rect 19716 17376 19732 17440
rect 19796 17376 19812 17440
rect 19876 17376 19892 17440
rect 19956 17376 19972 17440
rect 20036 17376 20042 17440
rect 19646 17375 20042 17376
rect 27646 17440 28042 17441
rect 27646 17376 27652 17440
rect 27716 17376 27732 17440
rect 27796 17376 27812 17440
rect 27876 17376 27892 17440
rect 27956 17376 27972 17440
rect 28036 17376 28042 17440
rect 27646 17375 28042 17376
rect 1393 17370 1459 17373
rect 798 17368 1459 17370
rect 798 17312 1398 17368
rect 1454 17312 1459 17368
rect 798 17310 1459 17312
rect 798 17264 858 17310
rect 1393 17307 1459 17310
rect 0 17174 858 17264
rect 0 17144 800 17174
rect 28349 16962 28415 16965
rect 29200 16962 30000 16992
rect 28349 16960 30000 16962
rect 28349 16904 28354 16960
rect 28410 16904 30000 16960
rect 28349 16902 30000 16904
rect 28349 16899 28415 16902
rect 2906 16896 3302 16897
rect 2906 16832 2912 16896
rect 2976 16832 2992 16896
rect 3056 16832 3072 16896
rect 3136 16832 3152 16896
rect 3216 16832 3232 16896
rect 3296 16832 3302 16896
rect 2906 16831 3302 16832
rect 10906 16896 11302 16897
rect 10906 16832 10912 16896
rect 10976 16832 10992 16896
rect 11056 16832 11072 16896
rect 11136 16832 11152 16896
rect 11216 16832 11232 16896
rect 11296 16832 11302 16896
rect 10906 16831 11302 16832
rect 18906 16896 19302 16897
rect 18906 16832 18912 16896
rect 18976 16832 18992 16896
rect 19056 16832 19072 16896
rect 19136 16832 19152 16896
rect 19216 16832 19232 16896
rect 19296 16832 19302 16896
rect 18906 16831 19302 16832
rect 26906 16896 27302 16897
rect 26906 16832 26912 16896
rect 26976 16832 26992 16896
rect 27056 16832 27072 16896
rect 27136 16832 27152 16896
rect 27216 16832 27232 16896
rect 27296 16832 27302 16896
rect 29200 16872 30000 16902
rect 26906 16831 27302 16832
rect 1393 16554 1459 16557
rect 798 16552 1459 16554
rect 798 16496 1398 16552
rect 1454 16496 1459 16552
rect 798 16494 1459 16496
rect 798 16448 858 16494
rect 1393 16491 1459 16494
rect 0 16358 858 16448
rect 0 16328 800 16358
rect 3646 16352 4042 16353
rect 3646 16288 3652 16352
rect 3716 16288 3732 16352
rect 3796 16288 3812 16352
rect 3876 16288 3892 16352
rect 3956 16288 3972 16352
rect 4036 16288 4042 16352
rect 3646 16287 4042 16288
rect 11646 16352 12042 16353
rect 11646 16288 11652 16352
rect 11716 16288 11732 16352
rect 11796 16288 11812 16352
rect 11876 16288 11892 16352
rect 11956 16288 11972 16352
rect 12036 16288 12042 16352
rect 11646 16287 12042 16288
rect 19646 16352 20042 16353
rect 19646 16288 19652 16352
rect 19716 16288 19732 16352
rect 19796 16288 19812 16352
rect 19876 16288 19892 16352
rect 19956 16288 19972 16352
rect 20036 16288 20042 16352
rect 19646 16287 20042 16288
rect 27646 16352 28042 16353
rect 27646 16288 27652 16352
rect 27716 16288 27732 16352
rect 27796 16288 27812 16352
rect 27876 16288 27892 16352
rect 27956 16288 27972 16352
rect 28036 16288 28042 16352
rect 27646 16287 28042 16288
rect 28349 16146 28415 16149
rect 29200 16146 30000 16176
rect 28349 16144 30000 16146
rect 28349 16088 28354 16144
rect 28410 16088 30000 16144
rect 28349 16086 30000 16088
rect 28349 16083 28415 16086
rect 29200 16056 30000 16086
rect 2906 15808 3302 15809
rect 2906 15744 2912 15808
rect 2976 15744 2992 15808
rect 3056 15744 3072 15808
rect 3136 15744 3152 15808
rect 3216 15744 3232 15808
rect 3296 15744 3302 15808
rect 2906 15743 3302 15744
rect 10906 15808 11302 15809
rect 10906 15744 10912 15808
rect 10976 15744 10992 15808
rect 11056 15744 11072 15808
rect 11136 15744 11152 15808
rect 11216 15744 11232 15808
rect 11296 15744 11302 15808
rect 10906 15743 11302 15744
rect 18906 15808 19302 15809
rect 18906 15744 18912 15808
rect 18976 15744 18992 15808
rect 19056 15744 19072 15808
rect 19136 15744 19152 15808
rect 19216 15744 19232 15808
rect 19296 15744 19302 15808
rect 18906 15743 19302 15744
rect 26906 15808 27302 15809
rect 26906 15744 26912 15808
rect 26976 15744 26992 15808
rect 27056 15744 27072 15808
rect 27136 15744 27152 15808
rect 27216 15744 27232 15808
rect 27296 15744 27302 15808
rect 26906 15743 27302 15744
rect 1393 15738 1459 15741
rect 798 15736 1459 15738
rect 798 15680 1398 15736
rect 1454 15680 1459 15736
rect 798 15678 1459 15680
rect 798 15632 858 15678
rect 1393 15675 1459 15678
rect 0 15542 858 15632
rect 0 15512 800 15542
rect 11462 15404 11468 15468
rect 11532 15466 11538 15468
rect 11605 15466 11671 15469
rect 11532 15464 11671 15466
rect 11532 15408 11610 15464
rect 11666 15408 11671 15464
rect 11532 15406 11671 15408
rect 11532 15404 11538 15406
rect 11605 15403 11671 15406
rect 28349 15330 28415 15333
rect 29200 15330 30000 15360
rect 28349 15328 30000 15330
rect 28349 15272 28354 15328
rect 28410 15272 30000 15328
rect 28349 15270 30000 15272
rect 28349 15267 28415 15270
rect 3646 15264 4042 15265
rect 3646 15200 3652 15264
rect 3716 15200 3732 15264
rect 3796 15200 3812 15264
rect 3876 15200 3892 15264
rect 3956 15200 3972 15264
rect 4036 15200 4042 15264
rect 3646 15199 4042 15200
rect 11646 15264 12042 15265
rect 11646 15200 11652 15264
rect 11716 15200 11732 15264
rect 11796 15200 11812 15264
rect 11876 15200 11892 15264
rect 11956 15200 11972 15264
rect 12036 15200 12042 15264
rect 11646 15199 12042 15200
rect 19646 15264 20042 15265
rect 19646 15200 19652 15264
rect 19716 15200 19732 15264
rect 19796 15200 19812 15264
rect 19876 15200 19892 15264
rect 19956 15200 19972 15264
rect 20036 15200 20042 15264
rect 19646 15199 20042 15200
rect 27646 15264 28042 15265
rect 27646 15200 27652 15264
rect 27716 15200 27732 15264
rect 27796 15200 27812 15264
rect 27876 15200 27892 15264
rect 27956 15200 27972 15264
rect 28036 15200 28042 15264
rect 29200 15240 30000 15270
rect 27646 15199 28042 15200
rect 1393 14922 1459 14925
rect 798 14920 1459 14922
rect 798 14864 1398 14920
rect 1454 14864 1459 14920
rect 798 14862 1459 14864
rect 798 14816 858 14862
rect 1393 14859 1459 14862
rect 0 14726 858 14816
rect 0 14696 800 14726
rect 2906 14720 3302 14721
rect 2906 14656 2912 14720
rect 2976 14656 2992 14720
rect 3056 14656 3072 14720
rect 3136 14656 3152 14720
rect 3216 14656 3232 14720
rect 3296 14656 3302 14720
rect 2906 14655 3302 14656
rect 10906 14720 11302 14721
rect 10906 14656 10912 14720
rect 10976 14656 10992 14720
rect 11056 14656 11072 14720
rect 11136 14656 11152 14720
rect 11216 14656 11232 14720
rect 11296 14656 11302 14720
rect 10906 14655 11302 14656
rect 18906 14720 19302 14721
rect 18906 14656 18912 14720
rect 18976 14656 18992 14720
rect 19056 14656 19072 14720
rect 19136 14656 19152 14720
rect 19216 14656 19232 14720
rect 19296 14656 19302 14720
rect 18906 14655 19302 14656
rect 26906 14720 27302 14721
rect 26906 14656 26912 14720
rect 26976 14656 26992 14720
rect 27056 14656 27072 14720
rect 27136 14656 27152 14720
rect 27216 14656 27232 14720
rect 27296 14656 27302 14720
rect 26906 14655 27302 14656
rect 28349 14514 28415 14517
rect 29200 14514 30000 14544
rect 28349 14512 30000 14514
rect 28349 14456 28354 14512
rect 28410 14456 30000 14512
rect 28349 14454 30000 14456
rect 28349 14451 28415 14454
rect 29200 14424 30000 14454
rect 3646 14176 4042 14177
rect 3646 14112 3652 14176
rect 3716 14112 3732 14176
rect 3796 14112 3812 14176
rect 3876 14112 3892 14176
rect 3956 14112 3972 14176
rect 4036 14112 4042 14176
rect 3646 14111 4042 14112
rect 11646 14176 12042 14177
rect 11646 14112 11652 14176
rect 11716 14112 11732 14176
rect 11796 14112 11812 14176
rect 11876 14112 11892 14176
rect 11956 14112 11972 14176
rect 12036 14112 12042 14176
rect 11646 14111 12042 14112
rect 19646 14176 20042 14177
rect 19646 14112 19652 14176
rect 19716 14112 19732 14176
rect 19796 14112 19812 14176
rect 19876 14112 19892 14176
rect 19956 14112 19972 14176
rect 20036 14112 20042 14176
rect 19646 14111 20042 14112
rect 27646 14176 28042 14177
rect 27646 14112 27652 14176
rect 27716 14112 27732 14176
rect 27796 14112 27812 14176
rect 27876 14112 27892 14176
rect 27956 14112 27972 14176
rect 28036 14112 28042 14176
rect 27646 14111 28042 14112
rect 1393 14106 1459 14109
rect 798 14104 1459 14106
rect 798 14048 1398 14104
rect 1454 14048 1459 14104
rect 798 14046 1459 14048
rect 798 14000 858 14046
rect 1393 14043 1459 14046
rect 0 13910 858 14000
rect 0 13880 800 13910
rect 28349 13698 28415 13701
rect 29200 13698 30000 13728
rect 28349 13696 30000 13698
rect 28349 13640 28354 13696
rect 28410 13640 30000 13696
rect 28349 13638 30000 13640
rect 28349 13635 28415 13638
rect 2906 13632 3302 13633
rect 2906 13568 2912 13632
rect 2976 13568 2992 13632
rect 3056 13568 3072 13632
rect 3136 13568 3152 13632
rect 3216 13568 3232 13632
rect 3296 13568 3302 13632
rect 2906 13567 3302 13568
rect 10906 13632 11302 13633
rect 10906 13568 10912 13632
rect 10976 13568 10992 13632
rect 11056 13568 11072 13632
rect 11136 13568 11152 13632
rect 11216 13568 11232 13632
rect 11296 13568 11302 13632
rect 10906 13567 11302 13568
rect 18906 13632 19302 13633
rect 18906 13568 18912 13632
rect 18976 13568 18992 13632
rect 19056 13568 19072 13632
rect 19136 13568 19152 13632
rect 19216 13568 19232 13632
rect 19296 13568 19302 13632
rect 18906 13567 19302 13568
rect 26906 13632 27302 13633
rect 26906 13568 26912 13632
rect 26976 13568 26992 13632
rect 27056 13568 27072 13632
rect 27136 13568 27152 13632
rect 27216 13568 27232 13632
rect 27296 13568 27302 13632
rect 29200 13608 30000 13638
rect 26906 13567 27302 13568
rect 1393 13290 1459 13293
rect 798 13288 1459 13290
rect 798 13232 1398 13288
rect 1454 13232 1459 13288
rect 798 13230 1459 13232
rect 798 13184 858 13230
rect 1393 13227 1459 13230
rect 0 13094 858 13184
rect 0 13064 800 13094
rect 3646 13088 4042 13089
rect 3646 13024 3652 13088
rect 3716 13024 3732 13088
rect 3796 13024 3812 13088
rect 3876 13024 3892 13088
rect 3956 13024 3972 13088
rect 4036 13024 4042 13088
rect 3646 13023 4042 13024
rect 11646 13088 12042 13089
rect 11646 13024 11652 13088
rect 11716 13024 11732 13088
rect 11796 13024 11812 13088
rect 11876 13024 11892 13088
rect 11956 13024 11972 13088
rect 12036 13024 12042 13088
rect 11646 13023 12042 13024
rect 19646 13088 20042 13089
rect 19646 13024 19652 13088
rect 19716 13024 19732 13088
rect 19796 13024 19812 13088
rect 19876 13024 19892 13088
rect 19956 13024 19972 13088
rect 20036 13024 20042 13088
rect 19646 13023 20042 13024
rect 27646 13088 28042 13089
rect 27646 13024 27652 13088
rect 27716 13024 27732 13088
rect 27796 13024 27812 13088
rect 27876 13024 27892 13088
rect 27956 13024 27972 13088
rect 28036 13024 28042 13088
rect 27646 13023 28042 13024
rect 28349 12882 28415 12885
rect 29200 12882 30000 12912
rect 28349 12880 30000 12882
rect 28349 12824 28354 12880
rect 28410 12824 30000 12880
rect 28349 12822 30000 12824
rect 28349 12819 28415 12822
rect 29200 12792 30000 12822
rect 2906 12544 3302 12545
rect 2906 12480 2912 12544
rect 2976 12480 2992 12544
rect 3056 12480 3072 12544
rect 3136 12480 3152 12544
rect 3216 12480 3232 12544
rect 3296 12480 3302 12544
rect 2906 12479 3302 12480
rect 10906 12544 11302 12545
rect 10906 12480 10912 12544
rect 10976 12480 10992 12544
rect 11056 12480 11072 12544
rect 11136 12480 11152 12544
rect 11216 12480 11232 12544
rect 11296 12480 11302 12544
rect 10906 12479 11302 12480
rect 18906 12544 19302 12545
rect 18906 12480 18912 12544
rect 18976 12480 18992 12544
rect 19056 12480 19072 12544
rect 19136 12480 19152 12544
rect 19216 12480 19232 12544
rect 19296 12480 19302 12544
rect 18906 12479 19302 12480
rect 26906 12544 27302 12545
rect 26906 12480 26912 12544
rect 26976 12480 26992 12544
rect 27056 12480 27072 12544
rect 27136 12480 27152 12544
rect 27216 12480 27232 12544
rect 27296 12480 27302 12544
rect 26906 12479 27302 12480
rect 1393 12474 1459 12477
rect 798 12472 1459 12474
rect 798 12416 1398 12472
rect 1454 12416 1459 12472
rect 798 12414 1459 12416
rect 798 12368 858 12414
rect 1393 12411 1459 12414
rect 0 12278 858 12368
rect 0 12248 800 12278
rect 28349 12066 28415 12069
rect 29200 12066 30000 12096
rect 28349 12064 30000 12066
rect 28349 12008 28354 12064
rect 28410 12008 30000 12064
rect 28349 12006 30000 12008
rect 28349 12003 28415 12006
rect 3646 12000 4042 12001
rect 3646 11936 3652 12000
rect 3716 11936 3732 12000
rect 3796 11936 3812 12000
rect 3876 11936 3892 12000
rect 3956 11936 3972 12000
rect 4036 11936 4042 12000
rect 3646 11935 4042 11936
rect 11646 12000 12042 12001
rect 11646 11936 11652 12000
rect 11716 11936 11732 12000
rect 11796 11936 11812 12000
rect 11876 11936 11892 12000
rect 11956 11936 11972 12000
rect 12036 11936 12042 12000
rect 11646 11935 12042 11936
rect 19646 12000 20042 12001
rect 19646 11936 19652 12000
rect 19716 11936 19732 12000
rect 19796 11936 19812 12000
rect 19876 11936 19892 12000
rect 19956 11936 19972 12000
rect 20036 11936 20042 12000
rect 19646 11935 20042 11936
rect 27646 12000 28042 12001
rect 27646 11936 27652 12000
rect 27716 11936 27732 12000
rect 27796 11936 27812 12000
rect 27876 11936 27892 12000
rect 27956 11936 27972 12000
rect 28036 11936 28042 12000
rect 29200 11976 30000 12006
rect 27646 11935 28042 11936
rect 1393 11658 1459 11661
rect 798 11656 1459 11658
rect 798 11600 1398 11656
rect 1454 11600 1459 11656
rect 798 11598 1459 11600
rect 798 11552 858 11598
rect 1393 11595 1459 11598
rect 0 11462 858 11552
rect 0 11432 800 11462
rect 2906 11456 3302 11457
rect 2906 11392 2912 11456
rect 2976 11392 2992 11456
rect 3056 11392 3072 11456
rect 3136 11392 3152 11456
rect 3216 11392 3232 11456
rect 3296 11392 3302 11456
rect 2906 11391 3302 11392
rect 10906 11456 11302 11457
rect 10906 11392 10912 11456
rect 10976 11392 10992 11456
rect 11056 11392 11072 11456
rect 11136 11392 11152 11456
rect 11216 11392 11232 11456
rect 11296 11392 11302 11456
rect 10906 11391 11302 11392
rect 18906 11456 19302 11457
rect 18906 11392 18912 11456
rect 18976 11392 18992 11456
rect 19056 11392 19072 11456
rect 19136 11392 19152 11456
rect 19216 11392 19232 11456
rect 19296 11392 19302 11456
rect 18906 11391 19302 11392
rect 26906 11456 27302 11457
rect 26906 11392 26912 11456
rect 26976 11392 26992 11456
rect 27056 11392 27072 11456
rect 27136 11392 27152 11456
rect 27216 11392 27232 11456
rect 27296 11392 27302 11456
rect 26906 11391 27302 11392
rect 28349 11250 28415 11253
rect 29200 11250 30000 11280
rect 28349 11248 30000 11250
rect 28349 11192 28354 11248
rect 28410 11192 30000 11248
rect 28349 11190 30000 11192
rect 28349 11187 28415 11190
rect 29200 11160 30000 11190
rect 3646 10912 4042 10913
rect 3646 10848 3652 10912
rect 3716 10848 3732 10912
rect 3796 10848 3812 10912
rect 3876 10848 3892 10912
rect 3956 10848 3972 10912
rect 4036 10848 4042 10912
rect 3646 10847 4042 10848
rect 11646 10912 12042 10913
rect 11646 10848 11652 10912
rect 11716 10848 11732 10912
rect 11796 10848 11812 10912
rect 11876 10848 11892 10912
rect 11956 10848 11972 10912
rect 12036 10848 12042 10912
rect 11646 10847 12042 10848
rect 19646 10912 20042 10913
rect 19646 10848 19652 10912
rect 19716 10848 19732 10912
rect 19796 10848 19812 10912
rect 19876 10848 19892 10912
rect 19956 10848 19972 10912
rect 20036 10848 20042 10912
rect 19646 10847 20042 10848
rect 27646 10912 28042 10913
rect 27646 10848 27652 10912
rect 27716 10848 27732 10912
rect 27796 10848 27812 10912
rect 27876 10848 27892 10912
rect 27956 10848 27972 10912
rect 28036 10848 28042 10912
rect 27646 10847 28042 10848
rect 1393 10842 1459 10845
rect 798 10840 1459 10842
rect 798 10784 1398 10840
rect 1454 10784 1459 10840
rect 798 10782 1459 10784
rect 798 10736 858 10782
rect 1393 10779 1459 10782
rect 0 10646 858 10736
rect 0 10616 800 10646
rect 11513 10436 11579 10437
rect 11462 10372 11468 10436
rect 11532 10434 11579 10436
rect 28349 10434 28415 10437
rect 29200 10434 30000 10464
rect 11532 10432 11624 10434
rect 11574 10376 11624 10432
rect 11532 10374 11624 10376
rect 28349 10432 30000 10434
rect 28349 10376 28354 10432
rect 28410 10376 30000 10432
rect 28349 10374 30000 10376
rect 11532 10372 11579 10374
rect 11513 10371 11579 10372
rect 28349 10371 28415 10374
rect 2906 10368 3302 10369
rect 2906 10304 2912 10368
rect 2976 10304 2992 10368
rect 3056 10304 3072 10368
rect 3136 10304 3152 10368
rect 3216 10304 3232 10368
rect 3296 10304 3302 10368
rect 2906 10303 3302 10304
rect 10906 10368 11302 10369
rect 10906 10304 10912 10368
rect 10976 10304 10992 10368
rect 11056 10304 11072 10368
rect 11136 10304 11152 10368
rect 11216 10304 11232 10368
rect 11296 10304 11302 10368
rect 10906 10303 11302 10304
rect 18906 10368 19302 10369
rect 18906 10304 18912 10368
rect 18976 10304 18992 10368
rect 19056 10304 19072 10368
rect 19136 10304 19152 10368
rect 19216 10304 19232 10368
rect 19296 10304 19302 10368
rect 18906 10303 19302 10304
rect 26906 10368 27302 10369
rect 26906 10304 26912 10368
rect 26976 10304 26992 10368
rect 27056 10304 27072 10368
rect 27136 10304 27152 10368
rect 27216 10304 27232 10368
rect 27296 10304 27302 10368
rect 29200 10344 30000 10374
rect 26906 10303 27302 10304
rect 0 9890 800 9920
rect 1393 9890 1459 9893
rect 0 9888 1459 9890
rect 0 9832 1398 9888
rect 1454 9832 1459 9888
rect 0 9830 1459 9832
rect 0 9800 800 9830
rect 1393 9827 1459 9830
rect 3646 9824 4042 9825
rect 3646 9760 3652 9824
rect 3716 9760 3732 9824
rect 3796 9760 3812 9824
rect 3876 9760 3892 9824
rect 3956 9760 3972 9824
rect 4036 9760 4042 9824
rect 3646 9759 4042 9760
rect 11646 9824 12042 9825
rect 11646 9760 11652 9824
rect 11716 9760 11732 9824
rect 11796 9760 11812 9824
rect 11876 9760 11892 9824
rect 11956 9760 11972 9824
rect 12036 9760 12042 9824
rect 11646 9759 12042 9760
rect 19646 9824 20042 9825
rect 19646 9760 19652 9824
rect 19716 9760 19732 9824
rect 19796 9760 19812 9824
rect 19876 9760 19892 9824
rect 19956 9760 19972 9824
rect 20036 9760 20042 9824
rect 19646 9759 20042 9760
rect 27646 9824 28042 9825
rect 27646 9760 27652 9824
rect 27716 9760 27732 9824
rect 27796 9760 27812 9824
rect 27876 9760 27892 9824
rect 27956 9760 27972 9824
rect 28036 9760 28042 9824
rect 27646 9759 28042 9760
rect 28349 9618 28415 9621
rect 29200 9618 30000 9648
rect 28349 9616 30000 9618
rect 28349 9560 28354 9616
rect 28410 9560 30000 9616
rect 28349 9558 30000 9560
rect 28349 9555 28415 9558
rect 29200 9528 30000 9558
rect 2906 9280 3302 9281
rect 2906 9216 2912 9280
rect 2976 9216 2992 9280
rect 3056 9216 3072 9280
rect 3136 9216 3152 9280
rect 3216 9216 3232 9280
rect 3296 9216 3302 9280
rect 2906 9215 3302 9216
rect 10906 9280 11302 9281
rect 10906 9216 10912 9280
rect 10976 9216 10992 9280
rect 11056 9216 11072 9280
rect 11136 9216 11152 9280
rect 11216 9216 11232 9280
rect 11296 9216 11302 9280
rect 10906 9215 11302 9216
rect 18906 9280 19302 9281
rect 18906 9216 18912 9280
rect 18976 9216 18992 9280
rect 19056 9216 19072 9280
rect 19136 9216 19152 9280
rect 19216 9216 19232 9280
rect 19296 9216 19302 9280
rect 18906 9215 19302 9216
rect 26906 9280 27302 9281
rect 26906 9216 26912 9280
rect 26976 9216 26992 9280
rect 27056 9216 27072 9280
rect 27136 9216 27152 9280
rect 27216 9216 27232 9280
rect 27296 9216 27302 9280
rect 26906 9215 27302 9216
rect 1393 9210 1459 9213
rect 798 9208 1459 9210
rect 798 9152 1398 9208
rect 1454 9152 1459 9208
rect 798 9150 1459 9152
rect 798 9104 858 9150
rect 1393 9147 1459 9150
rect 0 9014 858 9104
rect 0 8984 800 9014
rect 28349 8802 28415 8805
rect 29200 8802 30000 8832
rect 28349 8800 30000 8802
rect 28349 8744 28354 8800
rect 28410 8744 30000 8800
rect 28349 8742 30000 8744
rect 28349 8739 28415 8742
rect 3646 8736 4042 8737
rect 3646 8672 3652 8736
rect 3716 8672 3732 8736
rect 3796 8672 3812 8736
rect 3876 8672 3892 8736
rect 3956 8672 3972 8736
rect 4036 8672 4042 8736
rect 3646 8671 4042 8672
rect 11646 8736 12042 8737
rect 11646 8672 11652 8736
rect 11716 8672 11732 8736
rect 11796 8672 11812 8736
rect 11876 8672 11892 8736
rect 11956 8672 11972 8736
rect 12036 8672 12042 8736
rect 11646 8671 12042 8672
rect 19646 8736 20042 8737
rect 19646 8672 19652 8736
rect 19716 8672 19732 8736
rect 19796 8672 19812 8736
rect 19876 8672 19892 8736
rect 19956 8672 19972 8736
rect 20036 8672 20042 8736
rect 19646 8671 20042 8672
rect 27646 8736 28042 8737
rect 27646 8672 27652 8736
rect 27716 8672 27732 8736
rect 27796 8672 27812 8736
rect 27876 8672 27892 8736
rect 27956 8672 27972 8736
rect 28036 8672 28042 8736
rect 29200 8712 30000 8742
rect 27646 8671 28042 8672
rect 1393 8394 1459 8397
rect 798 8392 1459 8394
rect 798 8336 1398 8392
rect 1454 8336 1459 8392
rect 798 8334 1459 8336
rect 798 8288 858 8334
rect 1393 8331 1459 8334
rect 0 8198 858 8288
rect 0 8168 800 8198
rect 2906 8192 3302 8193
rect 2906 8128 2912 8192
rect 2976 8128 2992 8192
rect 3056 8128 3072 8192
rect 3136 8128 3152 8192
rect 3216 8128 3232 8192
rect 3296 8128 3302 8192
rect 2906 8127 3302 8128
rect 10906 8192 11302 8193
rect 10906 8128 10912 8192
rect 10976 8128 10992 8192
rect 11056 8128 11072 8192
rect 11136 8128 11152 8192
rect 11216 8128 11232 8192
rect 11296 8128 11302 8192
rect 10906 8127 11302 8128
rect 18906 8192 19302 8193
rect 18906 8128 18912 8192
rect 18976 8128 18992 8192
rect 19056 8128 19072 8192
rect 19136 8128 19152 8192
rect 19216 8128 19232 8192
rect 19296 8128 19302 8192
rect 18906 8127 19302 8128
rect 26906 8192 27302 8193
rect 26906 8128 26912 8192
rect 26976 8128 26992 8192
rect 27056 8128 27072 8192
rect 27136 8128 27152 8192
rect 27216 8128 27232 8192
rect 27296 8128 27302 8192
rect 26906 8127 27302 8128
rect 28349 7986 28415 7989
rect 29200 7986 30000 8016
rect 28349 7984 30000 7986
rect 28349 7928 28354 7984
rect 28410 7928 30000 7984
rect 28349 7926 30000 7928
rect 28349 7923 28415 7926
rect 29200 7896 30000 7926
rect 3646 7648 4042 7649
rect 3646 7584 3652 7648
rect 3716 7584 3732 7648
rect 3796 7584 3812 7648
rect 3876 7584 3892 7648
rect 3956 7584 3972 7648
rect 4036 7584 4042 7648
rect 3646 7583 4042 7584
rect 11646 7648 12042 7649
rect 11646 7584 11652 7648
rect 11716 7584 11732 7648
rect 11796 7584 11812 7648
rect 11876 7584 11892 7648
rect 11956 7584 11972 7648
rect 12036 7584 12042 7648
rect 11646 7583 12042 7584
rect 19646 7648 20042 7649
rect 19646 7584 19652 7648
rect 19716 7584 19732 7648
rect 19796 7584 19812 7648
rect 19876 7584 19892 7648
rect 19956 7584 19972 7648
rect 20036 7584 20042 7648
rect 19646 7583 20042 7584
rect 27646 7648 28042 7649
rect 27646 7584 27652 7648
rect 27716 7584 27732 7648
rect 27796 7584 27812 7648
rect 27876 7584 27892 7648
rect 27956 7584 27972 7648
rect 28036 7584 28042 7648
rect 27646 7583 28042 7584
rect 1393 7578 1459 7581
rect 798 7576 1459 7578
rect 798 7520 1398 7576
rect 1454 7520 1459 7576
rect 798 7518 1459 7520
rect 798 7472 858 7518
rect 1393 7515 1459 7518
rect 0 7382 858 7472
rect 0 7352 800 7382
rect 28349 7170 28415 7173
rect 29200 7170 30000 7200
rect 28349 7168 30000 7170
rect 28349 7112 28354 7168
rect 28410 7112 30000 7168
rect 28349 7110 30000 7112
rect 28349 7107 28415 7110
rect 2906 7104 3302 7105
rect 2906 7040 2912 7104
rect 2976 7040 2992 7104
rect 3056 7040 3072 7104
rect 3136 7040 3152 7104
rect 3216 7040 3232 7104
rect 3296 7040 3302 7104
rect 2906 7039 3302 7040
rect 10906 7104 11302 7105
rect 10906 7040 10912 7104
rect 10976 7040 10992 7104
rect 11056 7040 11072 7104
rect 11136 7040 11152 7104
rect 11216 7040 11232 7104
rect 11296 7040 11302 7104
rect 10906 7039 11302 7040
rect 18906 7104 19302 7105
rect 18906 7040 18912 7104
rect 18976 7040 18992 7104
rect 19056 7040 19072 7104
rect 19136 7040 19152 7104
rect 19216 7040 19232 7104
rect 19296 7040 19302 7104
rect 18906 7039 19302 7040
rect 26906 7104 27302 7105
rect 26906 7040 26912 7104
rect 26976 7040 26992 7104
rect 27056 7040 27072 7104
rect 27136 7040 27152 7104
rect 27216 7040 27232 7104
rect 27296 7040 27302 7104
rect 29200 7080 30000 7110
rect 26906 7039 27302 7040
rect 0 6626 800 6656
rect 0 6536 858 6626
rect 798 6490 858 6536
rect 3646 6560 4042 6561
rect 3646 6496 3652 6560
rect 3716 6496 3732 6560
rect 3796 6496 3812 6560
rect 3876 6496 3892 6560
rect 3956 6496 3972 6560
rect 4036 6496 4042 6560
rect 3646 6495 4042 6496
rect 11646 6560 12042 6561
rect 11646 6496 11652 6560
rect 11716 6496 11732 6560
rect 11796 6496 11812 6560
rect 11876 6496 11892 6560
rect 11956 6496 11972 6560
rect 12036 6496 12042 6560
rect 11646 6495 12042 6496
rect 19646 6560 20042 6561
rect 19646 6496 19652 6560
rect 19716 6496 19732 6560
rect 19796 6496 19812 6560
rect 19876 6496 19892 6560
rect 19956 6496 19972 6560
rect 20036 6496 20042 6560
rect 19646 6495 20042 6496
rect 27646 6560 28042 6561
rect 27646 6496 27652 6560
rect 27716 6496 27732 6560
rect 27796 6496 27812 6560
rect 27876 6496 27892 6560
rect 27956 6496 27972 6560
rect 28036 6496 28042 6560
rect 27646 6495 28042 6496
rect 1393 6490 1459 6493
rect 798 6488 1459 6490
rect 798 6432 1398 6488
rect 1454 6432 1459 6488
rect 798 6430 1459 6432
rect 1393 6427 1459 6430
rect 28349 6354 28415 6357
rect 29200 6354 30000 6384
rect 28349 6352 30000 6354
rect 28349 6296 28354 6352
rect 28410 6296 30000 6352
rect 28349 6294 30000 6296
rect 28349 6291 28415 6294
rect 29200 6264 30000 6294
rect 2906 6016 3302 6017
rect 2906 5952 2912 6016
rect 2976 5952 2992 6016
rect 3056 5952 3072 6016
rect 3136 5952 3152 6016
rect 3216 5952 3232 6016
rect 3296 5952 3302 6016
rect 2906 5951 3302 5952
rect 10906 6016 11302 6017
rect 10906 5952 10912 6016
rect 10976 5952 10992 6016
rect 11056 5952 11072 6016
rect 11136 5952 11152 6016
rect 11216 5952 11232 6016
rect 11296 5952 11302 6016
rect 10906 5951 11302 5952
rect 18906 6016 19302 6017
rect 18906 5952 18912 6016
rect 18976 5952 18992 6016
rect 19056 5952 19072 6016
rect 19136 5952 19152 6016
rect 19216 5952 19232 6016
rect 19296 5952 19302 6016
rect 18906 5951 19302 5952
rect 26906 6016 27302 6017
rect 26906 5952 26912 6016
rect 26976 5952 26992 6016
rect 27056 5952 27072 6016
rect 27136 5952 27152 6016
rect 27216 5952 27232 6016
rect 27296 5952 27302 6016
rect 26906 5951 27302 5952
rect 1393 5946 1459 5949
rect 798 5944 1459 5946
rect 798 5888 1398 5944
rect 1454 5888 1459 5944
rect 798 5886 1459 5888
rect 798 5840 858 5886
rect 1393 5883 1459 5886
rect 0 5750 858 5840
rect 0 5720 800 5750
rect 28349 5538 28415 5541
rect 29200 5538 30000 5568
rect 28349 5536 30000 5538
rect 28349 5480 28354 5536
rect 28410 5480 30000 5536
rect 28349 5478 30000 5480
rect 28349 5475 28415 5478
rect 3646 5472 4042 5473
rect 3646 5408 3652 5472
rect 3716 5408 3732 5472
rect 3796 5408 3812 5472
rect 3876 5408 3892 5472
rect 3956 5408 3972 5472
rect 4036 5408 4042 5472
rect 3646 5407 4042 5408
rect 11646 5472 12042 5473
rect 11646 5408 11652 5472
rect 11716 5408 11732 5472
rect 11796 5408 11812 5472
rect 11876 5408 11892 5472
rect 11956 5408 11972 5472
rect 12036 5408 12042 5472
rect 11646 5407 12042 5408
rect 19646 5472 20042 5473
rect 19646 5408 19652 5472
rect 19716 5408 19732 5472
rect 19796 5408 19812 5472
rect 19876 5408 19892 5472
rect 19956 5408 19972 5472
rect 20036 5408 20042 5472
rect 19646 5407 20042 5408
rect 27646 5472 28042 5473
rect 27646 5408 27652 5472
rect 27716 5408 27732 5472
rect 27796 5408 27812 5472
rect 27876 5408 27892 5472
rect 27956 5408 27972 5472
rect 28036 5408 28042 5472
rect 29200 5448 30000 5478
rect 27646 5407 28042 5408
rect 790 5204 796 5268
rect 860 5266 866 5268
rect 1393 5266 1459 5269
rect 860 5264 1459 5266
rect 860 5208 1398 5264
rect 1454 5208 1459 5264
rect 860 5206 1459 5208
rect 860 5204 866 5206
rect 1393 5203 1459 5206
rect 0 4996 800 5024
rect 0 4932 796 4996
rect 860 4932 866 4996
rect 0 4904 800 4932
rect 2906 4928 3302 4929
rect 2906 4864 2912 4928
rect 2976 4864 2992 4928
rect 3056 4864 3072 4928
rect 3136 4864 3152 4928
rect 3216 4864 3232 4928
rect 3296 4864 3302 4928
rect 2906 4863 3302 4864
rect 10906 4928 11302 4929
rect 10906 4864 10912 4928
rect 10976 4864 10992 4928
rect 11056 4864 11072 4928
rect 11136 4864 11152 4928
rect 11216 4864 11232 4928
rect 11296 4864 11302 4928
rect 10906 4863 11302 4864
rect 18906 4928 19302 4929
rect 18906 4864 18912 4928
rect 18976 4864 18992 4928
rect 19056 4864 19072 4928
rect 19136 4864 19152 4928
rect 19216 4864 19232 4928
rect 19296 4864 19302 4928
rect 18906 4863 19302 4864
rect 26906 4928 27302 4929
rect 26906 4864 26912 4928
rect 26976 4864 26992 4928
rect 27056 4864 27072 4928
rect 27136 4864 27152 4928
rect 27216 4864 27232 4928
rect 27296 4864 27302 4928
rect 26906 4863 27302 4864
rect 28349 4722 28415 4725
rect 29200 4722 30000 4752
rect 28349 4720 30000 4722
rect 28349 4664 28354 4720
rect 28410 4664 30000 4720
rect 28349 4662 30000 4664
rect 28349 4659 28415 4662
rect 29200 4632 30000 4662
rect 3646 4384 4042 4385
rect 3646 4320 3652 4384
rect 3716 4320 3732 4384
rect 3796 4320 3812 4384
rect 3876 4320 3892 4384
rect 3956 4320 3972 4384
rect 4036 4320 4042 4384
rect 3646 4319 4042 4320
rect 11646 4384 12042 4385
rect 11646 4320 11652 4384
rect 11716 4320 11732 4384
rect 11796 4320 11812 4384
rect 11876 4320 11892 4384
rect 11956 4320 11972 4384
rect 12036 4320 12042 4384
rect 11646 4319 12042 4320
rect 19646 4384 20042 4385
rect 19646 4320 19652 4384
rect 19716 4320 19732 4384
rect 19796 4320 19812 4384
rect 19876 4320 19892 4384
rect 19956 4320 19972 4384
rect 20036 4320 20042 4384
rect 19646 4319 20042 4320
rect 27646 4384 28042 4385
rect 27646 4320 27652 4384
rect 27716 4320 27732 4384
rect 27796 4320 27812 4384
rect 27876 4320 27892 4384
rect 27956 4320 27972 4384
rect 28036 4320 28042 4384
rect 27646 4319 28042 4320
rect 1393 4314 1459 4317
rect 798 4312 1459 4314
rect 798 4256 1398 4312
rect 1454 4256 1459 4312
rect 798 4254 1459 4256
rect 798 4208 858 4254
rect 1393 4251 1459 4254
rect 0 4118 858 4208
rect 0 4088 800 4118
rect 28349 3906 28415 3909
rect 29200 3906 30000 3936
rect 28349 3904 30000 3906
rect 28349 3848 28354 3904
rect 28410 3848 30000 3904
rect 28349 3846 30000 3848
rect 28349 3843 28415 3846
rect 2906 3840 3302 3841
rect 2906 3776 2912 3840
rect 2976 3776 2992 3840
rect 3056 3776 3072 3840
rect 3136 3776 3152 3840
rect 3216 3776 3232 3840
rect 3296 3776 3302 3840
rect 2906 3775 3302 3776
rect 10906 3840 11302 3841
rect 10906 3776 10912 3840
rect 10976 3776 10992 3840
rect 11056 3776 11072 3840
rect 11136 3776 11152 3840
rect 11216 3776 11232 3840
rect 11296 3776 11302 3840
rect 10906 3775 11302 3776
rect 18906 3840 19302 3841
rect 18906 3776 18912 3840
rect 18976 3776 18992 3840
rect 19056 3776 19072 3840
rect 19136 3776 19152 3840
rect 19216 3776 19232 3840
rect 19296 3776 19302 3840
rect 18906 3775 19302 3776
rect 26906 3840 27302 3841
rect 26906 3776 26912 3840
rect 26976 3776 26992 3840
rect 27056 3776 27072 3840
rect 27136 3776 27152 3840
rect 27216 3776 27232 3840
rect 27296 3776 27302 3840
rect 29200 3816 30000 3846
rect 26906 3775 27302 3776
rect 1393 3498 1459 3501
rect 798 3496 1459 3498
rect 798 3440 1398 3496
rect 1454 3440 1459 3496
rect 798 3438 1459 3440
rect 798 3392 858 3438
rect 1393 3435 1459 3438
rect 0 3302 858 3392
rect 0 3272 800 3302
rect 3646 3296 4042 3297
rect 3646 3232 3652 3296
rect 3716 3232 3732 3296
rect 3796 3232 3812 3296
rect 3876 3232 3892 3296
rect 3956 3232 3972 3296
rect 4036 3232 4042 3296
rect 3646 3231 4042 3232
rect 11646 3296 12042 3297
rect 11646 3232 11652 3296
rect 11716 3232 11732 3296
rect 11796 3232 11812 3296
rect 11876 3232 11892 3296
rect 11956 3232 11972 3296
rect 12036 3232 12042 3296
rect 11646 3231 12042 3232
rect 19646 3296 20042 3297
rect 19646 3232 19652 3296
rect 19716 3232 19732 3296
rect 19796 3232 19812 3296
rect 19876 3232 19892 3296
rect 19956 3232 19972 3296
rect 20036 3232 20042 3296
rect 19646 3231 20042 3232
rect 27646 3296 28042 3297
rect 27646 3232 27652 3296
rect 27716 3232 27732 3296
rect 27796 3232 27812 3296
rect 27876 3232 27892 3296
rect 27956 3232 27972 3296
rect 28036 3232 28042 3296
rect 27646 3231 28042 3232
rect 28349 3090 28415 3093
rect 29200 3090 30000 3120
rect 28349 3088 30000 3090
rect 28349 3032 28354 3088
rect 28410 3032 30000 3088
rect 28349 3030 30000 3032
rect 28349 3027 28415 3030
rect 29200 3000 30000 3030
rect 2906 2752 3302 2753
rect 2906 2688 2912 2752
rect 2976 2688 2992 2752
rect 3056 2688 3072 2752
rect 3136 2688 3152 2752
rect 3216 2688 3232 2752
rect 3296 2688 3302 2752
rect 2906 2687 3302 2688
rect 10906 2752 11302 2753
rect 10906 2688 10912 2752
rect 10976 2688 10992 2752
rect 11056 2688 11072 2752
rect 11136 2688 11152 2752
rect 11216 2688 11232 2752
rect 11296 2688 11302 2752
rect 10906 2687 11302 2688
rect 18906 2752 19302 2753
rect 18906 2688 18912 2752
rect 18976 2688 18992 2752
rect 19056 2688 19072 2752
rect 19136 2688 19152 2752
rect 19216 2688 19232 2752
rect 19296 2688 19302 2752
rect 18906 2687 19302 2688
rect 26906 2752 27302 2753
rect 26906 2688 26912 2752
rect 26976 2688 26992 2752
rect 27056 2688 27072 2752
rect 27136 2688 27152 2752
rect 27216 2688 27232 2752
rect 27296 2688 27302 2752
rect 26906 2687 27302 2688
rect 841 2682 907 2685
rect 798 2680 907 2682
rect 798 2624 846 2680
rect 902 2624 907 2680
rect 798 2619 907 2624
rect 798 2576 858 2619
rect 0 2486 858 2576
rect 0 2456 800 2486
rect 28349 2274 28415 2277
rect 29200 2274 30000 2304
rect 28349 2272 30000 2274
rect 28349 2216 28354 2272
rect 28410 2216 30000 2272
rect 28349 2214 30000 2216
rect 28349 2211 28415 2214
rect 3646 2208 4042 2209
rect 3646 2144 3652 2208
rect 3716 2144 3732 2208
rect 3796 2144 3812 2208
rect 3876 2144 3892 2208
rect 3956 2144 3972 2208
rect 4036 2144 4042 2208
rect 3646 2143 4042 2144
rect 11646 2208 12042 2209
rect 11646 2144 11652 2208
rect 11716 2144 11732 2208
rect 11796 2144 11812 2208
rect 11876 2144 11892 2208
rect 11956 2144 11972 2208
rect 12036 2144 12042 2208
rect 11646 2143 12042 2144
rect 19646 2208 20042 2209
rect 19646 2144 19652 2208
rect 19716 2144 19732 2208
rect 19796 2144 19812 2208
rect 19876 2144 19892 2208
rect 19956 2144 19972 2208
rect 20036 2144 20042 2208
rect 19646 2143 20042 2144
rect 27646 2208 28042 2209
rect 27646 2144 27652 2208
rect 27716 2144 27732 2208
rect 27796 2144 27812 2208
rect 27876 2144 27892 2208
rect 27956 2144 27972 2208
rect 28036 2144 28042 2208
rect 29200 2184 30000 2214
rect 27646 2143 28042 2144
rect 841 1866 907 1869
rect 798 1864 907 1866
rect 798 1808 846 1864
rect 902 1808 907 1864
rect 798 1803 907 1808
rect 798 1760 858 1803
rect 0 1670 858 1760
rect 0 1640 800 1670
rect 105 1186 171 1189
rect 105 1184 1042 1186
rect 105 1128 110 1184
rect 166 1128 1042 1184
rect 105 1126 1042 1128
rect 105 1123 171 1126
rect 0 914 800 944
rect 982 914 1042 1126
rect 0 854 1042 914
rect 0 824 800 854
<< via3 >>
rect 2912 27772 2976 27776
rect 2912 27716 2916 27772
rect 2916 27716 2972 27772
rect 2972 27716 2976 27772
rect 2912 27712 2976 27716
rect 2992 27772 3056 27776
rect 2992 27716 2996 27772
rect 2996 27716 3052 27772
rect 3052 27716 3056 27772
rect 2992 27712 3056 27716
rect 3072 27772 3136 27776
rect 3072 27716 3076 27772
rect 3076 27716 3132 27772
rect 3132 27716 3136 27772
rect 3072 27712 3136 27716
rect 3152 27772 3216 27776
rect 3152 27716 3156 27772
rect 3156 27716 3212 27772
rect 3212 27716 3216 27772
rect 3152 27712 3216 27716
rect 3232 27772 3296 27776
rect 3232 27716 3236 27772
rect 3236 27716 3292 27772
rect 3292 27716 3296 27772
rect 3232 27712 3296 27716
rect 10912 27772 10976 27776
rect 10912 27716 10916 27772
rect 10916 27716 10972 27772
rect 10972 27716 10976 27772
rect 10912 27712 10976 27716
rect 10992 27772 11056 27776
rect 10992 27716 10996 27772
rect 10996 27716 11052 27772
rect 11052 27716 11056 27772
rect 10992 27712 11056 27716
rect 11072 27772 11136 27776
rect 11072 27716 11076 27772
rect 11076 27716 11132 27772
rect 11132 27716 11136 27772
rect 11072 27712 11136 27716
rect 11152 27772 11216 27776
rect 11152 27716 11156 27772
rect 11156 27716 11212 27772
rect 11212 27716 11216 27772
rect 11152 27712 11216 27716
rect 11232 27772 11296 27776
rect 11232 27716 11236 27772
rect 11236 27716 11292 27772
rect 11292 27716 11296 27772
rect 11232 27712 11296 27716
rect 18912 27772 18976 27776
rect 18912 27716 18916 27772
rect 18916 27716 18972 27772
rect 18972 27716 18976 27772
rect 18912 27712 18976 27716
rect 18992 27772 19056 27776
rect 18992 27716 18996 27772
rect 18996 27716 19052 27772
rect 19052 27716 19056 27772
rect 18992 27712 19056 27716
rect 19072 27772 19136 27776
rect 19072 27716 19076 27772
rect 19076 27716 19132 27772
rect 19132 27716 19136 27772
rect 19072 27712 19136 27716
rect 19152 27772 19216 27776
rect 19152 27716 19156 27772
rect 19156 27716 19212 27772
rect 19212 27716 19216 27772
rect 19152 27712 19216 27716
rect 19232 27772 19296 27776
rect 19232 27716 19236 27772
rect 19236 27716 19292 27772
rect 19292 27716 19296 27772
rect 19232 27712 19296 27716
rect 26912 27772 26976 27776
rect 26912 27716 26916 27772
rect 26916 27716 26972 27772
rect 26972 27716 26976 27772
rect 26912 27712 26976 27716
rect 26992 27772 27056 27776
rect 26992 27716 26996 27772
rect 26996 27716 27052 27772
rect 27052 27716 27056 27772
rect 26992 27712 27056 27716
rect 27072 27772 27136 27776
rect 27072 27716 27076 27772
rect 27076 27716 27132 27772
rect 27132 27716 27136 27772
rect 27072 27712 27136 27716
rect 27152 27772 27216 27776
rect 27152 27716 27156 27772
rect 27156 27716 27212 27772
rect 27212 27716 27216 27772
rect 27152 27712 27216 27716
rect 27232 27772 27296 27776
rect 27232 27716 27236 27772
rect 27236 27716 27292 27772
rect 27292 27716 27296 27772
rect 27232 27712 27296 27716
rect 3652 27228 3716 27232
rect 3652 27172 3656 27228
rect 3656 27172 3712 27228
rect 3712 27172 3716 27228
rect 3652 27168 3716 27172
rect 3732 27228 3796 27232
rect 3732 27172 3736 27228
rect 3736 27172 3792 27228
rect 3792 27172 3796 27228
rect 3732 27168 3796 27172
rect 3812 27228 3876 27232
rect 3812 27172 3816 27228
rect 3816 27172 3872 27228
rect 3872 27172 3876 27228
rect 3812 27168 3876 27172
rect 3892 27228 3956 27232
rect 3892 27172 3896 27228
rect 3896 27172 3952 27228
rect 3952 27172 3956 27228
rect 3892 27168 3956 27172
rect 3972 27228 4036 27232
rect 3972 27172 3976 27228
rect 3976 27172 4032 27228
rect 4032 27172 4036 27228
rect 3972 27168 4036 27172
rect 11652 27228 11716 27232
rect 11652 27172 11656 27228
rect 11656 27172 11712 27228
rect 11712 27172 11716 27228
rect 11652 27168 11716 27172
rect 11732 27228 11796 27232
rect 11732 27172 11736 27228
rect 11736 27172 11792 27228
rect 11792 27172 11796 27228
rect 11732 27168 11796 27172
rect 11812 27228 11876 27232
rect 11812 27172 11816 27228
rect 11816 27172 11872 27228
rect 11872 27172 11876 27228
rect 11812 27168 11876 27172
rect 11892 27228 11956 27232
rect 11892 27172 11896 27228
rect 11896 27172 11952 27228
rect 11952 27172 11956 27228
rect 11892 27168 11956 27172
rect 11972 27228 12036 27232
rect 11972 27172 11976 27228
rect 11976 27172 12032 27228
rect 12032 27172 12036 27228
rect 11972 27168 12036 27172
rect 19652 27228 19716 27232
rect 19652 27172 19656 27228
rect 19656 27172 19712 27228
rect 19712 27172 19716 27228
rect 19652 27168 19716 27172
rect 19732 27228 19796 27232
rect 19732 27172 19736 27228
rect 19736 27172 19792 27228
rect 19792 27172 19796 27228
rect 19732 27168 19796 27172
rect 19812 27228 19876 27232
rect 19812 27172 19816 27228
rect 19816 27172 19872 27228
rect 19872 27172 19876 27228
rect 19812 27168 19876 27172
rect 19892 27228 19956 27232
rect 19892 27172 19896 27228
rect 19896 27172 19952 27228
rect 19952 27172 19956 27228
rect 19892 27168 19956 27172
rect 19972 27228 20036 27232
rect 19972 27172 19976 27228
rect 19976 27172 20032 27228
rect 20032 27172 20036 27228
rect 19972 27168 20036 27172
rect 27652 27228 27716 27232
rect 27652 27172 27656 27228
rect 27656 27172 27712 27228
rect 27712 27172 27716 27228
rect 27652 27168 27716 27172
rect 27732 27228 27796 27232
rect 27732 27172 27736 27228
rect 27736 27172 27792 27228
rect 27792 27172 27796 27228
rect 27732 27168 27796 27172
rect 27812 27228 27876 27232
rect 27812 27172 27816 27228
rect 27816 27172 27872 27228
rect 27872 27172 27876 27228
rect 27812 27168 27876 27172
rect 27892 27228 27956 27232
rect 27892 27172 27896 27228
rect 27896 27172 27952 27228
rect 27952 27172 27956 27228
rect 27892 27168 27956 27172
rect 27972 27228 28036 27232
rect 27972 27172 27976 27228
rect 27976 27172 28032 27228
rect 28032 27172 28036 27228
rect 27972 27168 28036 27172
rect 2912 26684 2976 26688
rect 2912 26628 2916 26684
rect 2916 26628 2972 26684
rect 2972 26628 2976 26684
rect 2912 26624 2976 26628
rect 2992 26684 3056 26688
rect 2992 26628 2996 26684
rect 2996 26628 3052 26684
rect 3052 26628 3056 26684
rect 2992 26624 3056 26628
rect 3072 26684 3136 26688
rect 3072 26628 3076 26684
rect 3076 26628 3132 26684
rect 3132 26628 3136 26684
rect 3072 26624 3136 26628
rect 3152 26684 3216 26688
rect 3152 26628 3156 26684
rect 3156 26628 3212 26684
rect 3212 26628 3216 26684
rect 3152 26624 3216 26628
rect 3232 26684 3296 26688
rect 3232 26628 3236 26684
rect 3236 26628 3292 26684
rect 3292 26628 3296 26684
rect 3232 26624 3296 26628
rect 10912 26684 10976 26688
rect 10912 26628 10916 26684
rect 10916 26628 10972 26684
rect 10972 26628 10976 26684
rect 10912 26624 10976 26628
rect 10992 26684 11056 26688
rect 10992 26628 10996 26684
rect 10996 26628 11052 26684
rect 11052 26628 11056 26684
rect 10992 26624 11056 26628
rect 11072 26684 11136 26688
rect 11072 26628 11076 26684
rect 11076 26628 11132 26684
rect 11132 26628 11136 26684
rect 11072 26624 11136 26628
rect 11152 26684 11216 26688
rect 11152 26628 11156 26684
rect 11156 26628 11212 26684
rect 11212 26628 11216 26684
rect 11152 26624 11216 26628
rect 11232 26684 11296 26688
rect 11232 26628 11236 26684
rect 11236 26628 11292 26684
rect 11292 26628 11296 26684
rect 11232 26624 11296 26628
rect 18912 26684 18976 26688
rect 18912 26628 18916 26684
rect 18916 26628 18972 26684
rect 18972 26628 18976 26684
rect 18912 26624 18976 26628
rect 18992 26684 19056 26688
rect 18992 26628 18996 26684
rect 18996 26628 19052 26684
rect 19052 26628 19056 26684
rect 18992 26624 19056 26628
rect 19072 26684 19136 26688
rect 19072 26628 19076 26684
rect 19076 26628 19132 26684
rect 19132 26628 19136 26684
rect 19072 26624 19136 26628
rect 19152 26684 19216 26688
rect 19152 26628 19156 26684
rect 19156 26628 19212 26684
rect 19212 26628 19216 26684
rect 19152 26624 19216 26628
rect 19232 26684 19296 26688
rect 19232 26628 19236 26684
rect 19236 26628 19292 26684
rect 19292 26628 19296 26684
rect 19232 26624 19296 26628
rect 26912 26684 26976 26688
rect 26912 26628 26916 26684
rect 26916 26628 26972 26684
rect 26972 26628 26976 26684
rect 26912 26624 26976 26628
rect 26992 26684 27056 26688
rect 26992 26628 26996 26684
rect 26996 26628 27052 26684
rect 27052 26628 27056 26684
rect 26992 26624 27056 26628
rect 27072 26684 27136 26688
rect 27072 26628 27076 26684
rect 27076 26628 27132 26684
rect 27132 26628 27136 26684
rect 27072 26624 27136 26628
rect 27152 26684 27216 26688
rect 27152 26628 27156 26684
rect 27156 26628 27212 26684
rect 27212 26628 27216 26684
rect 27152 26624 27216 26628
rect 27232 26684 27296 26688
rect 27232 26628 27236 26684
rect 27236 26628 27292 26684
rect 27292 26628 27296 26684
rect 27232 26624 27296 26628
rect 3652 26140 3716 26144
rect 3652 26084 3656 26140
rect 3656 26084 3712 26140
rect 3712 26084 3716 26140
rect 3652 26080 3716 26084
rect 3732 26140 3796 26144
rect 3732 26084 3736 26140
rect 3736 26084 3792 26140
rect 3792 26084 3796 26140
rect 3732 26080 3796 26084
rect 3812 26140 3876 26144
rect 3812 26084 3816 26140
rect 3816 26084 3872 26140
rect 3872 26084 3876 26140
rect 3812 26080 3876 26084
rect 3892 26140 3956 26144
rect 3892 26084 3896 26140
rect 3896 26084 3952 26140
rect 3952 26084 3956 26140
rect 3892 26080 3956 26084
rect 3972 26140 4036 26144
rect 3972 26084 3976 26140
rect 3976 26084 4032 26140
rect 4032 26084 4036 26140
rect 3972 26080 4036 26084
rect 11652 26140 11716 26144
rect 11652 26084 11656 26140
rect 11656 26084 11712 26140
rect 11712 26084 11716 26140
rect 11652 26080 11716 26084
rect 11732 26140 11796 26144
rect 11732 26084 11736 26140
rect 11736 26084 11792 26140
rect 11792 26084 11796 26140
rect 11732 26080 11796 26084
rect 11812 26140 11876 26144
rect 11812 26084 11816 26140
rect 11816 26084 11872 26140
rect 11872 26084 11876 26140
rect 11812 26080 11876 26084
rect 11892 26140 11956 26144
rect 11892 26084 11896 26140
rect 11896 26084 11952 26140
rect 11952 26084 11956 26140
rect 11892 26080 11956 26084
rect 11972 26140 12036 26144
rect 11972 26084 11976 26140
rect 11976 26084 12032 26140
rect 12032 26084 12036 26140
rect 11972 26080 12036 26084
rect 19652 26140 19716 26144
rect 19652 26084 19656 26140
rect 19656 26084 19712 26140
rect 19712 26084 19716 26140
rect 19652 26080 19716 26084
rect 19732 26140 19796 26144
rect 19732 26084 19736 26140
rect 19736 26084 19792 26140
rect 19792 26084 19796 26140
rect 19732 26080 19796 26084
rect 19812 26140 19876 26144
rect 19812 26084 19816 26140
rect 19816 26084 19872 26140
rect 19872 26084 19876 26140
rect 19812 26080 19876 26084
rect 19892 26140 19956 26144
rect 19892 26084 19896 26140
rect 19896 26084 19952 26140
rect 19952 26084 19956 26140
rect 19892 26080 19956 26084
rect 19972 26140 20036 26144
rect 19972 26084 19976 26140
rect 19976 26084 20032 26140
rect 20032 26084 20036 26140
rect 19972 26080 20036 26084
rect 27652 26140 27716 26144
rect 27652 26084 27656 26140
rect 27656 26084 27712 26140
rect 27712 26084 27716 26140
rect 27652 26080 27716 26084
rect 27732 26140 27796 26144
rect 27732 26084 27736 26140
rect 27736 26084 27792 26140
rect 27792 26084 27796 26140
rect 27732 26080 27796 26084
rect 27812 26140 27876 26144
rect 27812 26084 27816 26140
rect 27816 26084 27872 26140
rect 27872 26084 27876 26140
rect 27812 26080 27876 26084
rect 27892 26140 27956 26144
rect 27892 26084 27896 26140
rect 27896 26084 27952 26140
rect 27952 26084 27956 26140
rect 27892 26080 27956 26084
rect 27972 26140 28036 26144
rect 27972 26084 27976 26140
rect 27976 26084 28032 26140
rect 28032 26084 28036 26140
rect 27972 26080 28036 26084
rect 2912 25596 2976 25600
rect 2912 25540 2916 25596
rect 2916 25540 2972 25596
rect 2972 25540 2976 25596
rect 2912 25536 2976 25540
rect 2992 25596 3056 25600
rect 2992 25540 2996 25596
rect 2996 25540 3052 25596
rect 3052 25540 3056 25596
rect 2992 25536 3056 25540
rect 3072 25596 3136 25600
rect 3072 25540 3076 25596
rect 3076 25540 3132 25596
rect 3132 25540 3136 25596
rect 3072 25536 3136 25540
rect 3152 25596 3216 25600
rect 3152 25540 3156 25596
rect 3156 25540 3212 25596
rect 3212 25540 3216 25596
rect 3152 25536 3216 25540
rect 3232 25596 3296 25600
rect 3232 25540 3236 25596
rect 3236 25540 3292 25596
rect 3292 25540 3296 25596
rect 3232 25536 3296 25540
rect 10912 25596 10976 25600
rect 10912 25540 10916 25596
rect 10916 25540 10972 25596
rect 10972 25540 10976 25596
rect 10912 25536 10976 25540
rect 10992 25596 11056 25600
rect 10992 25540 10996 25596
rect 10996 25540 11052 25596
rect 11052 25540 11056 25596
rect 10992 25536 11056 25540
rect 11072 25596 11136 25600
rect 11072 25540 11076 25596
rect 11076 25540 11132 25596
rect 11132 25540 11136 25596
rect 11072 25536 11136 25540
rect 11152 25596 11216 25600
rect 11152 25540 11156 25596
rect 11156 25540 11212 25596
rect 11212 25540 11216 25596
rect 11152 25536 11216 25540
rect 11232 25596 11296 25600
rect 11232 25540 11236 25596
rect 11236 25540 11292 25596
rect 11292 25540 11296 25596
rect 11232 25536 11296 25540
rect 18912 25596 18976 25600
rect 18912 25540 18916 25596
rect 18916 25540 18972 25596
rect 18972 25540 18976 25596
rect 18912 25536 18976 25540
rect 18992 25596 19056 25600
rect 18992 25540 18996 25596
rect 18996 25540 19052 25596
rect 19052 25540 19056 25596
rect 18992 25536 19056 25540
rect 19072 25596 19136 25600
rect 19072 25540 19076 25596
rect 19076 25540 19132 25596
rect 19132 25540 19136 25596
rect 19072 25536 19136 25540
rect 19152 25596 19216 25600
rect 19152 25540 19156 25596
rect 19156 25540 19212 25596
rect 19212 25540 19216 25596
rect 19152 25536 19216 25540
rect 19232 25596 19296 25600
rect 19232 25540 19236 25596
rect 19236 25540 19292 25596
rect 19292 25540 19296 25596
rect 19232 25536 19296 25540
rect 26912 25596 26976 25600
rect 26912 25540 26916 25596
rect 26916 25540 26972 25596
rect 26972 25540 26976 25596
rect 26912 25536 26976 25540
rect 26992 25596 27056 25600
rect 26992 25540 26996 25596
rect 26996 25540 27052 25596
rect 27052 25540 27056 25596
rect 26992 25536 27056 25540
rect 27072 25596 27136 25600
rect 27072 25540 27076 25596
rect 27076 25540 27132 25596
rect 27132 25540 27136 25596
rect 27072 25536 27136 25540
rect 27152 25596 27216 25600
rect 27152 25540 27156 25596
rect 27156 25540 27212 25596
rect 27212 25540 27216 25596
rect 27152 25536 27216 25540
rect 27232 25596 27296 25600
rect 27232 25540 27236 25596
rect 27236 25540 27292 25596
rect 27292 25540 27296 25596
rect 27232 25536 27296 25540
rect 3652 25052 3716 25056
rect 3652 24996 3656 25052
rect 3656 24996 3712 25052
rect 3712 24996 3716 25052
rect 3652 24992 3716 24996
rect 3732 25052 3796 25056
rect 3732 24996 3736 25052
rect 3736 24996 3792 25052
rect 3792 24996 3796 25052
rect 3732 24992 3796 24996
rect 3812 25052 3876 25056
rect 3812 24996 3816 25052
rect 3816 24996 3872 25052
rect 3872 24996 3876 25052
rect 3812 24992 3876 24996
rect 3892 25052 3956 25056
rect 3892 24996 3896 25052
rect 3896 24996 3952 25052
rect 3952 24996 3956 25052
rect 3892 24992 3956 24996
rect 3972 25052 4036 25056
rect 3972 24996 3976 25052
rect 3976 24996 4032 25052
rect 4032 24996 4036 25052
rect 3972 24992 4036 24996
rect 11652 25052 11716 25056
rect 11652 24996 11656 25052
rect 11656 24996 11712 25052
rect 11712 24996 11716 25052
rect 11652 24992 11716 24996
rect 11732 25052 11796 25056
rect 11732 24996 11736 25052
rect 11736 24996 11792 25052
rect 11792 24996 11796 25052
rect 11732 24992 11796 24996
rect 11812 25052 11876 25056
rect 11812 24996 11816 25052
rect 11816 24996 11872 25052
rect 11872 24996 11876 25052
rect 11812 24992 11876 24996
rect 11892 25052 11956 25056
rect 11892 24996 11896 25052
rect 11896 24996 11952 25052
rect 11952 24996 11956 25052
rect 11892 24992 11956 24996
rect 11972 25052 12036 25056
rect 11972 24996 11976 25052
rect 11976 24996 12032 25052
rect 12032 24996 12036 25052
rect 11972 24992 12036 24996
rect 19652 25052 19716 25056
rect 19652 24996 19656 25052
rect 19656 24996 19712 25052
rect 19712 24996 19716 25052
rect 19652 24992 19716 24996
rect 19732 25052 19796 25056
rect 19732 24996 19736 25052
rect 19736 24996 19792 25052
rect 19792 24996 19796 25052
rect 19732 24992 19796 24996
rect 19812 25052 19876 25056
rect 19812 24996 19816 25052
rect 19816 24996 19872 25052
rect 19872 24996 19876 25052
rect 19812 24992 19876 24996
rect 19892 25052 19956 25056
rect 19892 24996 19896 25052
rect 19896 24996 19952 25052
rect 19952 24996 19956 25052
rect 19892 24992 19956 24996
rect 19972 25052 20036 25056
rect 19972 24996 19976 25052
rect 19976 24996 20032 25052
rect 20032 24996 20036 25052
rect 19972 24992 20036 24996
rect 27652 25052 27716 25056
rect 27652 24996 27656 25052
rect 27656 24996 27712 25052
rect 27712 24996 27716 25052
rect 27652 24992 27716 24996
rect 27732 25052 27796 25056
rect 27732 24996 27736 25052
rect 27736 24996 27792 25052
rect 27792 24996 27796 25052
rect 27732 24992 27796 24996
rect 27812 25052 27876 25056
rect 27812 24996 27816 25052
rect 27816 24996 27872 25052
rect 27872 24996 27876 25052
rect 27812 24992 27876 24996
rect 27892 25052 27956 25056
rect 27892 24996 27896 25052
rect 27896 24996 27952 25052
rect 27952 24996 27956 25052
rect 27892 24992 27956 24996
rect 27972 25052 28036 25056
rect 27972 24996 27976 25052
rect 27976 24996 28032 25052
rect 28032 24996 28036 25052
rect 27972 24992 28036 24996
rect 2912 24508 2976 24512
rect 2912 24452 2916 24508
rect 2916 24452 2972 24508
rect 2972 24452 2976 24508
rect 2912 24448 2976 24452
rect 2992 24508 3056 24512
rect 2992 24452 2996 24508
rect 2996 24452 3052 24508
rect 3052 24452 3056 24508
rect 2992 24448 3056 24452
rect 3072 24508 3136 24512
rect 3072 24452 3076 24508
rect 3076 24452 3132 24508
rect 3132 24452 3136 24508
rect 3072 24448 3136 24452
rect 3152 24508 3216 24512
rect 3152 24452 3156 24508
rect 3156 24452 3212 24508
rect 3212 24452 3216 24508
rect 3152 24448 3216 24452
rect 3232 24508 3296 24512
rect 3232 24452 3236 24508
rect 3236 24452 3292 24508
rect 3292 24452 3296 24508
rect 3232 24448 3296 24452
rect 10912 24508 10976 24512
rect 10912 24452 10916 24508
rect 10916 24452 10972 24508
rect 10972 24452 10976 24508
rect 10912 24448 10976 24452
rect 10992 24508 11056 24512
rect 10992 24452 10996 24508
rect 10996 24452 11052 24508
rect 11052 24452 11056 24508
rect 10992 24448 11056 24452
rect 11072 24508 11136 24512
rect 11072 24452 11076 24508
rect 11076 24452 11132 24508
rect 11132 24452 11136 24508
rect 11072 24448 11136 24452
rect 11152 24508 11216 24512
rect 11152 24452 11156 24508
rect 11156 24452 11212 24508
rect 11212 24452 11216 24508
rect 11152 24448 11216 24452
rect 11232 24508 11296 24512
rect 11232 24452 11236 24508
rect 11236 24452 11292 24508
rect 11292 24452 11296 24508
rect 11232 24448 11296 24452
rect 18912 24508 18976 24512
rect 18912 24452 18916 24508
rect 18916 24452 18972 24508
rect 18972 24452 18976 24508
rect 18912 24448 18976 24452
rect 18992 24508 19056 24512
rect 18992 24452 18996 24508
rect 18996 24452 19052 24508
rect 19052 24452 19056 24508
rect 18992 24448 19056 24452
rect 19072 24508 19136 24512
rect 19072 24452 19076 24508
rect 19076 24452 19132 24508
rect 19132 24452 19136 24508
rect 19072 24448 19136 24452
rect 19152 24508 19216 24512
rect 19152 24452 19156 24508
rect 19156 24452 19212 24508
rect 19212 24452 19216 24508
rect 19152 24448 19216 24452
rect 19232 24508 19296 24512
rect 19232 24452 19236 24508
rect 19236 24452 19292 24508
rect 19292 24452 19296 24508
rect 19232 24448 19296 24452
rect 26912 24508 26976 24512
rect 26912 24452 26916 24508
rect 26916 24452 26972 24508
rect 26972 24452 26976 24508
rect 26912 24448 26976 24452
rect 26992 24508 27056 24512
rect 26992 24452 26996 24508
rect 26996 24452 27052 24508
rect 27052 24452 27056 24508
rect 26992 24448 27056 24452
rect 27072 24508 27136 24512
rect 27072 24452 27076 24508
rect 27076 24452 27132 24508
rect 27132 24452 27136 24508
rect 27072 24448 27136 24452
rect 27152 24508 27216 24512
rect 27152 24452 27156 24508
rect 27156 24452 27212 24508
rect 27212 24452 27216 24508
rect 27152 24448 27216 24452
rect 27232 24508 27296 24512
rect 27232 24452 27236 24508
rect 27236 24452 27292 24508
rect 27292 24452 27296 24508
rect 27232 24448 27296 24452
rect 3652 23964 3716 23968
rect 3652 23908 3656 23964
rect 3656 23908 3712 23964
rect 3712 23908 3716 23964
rect 3652 23904 3716 23908
rect 3732 23964 3796 23968
rect 3732 23908 3736 23964
rect 3736 23908 3792 23964
rect 3792 23908 3796 23964
rect 3732 23904 3796 23908
rect 3812 23964 3876 23968
rect 3812 23908 3816 23964
rect 3816 23908 3872 23964
rect 3872 23908 3876 23964
rect 3812 23904 3876 23908
rect 3892 23964 3956 23968
rect 3892 23908 3896 23964
rect 3896 23908 3952 23964
rect 3952 23908 3956 23964
rect 3892 23904 3956 23908
rect 3972 23964 4036 23968
rect 3972 23908 3976 23964
rect 3976 23908 4032 23964
rect 4032 23908 4036 23964
rect 3972 23904 4036 23908
rect 11652 23964 11716 23968
rect 11652 23908 11656 23964
rect 11656 23908 11712 23964
rect 11712 23908 11716 23964
rect 11652 23904 11716 23908
rect 11732 23964 11796 23968
rect 11732 23908 11736 23964
rect 11736 23908 11792 23964
rect 11792 23908 11796 23964
rect 11732 23904 11796 23908
rect 11812 23964 11876 23968
rect 11812 23908 11816 23964
rect 11816 23908 11872 23964
rect 11872 23908 11876 23964
rect 11812 23904 11876 23908
rect 11892 23964 11956 23968
rect 11892 23908 11896 23964
rect 11896 23908 11952 23964
rect 11952 23908 11956 23964
rect 11892 23904 11956 23908
rect 11972 23964 12036 23968
rect 11972 23908 11976 23964
rect 11976 23908 12032 23964
rect 12032 23908 12036 23964
rect 11972 23904 12036 23908
rect 19652 23964 19716 23968
rect 19652 23908 19656 23964
rect 19656 23908 19712 23964
rect 19712 23908 19716 23964
rect 19652 23904 19716 23908
rect 19732 23964 19796 23968
rect 19732 23908 19736 23964
rect 19736 23908 19792 23964
rect 19792 23908 19796 23964
rect 19732 23904 19796 23908
rect 19812 23964 19876 23968
rect 19812 23908 19816 23964
rect 19816 23908 19872 23964
rect 19872 23908 19876 23964
rect 19812 23904 19876 23908
rect 19892 23964 19956 23968
rect 19892 23908 19896 23964
rect 19896 23908 19952 23964
rect 19952 23908 19956 23964
rect 19892 23904 19956 23908
rect 19972 23964 20036 23968
rect 19972 23908 19976 23964
rect 19976 23908 20032 23964
rect 20032 23908 20036 23964
rect 19972 23904 20036 23908
rect 27652 23964 27716 23968
rect 27652 23908 27656 23964
rect 27656 23908 27712 23964
rect 27712 23908 27716 23964
rect 27652 23904 27716 23908
rect 27732 23964 27796 23968
rect 27732 23908 27736 23964
rect 27736 23908 27792 23964
rect 27792 23908 27796 23964
rect 27732 23904 27796 23908
rect 27812 23964 27876 23968
rect 27812 23908 27816 23964
rect 27816 23908 27872 23964
rect 27872 23908 27876 23964
rect 27812 23904 27876 23908
rect 27892 23964 27956 23968
rect 27892 23908 27896 23964
rect 27896 23908 27952 23964
rect 27952 23908 27956 23964
rect 27892 23904 27956 23908
rect 27972 23964 28036 23968
rect 27972 23908 27976 23964
rect 27976 23908 28032 23964
rect 28032 23908 28036 23964
rect 27972 23904 28036 23908
rect 2912 23420 2976 23424
rect 2912 23364 2916 23420
rect 2916 23364 2972 23420
rect 2972 23364 2976 23420
rect 2912 23360 2976 23364
rect 2992 23420 3056 23424
rect 2992 23364 2996 23420
rect 2996 23364 3052 23420
rect 3052 23364 3056 23420
rect 2992 23360 3056 23364
rect 3072 23420 3136 23424
rect 3072 23364 3076 23420
rect 3076 23364 3132 23420
rect 3132 23364 3136 23420
rect 3072 23360 3136 23364
rect 3152 23420 3216 23424
rect 3152 23364 3156 23420
rect 3156 23364 3212 23420
rect 3212 23364 3216 23420
rect 3152 23360 3216 23364
rect 3232 23420 3296 23424
rect 3232 23364 3236 23420
rect 3236 23364 3292 23420
rect 3292 23364 3296 23420
rect 3232 23360 3296 23364
rect 10912 23420 10976 23424
rect 10912 23364 10916 23420
rect 10916 23364 10972 23420
rect 10972 23364 10976 23420
rect 10912 23360 10976 23364
rect 10992 23420 11056 23424
rect 10992 23364 10996 23420
rect 10996 23364 11052 23420
rect 11052 23364 11056 23420
rect 10992 23360 11056 23364
rect 11072 23420 11136 23424
rect 11072 23364 11076 23420
rect 11076 23364 11132 23420
rect 11132 23364 11136 23420
rect 11072 23360 11136 23364
rect 11152 23420 11216 23424
rect 11152 23364 11156 23420
rect 11156 23364 11212 23420
rect 11212 23364 11216 23420
rect 11152 23360 11216 23364
rect 11232 23420 11296 23424
rect 11232 23364 11236 23420
rect 11236 23364 11292 23420
rect 11292 23364 11296 23420
rect 11232 23360 11296 23364
rect 18912 23420 18976 23424
rect 18912 23364 18916 23420
rect 18916 23364 18972 23420
rect 18972 23364 18976 23420
rect 18912 23360 18976 23364
rect 18992 23420 19056 23424
rect 18992 23364 18996 23420
rect 18996 23364 19052 23420
rect 19052 23364 19056 23420
rect 18992 23360 19056 23364
rect 19072 23420 19136 23424
rect 19072 23364 19076 23420
rect 19076 23364 19132 23420
rect 19132 23364 19136 23420
rect 19072 23360 19136 23364
rect 19152 23420 19216 23424
rect 19152 23364 19156 23420
rect 19156 23364 19212 23420
rect 19212 23364 19216 23420
rect 19152 23360 19216 23364
rect 19232 23420 19296 23424
rect 19232 23364 19236 23420
rect 19236 23364 19292 23420
rect 19292 23364 19296 23420
rect 19232 23360 19296 23364
rect 26912 23420 26976 23424
rect 26912 23364 26916 23420
rect 26916 23364 26972 23420
rect 26972 23364 26976 23420
rect 26912 23360 26976 23364
rect 26992 23420 27056 23424
rect 26992 23364 26996 23420
rect 26996 23364 27052 23420
rect 27052 23364 27056 23420
rect 26992 23360 27056 23364
rect 27072 23420 27136 23424
rect 27072 23364 27076 23420
rect 27076 23364 27132 23420
rect 27132 23364 27136 23420
rect 27072 23360 27136 23364
rect 27152 23420 27216 23424
rect 27152 23364 27156 23420
rect 27156 23364 27212 23420
rect 27212 23364 27216 23420
rect 27152 23360 27216 23364
rect 27232 23420 27296 23424
rect 27232 23364 27236 23420
rect 27236 23364 27292 23420
rect 27292 23364 27296 23420
rect 27232 23360 27296 23364
rect 3652 22876 3716 22880
rect 3652 22820 3656 22876
rect 3656 22820 3712 22876
rect 3712 22820 3716 22876
rect 3652 22816 3716 22820
rect 3732 22876 3796 22880
rect 3732 22820 3736 22876
rect 3736 22820 3792 22876
rect 3792 22820 3796 22876
rect 3732 22816 3796 22820
rect 3812 22876 3876 22880
rect 3812 22820 3816 22876
rect 3816 22820 3872 22876
rect 3872 22820 3876 22876
rect 3812 22816 3876 22820
rect 3892 22876 3956 22880
rect 3892 22820 3896 22876
rect 3896 22820 3952 22876
rect 3952 22820 3956 22876
rect 3892 22816 3956 22820
rect 3972 22876 4036 22880
rect 3972 22820 3976 22876
rect 3976 22820 4032 22876
rect 4032 22820 4036 22876
rect 3972 22816 4036 22820
rect 11652 22876 11716 22880
rect 11652 22820 11656 22876
rect 11656 22820 11712 22876
rect 11712 22820 11716 22876
rect 11652 22816 11716 22820
rect 11732 22876 11796 22880
rect 11732 22820 11736 22876
rect 11736 22820 11792 22876
rect 11792 22820 11796 22876
rect 11732 22816 11796 22820
rect 11812 22876 11876 22880
rect 11812 22820 11816 22876
rect 11816 22820 11872 22876
rect 11872 22820 11876 22876
rect 11812 22816 11876 22820
rect 11892 22876 11956 22880
rect 11892 22820 11896 22876
rect 11896 22820 11952 22876
rect 11952 22820 11956 22876
rect 11892 22816 11956 22820
rect 11972 22876 12036 22880
rect 11972 22820 11976 22876
rect 11976 22820 12032 22876
rect 12032 22820 12036 22876
rect 11972 22816 12036 22820
rect 19652 22876 19716 22880
rect 19652 22820 19656 22876
rect 19656 22820 19712 22876
rect 19712 22820 19716 22876
rect 19652 22816 19716 22820
rect 19732 22876 19796 22880
rect 19732 22820 19736 22876
rect 19736 22820 19792 22876
rect 19792 22820 19796 22876
rect 19732 22816 19796 22820
rect 19812 22876 19876 22880
rect 19812 22820 19816 22876
rect 19816 22820 19872 22876
rect 19872 22820 19876 22876
rect 19812 22816 19876 22820
rect 19892 22876 19956 22880
rect 19892 22820 19896 22876
rect 19896 22820 19952 22876
rect 19952 22820 19956 22876
rect 19892 22816 19956 22820
rect 19972 22876 20036 22880
rect 19972 22820 19976 22876
rect 19976 22820 20032 22876
rect 20032 22820 20036 22876
rect 19972 22816 20036 22820
rect 27652 22876 27716 22880
rect 27652 22820 27656 22876
rect 27656 22820 27712 22876
rect 27712 22820 27716 22876
rect 27652 22816 27716 22820
rect 27732 22876 27796 22880
rect 27732 22820 27736 22876
rect 27736 22820 27792 22876
rect 27792 22820 27796 22876
rect 27732 22816 27796 22820
rect 27812 22876 27876 22880
rect 27812 22820 27816 22876
rect 27816 22820 27872 22876
rect 27872 22820 27876 22876
rect 27812 22816 27876 22820
rect 27892 22876 27956 22880
rect 27892 22820 27896 22876
rect 27896 22820 27952 22876
rect 27952 22820 27956 22876
rect 27892 22816 27956 22820
rect 27972 22876 28036 22880
rect 27972 22820 27976 22876
rect 27976 22820 28032 22876
rect 28032 22820 28036 22876
rect 27972 22816 28036 22820
rect 2912 22332 2976 22336
rect 2912 22276 2916 22332
rect 2916 22276 2972 22332
rect 2972 22276 2976 22332
rect 2912 22272 2976 22276
rect 2992 22332 3056 22336
rect 2992 22276 2996 22332
rect 2996 22276 3052 22332
rect 3052 22276 3056 22332
rect 2992 22272 3056 22276
rect 3072 22332 3136 22336
rect 3072 22276 3076 22332
rect 3076 22276 3132 22332
rect 3132 22276 3136 22332
rect 3072 22272 3136 22276
rect 3152 22332 3216 22336
rect 3152 22276 3156 22332
rect 3156 22276 3212 22332
rect 3212 22276 3216 22332
rect 3152 22272 3216 22276
rect 3232 22332 3296 22336
rect 3232 22276 3236 22332
rect 3236 22276 3292 22332
rect 3292 22276 3296 22332
rect 3232 22272 3296 22276
rect 10912 22332 10976 22336
rect 10912 22276 10916 22332
rect 10916 22276 10972 22332
rect 10972 22276 10976 22332
rect 10912 22272 10976 22276
rect 10992 22332 11056 22336
rect 10992 22276 10996 22332
rect 10996 22276 11052 22332
rect 11052 22276 11056 22332
rect 10992 22272 11056 22276
rect 11072 22332 11136 22336
rect 11072 22276 11076 22332
rect 11076 22276 11132 22332
rect 11132 22276 11136 22332
rect 11072 22272 11136 22276
rect 11152 22332 11216 22336
rect 11152 22276 11156 22332
rect 11156 22276 11212 22332
rect 11212 22276 11216 22332
rect 11152 22272 11216 22276
rect 11232 22332 11296 22336
rect 11232 22276 11236 22332
rect 11236 22276 11292 22332
rect 11292 22276 11296 22332
rect 11232 22272 11296 22276
rect 18912 22332 18976 22336
rect 18912 22276 18916 22332
rect 18916 22276 18972 22332
rect 18972 22276 18976 22332
rect 18912 22272 18976 22276
rect 18992 22332 19056 22336
rect 18992 22276 18996 22332
rect 18996 22276 19052 22332
rect 19052 22276 19056 22332
rect 18992 22272 19056 22276
rect 19072 22332 19136 22336
rect 19072 22276 19076 22332
rect 19076 22276 19132 22332
rect 19132 22276 19136 22332
rect 19072 22272 19136 22276
rect 19152 22332 19216 22336
rect 19152 22276 19156 22332
rect 19156 22276 19212 22332
rect 19212 22276 19216 22332
rect 19152 22272 19216 22276
rect 19232 22332 19296 22336
rect 19232 22276 19236 22332
rect 19236 22276 19292 22332
rect 19292 22276 19296 22332
rect 19232 22272 19296 22276
rect 26912 22332 26976 22336
rect 26912 22276 26916 22332
rect 26916 22276 26972 22332
rect 26972 22276 26976 22332
rect 26912 22272 26976 22276
rect 26992 22332 27056 22336
rect 26992 22276 26996 22332
rect 26996 22276 27052 22332
rect 27052 22276 27056 22332
rect 26992 22272 27056 22276
rect 27072 22332 27136 22336
rect 27072 22276 27076 22332
rect 27076 22276 27132 22332
rect 27132 22276 27136 22332
rect 27072 22272 27136 22276
rect 27152 22332 27216 22336
rect 27152 22276 27156 22332
rect 27156 22276 27212 22332
rect 27212 22276 27216 22332
rect 27152 22272 27216 22276
rect 27232 22332 27296 22336
rect 27232 22276 27236 22332
rect 27236 22276 27292 22332
rect 27292 22276 27296 22332
rect 27232 22272 27296 22276
rect 3652 21788 3716 21792
rect 3652 21732 3656 21788
rect 3656 21732 3712 21788
rect 3712 21732 3716 21788
rect 3652 21728 3716 21732
rect 3732 21788 3796 21792
rect 3732 21732 3736 21788
rect 3736 21732 3792 21788
rect 3792 21732 3796 21788
rect 3732 21728 3796 21732
rect 3812 21788 3876 21792
rect 3812 21732 3816 21788
rect 3816 21732 3872 21788
rect 3872 21732 3876 21788
rect 3812 21728 3876 21732
rect 3892 21788 3956 21792
rect 3892 21732 3896 21788
rect 3896 21732 3952 21788
rect 3952 21732 3956 21788
rect 3892 21728 3956 21732
rect 3972 21788 4036 21792
rect 3972 21732 3976 21788
rect 3976 21732 4032 21788
rect 4032 21732 4036 21788
rect 3972 21728 4036 21732
rect 11652 21788 11716 21792
rect 11652 21732 11656 21788
rect 11656 21732 11712 21788
rect 11712 21732 11716 21788
rect 11652 21728 11716 21732
rect 11732 21788 11796 21792
rect 11732 21732 11736 21788
rect 11736 21732 11792 21788
rect 11792 21732 11796 21788
rect 11732 21728 11796 21732
rect 11812 21788 11876 21792
rect 11812 21732 11816 21788
rect 11816 21732 11872 21788
rect 11872 21732 11876 21788
rect 11812 21728 11876 21732
rect 11892 21788 11956 21792
rect 11892 21732 11896 21788
rect 11896 21732 11952 21788
rect 11952 21732 11956 21788
rect 11892 21728 11956 21732
rect 11972 21788 12036 21792
rect 11972 21732 11976 21788
rect 11976 21732 12032 21788
rect 12032 21732 12036 21788
rect 11972 21728 12036 21732
rect 19652 21788 19716 21792
rect 19652 21732 19656 21788
rect 19656 21732 19712 21788
rect 19712 21732 19716 21788
rect 19652 21728 19716 21732
rect 19732 21788 19796 21792
rect 19732 21732 19736 21788
rect 19736 21732 19792 21788
rect 19792 21732 19796 21788
rect 19732 21728 19796 21732
rect 19812 21788 19876 21792
rect 19812 21732 19816 21788
rect 19816 21732 19872 21788
rect 19872 21732 19876 21788
rect 19812 21728 19876 21732
rect 19892 21788 19956 21792
rect 19892 21732 19896 21788
rect 19896 21732 19952 21788
rect 19952 21732 19956 21788
rect 19892 21728 19956 21732
rect 19972 21788 20036 21792
rect 19972 21732 19976 21788
rect 19976 21732 20032 21788
rect 20032 21732 20036 21788
rect 19972 21728 20036 21732
rect 27652 21788 27716 21792
rect 27652 21732 27656 21788
rect 27656 21732 27712 21788
rect 27712 21732 27716 21788
rect 27652 21728 27716 21732
rect 27732 21788 27796 21792
rect 27732 21732 27736 21788
rect 27736 21732 27792 21788
rect 27792 21732 27796 21788
rect 27732 21728 27796 21732
rect 27812 21788 27876 21792
rect 27812 21732 27816 21788
rect 27816 21732 27872 21788
rect 27872 21732 27876 21788
rect 27812 21728 27876 21732
rect 27892 21788 27956 21792
rect 27892 21732 27896 21788
rect 27896 21732 27952 21788
rect 27952 21732 27956 21788
rect 27892 21728 27956 21732
rect 27972 21788 28036 21792
rect 27972 21732 27976 21788
rect 27976 21732 28032 21788
rect 28032 21732 28036 21788
rect 27972 21728 28036 21732
rect 2912 21244 2976 21248
rect 2912 21188 2916 21244
rect 2916 21188 2972 21244
rect 2972 21188 2976 21244
rect 2912 21184 2976 21188
rect 2992 21244 3056 21248
rect 2992 21188 2996 21244
rect 2996 21188 3052 21244
rect 3052 21188 3056 21244
rect 2992 21184 3056 21188
rect 3072 21244 3136 21248
rect 3072 21188 3076 21244
rect 3076 21188 3132 21244
rect 3132 21188 3136 21244
rect 3072 21184 3136 21188
rect 3152 21244 3216 21248
rect 3152 21188 3156 21244
rect 3156 21188 3212 21244
rect 3212 21188 3216 21244
rect 3152 21184 3216 21188
rect 3232 21244 3296 21248
rect 3232 21188 3236 21244
rect 3236 21188 3292 21244
rect 3292 21188 3296 21244
rect 3232 21184 3296 21188
rect 10912 21244 10976 21248
rect 10912 21188 10916 21244
rect 10916 21188 10972 21244
rect 10972 21188 10976 21244
rect 10912 21184 10976 21188
rect 10992 21244 11056 21248
rect 10992 21188 10996 21244
rect 10996 21188 11052 21244
rect 11052 21188 11056 21244
rect 10992 21184 11056 21188
rect 11072 21244 11136 21248
rect 11072 21188 11076 21244
rect 11076 21188 11132 21244
rect 11132 21188 11136 21244
rect 11072 21184 11136 21188
rect 11152 21244 11216 21248
rect 11152 21188 11156 21244
rect 11156 21188 11212 21244
rect 11212 21188 11216 21244
rect 11152 21184 11216 21188
rect 11232 21244 11296 21248
rect 11232 21188 11236 21244
rect 11236 21188 11292 21244
rect 11292 21188 11296 21244
rect 11232 21184 11296 21188
rect 18912 21244 18976 21248
rect 18912 21188 18916 21244
rect 18916 21188 18972 21244
rect 18972 21188 18976 21244
rect 18912 21184 18976 21188
rect 18992 21244 19056 21248
rect 18992 21188 18996 21244
rect 18996 21188 19052 21244
rect 19052 21188 19056 21244
rect 18992 21184 19056 21188
rect 19072 21244 19136 21248
rect 19072 21188 19076 21244
rect 19076 21188 19132 21244
rect 19132 21188 19136 21244
rect 19072 21184 19136 21188
rect 19152 21244 19216 21248
rect 19152 21188 19156 21244
rect 19156 21188 19212 21244
rect 19212 21188 19216 21244
rect 19152 21184 19216 21188
rect 19232 21244 19296 21248
rect 19232 21188 19236 21244
rect 19236 21188 19292 21244
rect 19292 21188 19296 21244
rect 19232 21184 19296 21188
rect 26912 21244 26976 21248
rect 26912 21188 26916 21244
rect 26916 21188 26972 21244
rect 26972 21188 26976 21244
rect 26912 21184 26976 21188
rect 26992 21244 27056 21248
rect 26992 21188 26996 21244
rect 26996 21188 27052 21244
rect 27052 21188 27056 21244
rect 26992 21184 27056 21188
rect 27072 21244 27136 21248
rect 27072 21188 27076 21244
rect 27076 21188 27132 21244
rect 27132 21188 27136 21244
rect 27072 21184 27136 21188
rect 27152 21244 27216 21248
rect 27152 21188 27156 21244
rect 27156 21188 27212 21244
rect 27212 21188 27216 21244
rect 27152 21184 27216 21188
rect 27232 21244 27296 21248
rect 27232 21188 27236 21244
rect 27236 21188 27292 21244
rect 27292 21188 27296 21244
rect 27232 21184 27296 21188
rect 3652 20700 3716 20704
rect 3652 20644 3656 20700
rect 3656 20644 3712 20700
rect 3712 20644 3716 20700
rect 3652 20640 3716 20644
rect 3732 20700 3796 20704
rect 3732 20644 3736 20700
rect 3736 20644 3792 20700
rect 3792 20644 3796 20700
rect 3732 20640 3796 20644
rect 3812 20700 3876 20704
rect 3812 20644 3816 20700
rect 3816 20644 3872 20700
rect 3872 20644 3876 20700
rect 3812 20640 3876 20644
rect 3892 20700 3956 20704
rect 3892 20644 3896 20700
rect 3896 20644 3952 20700
rect 3952 20644 3956 20700
rect 3892 20640 3956 20644
rect 3972 20700 4036 20704
rect 3972 20644 3976 20700
rect 3976 20644 4032 20700
rect 4032 20644 4036 20700
rect 3972 20640 4036 20644
rect 11652 20700 11716 20704
rect 11652 20644 11656 20700
rect 11656 20644 11712 20700
rect 11712 20644 11716 20700
rect 11652 20640 11716 20644
rect 11732 20700 11796 20704
rect 11732 20644 11736 20700
rect 11736 20644 11792 20700
rect 11792 20644 11796 20700
rect 11732 20640 11796 20644
rect 11812 20700 11876 20704
rect 11812 20644 11816 20700
rect 11816 20644 11872 20700
rect 11872 20644 11876 20700
rect 11812 20640 11876 20644
rect 11892 20700 11956 20704
rect 11892 20644 11896 20700
rect 11896 20644 11952 20700
rect 11952 20644 11956 20700
rect 11892 20640 11956 20644
rect 11972 20700 12036 20704
rect 11972 20644 11976 20700
rect 11976 20644 12032 20700
rect 12032 20644 12036 20700
rect 11972 20640 12036 20644
rect 19652 20700 19716 20704
rect 19652 20644 19656 20700
rect 19656 20644 19712 20700
rect 19712 20644 19716 20700
rect 19652 20640 19716 20644
rect 19732 20700 19796 20704
rect 19732 20644 19736 20700
rect 19736 20644 19792 20700
rect 19792 20644 19796 20700
rect 19732 20640 19796 20644
rect 19812 20700 19876 20704
rect 19812 20644 19816 20700
rect 19816 20644 19872 20700
rect 19872 20644 19876 20700
rect 19812 20640 19876 20644
rect 19892 20700 19956 20704
rect 19892 20644 19896 20700
rect 19896 20644 19952 20700
rect 19952 20644 19956 20700
rect 19892 20640 19956 20644
rect 19972 20700 20036 20704
rect 19972 20644 19976 20700
rect 19976 20644 20032 20700
rect 20032 20644 20036 20700
rect 19972 20640 20036 20644
rect 27652 20700 27716 20704
rect 27652 20644 27656 20700
rect 27656 20644 27712 20700
rect 27712 20644 27716 20700
rect 27652 20640 27716 20644
rect 27732 20700 27796 20704
rect 27732 20644 27736 20700
rect 27736 20644 27792 20700
rect 27792 20644 27796 20700
rect 27732 20640 27796 20644
rect 27812 20700 27876 20704
rect 27812 20644 27816 20700
rect 27816 20644 27872 20700
rect 27872 20644 27876 20700
rect 27812 20640 27876 20644
rect 27892 20700 27956 20704
rect 27892 20644 27896 20700
rect 27896 20644 27952 20700
rect 27952 20644 27956 20700
rect 27892 20640 27956 20644
rect 27972 20700 28036 20704
rect 27972 20644 27976 20700
rect 27976 20644 28032 20700
rect 28032 20644 28036 20700
rect 27972 20640 28036 20644
rect 2912 20156 2976 20160
rect 2912 20100 2916 20156
rect 2916 20100 2972 20156
rect 2972 20100 2976 20156
rect 2912 20096 2976 20100
rect 2992 20156 3056 20160
rect 2992 20100 2996 20156
rect 2996 20100 3052 20156
rect 3052 20100 3056 20156
rect 2992 20096 3056 20100
rect 3072 20156 3136 20160
rect 3072 20100 3076 20156
rect 3076 20100 3132 20156
rect 3132 20100 3136 20156
rect 3072 20096 3136 20100
rect 3152 20156 3216 20160
rect 3152 20100 3156 20156
rect 3156 20100 3212 20156
rect 3212 20100 3216 20156
rect 3152 20096 3216 20100
rect 3232 20156 3296 20160
rect 3232 20100 3236 20156
rect 3236 20100 3292 20156
rect 3292 20100 3296 20156
rect 3232 20096 3296 20100
rect 10912 20156 10976 20160
rect 10912 20100 10916 20156
rect 10916 20100 10972 20156
rect 10972 20100 10976 20156
rect 10912 20096 10976 20100
rect 10992 20156 11056 20160
rect 10992 20100 10996 20156
rect 10996 20100 11052 20156
rect 11052 20100 11056 20156
rect 10992 20096 11056 20100
rect 11072 20156 11136 20160
rect 11072 20100 11076 20156
rect 11076 20100 11132 20156
rect 11132 20100 11136 20156
rect 11072 20096 11136 20100
rect 11152 20156 11216 20160
rect 11152 20100 11156 20156
rect 11156 20100 11212 20156
rect 11212 20100 11216 20156
rect 11152 20096 11216 20100
rect 11232 20156 11296 20160
rect 11232 20100 11236 20156
rect 11236 20100 11292 20156
rect 11292 20100 11296 20156
rect 11232 20096 11296 20100
rect 18912 20156 18976 20160
rect 18912 20100 18916 20156
rect 18916 20100 18972 20156
rect 18972 20100 18976 20156
rect 18912 20096 18976 20100
rect 18992 20156 19056 20160
rect 18992 20100 18996 20156
rect 18996 20100 19052 20156
rect 19052 20100 19056 20156
rect 18992 20096 19056 20100
rect 19072 20156 19136 20160
rect 19072 20100 19076 20156
rect 19076 20100 19132 20156
rect 19132 20100 19136 20156
rect 19072 20096 19136 20100
rect 19152 20156 19216 20160
rect 19152 20100 19156 20156
rect 19156 20100 19212 20156
rect 19212 20100 19216 20156
rect 19152 20096 19216 20100
rect 19232 20156 19296 20160
rect 19232 20100 19236 20156
rect 19236 20100 19292 20156
rect 19292 20100 19296 20156
rect 19232 20096 19296 20100
rect 26912 20156 26976 20160
rect 26912 20100 26916 20156
rect 26916 20100 26972 20156
rect 26972 20100 26976 20156
rect 26912 20096 26976 20100
rect 26992 20156 27056 20160
rect 26992 20100 26996 20156
rect 26996 20100 27052 20156
rect 27052 20100 27056 20156
rect 26992 20096 27056 20100
rect 27072 20156 27136 20160
rect 27072 20100 27076 20156
rect 27076 20100 27132 20156
rect 27132 20100 27136 20156
rect 27072 20096 27136 20100
rect 27152 20156 27216 20160
rect 27152 20100 27156 20156
rect 27156 20100 27212 20156
rect 27212 20100 27216 20156
rect 27152 20096 27216 20100
rect 27232 20156 27296 20160
rect 27232 20100 27236 20156
rect 27236 20100 27292 20156
rect 27292 20100 27296 20156
rect 27232 20096 27296 20100
rect 3652 19612 3716 19616
rect 3652 19556 3656 19612
rect 3656 19556 3712 19612
rect 3712 19556 3716 19612
rect 3652 19552 3716 19556
rect 3732 19612 3796 19616
rect 3732 19556 3736 19612
rect 3736 19556 3792 19612
rect 3792 19556 3796 19612
rect 3732 19552 3796 19556
rect 3812 19612 3876 19616
rect 3812 19556 3816 19612
rect 3816 19556 3872 19612
rect 3872 19556 3876 19612
rect 3812 19552 3876 19556
rect 3892 19612 3956 19616
rect 3892 19556 3896 19612
rect 3896 19556 3952 19612
rect 3952 19556 3956 19612
rect 3892 19552 3956 19556
rect 3972 19612 4036 19616
rect 3972 19556 3976 19612
rect 3976 19556 4032 19612
rect 4032 19556 4036 19612
rect 3972 19552 4036 19556
rect 11652 19612 11716 19616
rect 11652 19556 11656 19612
rect 11656 19556 11712 19612
rect 11712 19556 11716 19612
rect 11652 19552 11716 19556
rect 11732 19612 11796 19616
rect 11732 19556 11736 19612
rect 11736 19556 11792 19612
rect 11792 19556 11796 19612
rect 11732 19552 11796 19556
rect 11812 19612 11876 19616
rect 11812 19556 11816 19612
rect 11816 19556 11872 19612
rect 11872 19556 11876 19612
rect 11812 19552 11876 19556
rect 11892 19612 11956 19616
rect 11892 19556 11896 19612
rect 11896 19556 11952 19612
rect 11952 19556 11956 19612
rect 11892 19552 11956 19556
rect 11972 19612 12036 19616
rect 11972 19556 11976 19612
rect 11976 19556 12032 19612
rect 12032 19556 12036 19612
rect 11972 19552 12036 19556
rect 19652 19612 19716 19616
rect 19652 19556 19656 19612
rect 19656 19556 19712 19612
rect 19712 19556 19716 19612
rect 19652 19552 19716 19556
rect 19732 19612 19796 19616
rect 19732 19556 19736 19612
rect 19736 19556 19792 19612
rect 19792 19556 19796 19612
rect 19732 19552 19796 19556
rect 19812 19612 19876 19616
rect 19812 19556 19816 19612
rect 19816 19556 19872 19612
rect 19872 19556 19876 19612
rect 19812 19552 19876 19556
rect 19892 19612 19956 19616
rect 19892 19556 19896 19612
rect 19896 19556 19952 19612
rect 19952 19556 19956 19612
rect 19892 19552 19956 19556
rect 19972 19612 20036 19616
rect 19972 19556 19976 19612
rect 19976 19556 20032 19612
rect 20032 19556 20036 19612
rect 19972 19552 20036 19556
rect 27652 19612 27716 19616
rect 27652 19556 27656 19612
rect 27656 19556 27712 19612
rect 27712 19556 27716 19612
rect 27652 19552 27716 19556
rect 27732 19612 27796 19616
rect 27732 19556 27736 19612
rect 27736 19556 27792 19612
rect 27792 19556 27796 19612
rect 27732 19552 27796 19556
rect 27812 19612 27876 19616
rect 27812 19556 27816 19612
rect 27816 19556 27872 19612
rect 27872 19556 27876 19612
rect 27812 19552 27876 19556
rect 27892 19612 27956 19616
rect 27892 19556 27896 19612
rect 27896 19556 27952 19612
rect 27952 19556 27956 19612
rect 27892 19552 27956 19556
rect 27972 19612 28036 19616
rect 27972 19556 27976 19612
rect 27976 19556 28032 19612
rect 28032 19556 28036 19612
rect 27972 19552 28036 19556
rect 2912 19068 2976 19072
rect 2912 19012 2916 19068
rect 2916 19012 2972 19068
rect 2972 19012 2976 19068
rect 2912 19008 2976 19012
rect 2992 19068 3056 19072
rect 2992 19012 2996 19068
rect 2996 19012 3052 19068
rect 3052 19012 3056 19068
rect 2992 19008 3056 19012
rect 3072 19068 3136 19072
rect 3072 19012 3076 19068
rect 3076 19012 3132 19068
rect 3132 19012 3136 19068
rect 3072 19008 3136 19012
rect 3152 19068 3216 19072
rect 3152 19012 3156 19068
rect 3156 19012 3212 19068
rect 3212 19012 3216 19068
rect 3152 19008 3216 19012
rect 3232 19068 3296 19072
rect 3232 19012 3236 19068
rect 3236 19012 3292 19068
rect 3292 19012 3296 19068
rect 3232 19008 3296 19012
rect 10912 19068 10976 19072
rect 10912 19012 10916 19068
rect 10916 19012 10972 19068
rect 10972 19012 10976 19068
rect 10912 19008 10976 19012
rect 10992 19068 11056 19072
rect 10992 19012 10996 19068
rect 10996 19012 11052 19068
rect 11052 19012 11056 19068
rect 10992 19008 11056 19012
rect 11072 19068 11136 19072
rect 11072 19012 11076 19068
rect 11076 19012 11132 19068
rect 11132 19012 11136 19068
rect 11072 19008 11136 19012
rect 11152 19068 11216 19072
rect 11152 19012 11156 19068
rect 11156 19012 11212 19068
rect 11212 19012 11216 19068
rect 11152 19008 11216 19012
rect 11232 19068 11296 19072
rect 11232 19012 11236 19068
rect 11236 19012 11292 19068
rect 11292 19012 11296 19068
rect 11232 19008 11296 19012
rect 18912 19068 18976 19072
rect 18912 19012 18916 19068
rect 18916 19012 18972 19068
rect 18972 19012 18976 19068
rect 18912 19008 18976 19012
rect 18992 19068 19056 19072
rect 18992 19012 18996 19068
rect 18996 19012 19052 19068
rect 19052 19012 19056 19068
rect 18992 19008 19056 19012
rect 19072 19068 19136 19072
rect 19072 19012 19076 19068
rect 19076 19012 19132 19068
rect 19132 19012 19136 19068
rect 19072 19008 19136 19012
rect 19152 19068 19216 19072
rect 19152 19012 19156 19068
rect 19156 19012 19212 19068
rect 19212 19012 19216 19068
rect 19152 19008 19216 19012
rect 19232 19068 19296 19072
rect 19232 19012 19236 19068
rect 19236 19012 19292 19068
rect 19292 19012 19296 19068
rect 19232 19008 19296 19012
rect 26912 19068 26976 19072
rect 26912 19012 26916 19068
rect 26916 19012 26972 19068
rect 26972 19012 26976 19068
rect 26912 19008 26976 19012
rect 26992 19068 27056 19072
rect 26992 19012 26996 19068
rect 26996 19012 27052 19068
rect 27052 19012 27056 19068
rect 26992 19008 27056 19012
rect 27072 19068 27136 19072
rect 27072 19012 27076 19068
rect 27076 19012 27132 19068
rect 27132 19012 27136 19068
rect 27072 19008 27136 19012
rect 27152 19068 27216 19072
rect 27152 19012 27156 19068
rect 27156 19012 27212 19068
rect 27212 19012 27216 19068
rect 27152 19008 27216 19012
rect 27232 19068 27296 19072
rect 27232 19012 27236 19068
rect 27236 19012 27292 19068
rect 27292 19012 27296 19068
rect 27232 19008 27296 19012
rect 3652 18524 3716 18528
rect 3652 18468 3656 18524
rect 3656 18468 3712 18524
rect 3712 18468 3716 18524
rect 3652 18464 3716 18468
rect 3732 18524 3796 18528
rect 3732 18468 3736 18524
rect 3736 18468 3792 18524
rect 3792 18468 3796 18524
rect 3732 18464 3796 18468
rect 3812 18524 3876 18528
rect 3812 18468 3816 18524
rect 3816 18468 3872 18524
rect 3872 18468 3876 18524
rect 3812 18464 3876 18468
rect 3892 18524 3956 18528
rect 3892 18468 3896 18524
rect 3896 18468 3952 18524
rect 3952 18468 3956 18524
rect 3892 18464 3956 18468
rect 3972 18524 4036 18528
rect 3972 18468 3976 18524
rect 3976 18468 4032 18524
rect 4032 18468 4036 18524
rect 3972 18464 4036 18468
rect 11652 18524 11716 18528
rect 11652 18468 11656 18524
rect 11656 18468 11712 18524
rect 11712 18468 11716 18524
rect 11652 18464 11716 18468
rect 11732 18524 11796 18528
rect 11732 18468 11736 18524
rect 11736 18468 11792 18524
rect 11792 18468 11796 18524
rect 11732 18464 11796 18468
rect 11812 18524 11876 18528
rect 11812 18468 11816 18524
rect 11816 18468 11872 18524
rect 11872 18468 11876 18524
rect 11812 18464 11876 18468
rect 11892 18524 11956 18528
rect 11892 18468 11896 18524
rect 11896 18468 11952 18524
rect 11952 18468 11956 18524
rect 11892 18464 11956 18468
rect 11972 18524 12036 18528
rect 11972 18468 11976 18524
rect 11976 18468 12032 18524
rect 12032 18468 12036 18524
rect 11972 18464 12036 18468
rect 19652 18524 19716 18528
rect 19652 18468 19656 18524
rect 19656 18468 19712 18524
rect 19712 18468 19716 18524
rect 19652 18464 19716 18468
rect 19732 18524 19796 18528
rect 19732 18468 19736 18524
rect 19736 18468 19792 18524
rect 19792 18468 19796 18524
rect 19732 18464 19796 18468
rect 19812 18524 19876 18528
rect 19812 18468 19816 18524
rect 19816 18468 19872 18524
rect 19872 18468 19876 18524
rect 19812 18464 19876 18468
rect 19892 18524 19956 18528
rect 19892 18468 19896 18524
rect 19896 18468 19952 18524
rect 19952 18468 19956 18524
rect 19892 18464 19956 18468
rect 19972 18524 20036 18528
rect 19972 18468 19976 18524
rect 19976 18468 20032 18524
rect 20032 18468 20036 18524
rect 19972 18464 20036 18468
rect 27652 18524 27716 18528
rect 27652 18468 27656 18524
rect 27656 18468 27712 18524
rect 27712 18468 27716 18524
rect 27652 18464 27716 18468
rect 27732 18524 27796 18528
rect 27732 18468 27736 18524
rect 27736 18468 27792 18524
rect 27792 18468 27796 18524
rect 27732 18464 27796 18468
rect 27812 18524 27876 18528
rect 27812 18468 27816 18524
rect 27816 18468 27872 18524
rect 27872 18468 27876 18524
rect 27812 18464 27876 18468
rect 27892 18524 27956 18528
rect 27892 18468 27896 18524
rect 27896 18468 27952 18524
rect 27952 18468 27956 18524
rect 27892 18464 27956 18468
rect 27972 18524 28036 18528
rect 27972 18468 27976 18524
rect 27976 18468 28032 18524
rect 28032 18468 28036 18524
rect 27972 18464 28036 18468
rect 2912 17980 2976 17984
rect 2912 17924 2916 17980
rect 2916 17924 2972 17980
rect 2972 17924 2976 17980
rect 2912 17920 2976 17924
rect 2992 17980 3056 17984
rect 2992 17924 2996 17980
rect 2996 17924 3052 17980
rect 3052 17924 3056 17980
rect 2992 17920 3056 17924
rect 3072 17980 3136 17984
rect 3072 17924 3076 17980
rect 3076 17924 3132 17980
rect 3132 17924 3136 17980
rect 3072 17920 3136 17924
rect 3152 17980 3216 17984
rect 3152 17924 3156 17980
rect 3156 17924 3212 17980
rect 3212 17924 3216 17980
rect 3152 17920 3216 17924
rect 3232 17980 3296 17984
rect 3232 17924 3236 17980
rect 3236 17924 3292 17980
rect 3292 17924 3296 17980
rect 3232 17920 3296 17924
rect 10912 17980 10976 17984
rect 10912 17924 10916 17980
rect 10916 17924 10972 17980
rect 10972 17924 10976 17980
rect 10912 17920 10976 17924
rect 10992 17980 11056 17984
rect 10992 17924 10996 17980
rect 10996 17924 11052 17980
rect 11052 17924 11056 17980
rect 10992 17920 11056 17924
rect 11072 17980 11136 17984
rect 11072 17924 11076 17980
rect 11076 17924 11132 17980
rect 11132 17924 11136 17980
rect 11072 17920 11136 17924
rect 11152 17980 11216 17984
rect 11152 17924 11156 17980
rect 11156 17924 11212 17980
rect 11212 17924 11216 17980
rect 11152 17920 11216 17924
rect 11232 17980 11296 17984
rect 11232 17924 11236 17980
rect 11236 17924 11292 17980
rect 11292 17924 11296 17980
rect 11232 17920 11296 17924
rect 18912 17980 18976 17984
rect 18912 17924 18916 17980
rect 18916 17924 18972 17980
rect 18972 17924 18976 17980
rect 18912 17920 18976 17924
rect 18992 17980 19056 17984
rect 18992 17924 18996 17980
rect 18996 17924 19052 17980
rect 19052 17924 19056 17980
rect 18992 17920 19056 17924
rect 19072 17980 19136 17984
rect 19072 17924 19076 17980
rect 19076 17924 19132 17980
rect 19132 17924 19136 17980
rect 19072 17920 19136 17924
rect 19152 17980 19216 17984
rect 19152 17924 19156 17980
rect 19156 17924 19212 17980
rect 19212 17924 19216 17980
rect 19152 17920 19216 17924
rect 19232 17980 19296 17984
rect 19232 17924 19236 17980
rect 19236 17924 19292 17980
rect 19292 17924 19296 17980
rect 19232 17920 19296 17924
rect 26912 17980 26976 17984
rect 26912 17924 26916 17980
rect 26916 17924 26972 17980
rect 26972 17924 26976 17980
rect 26912 17920 26976 17924
rect 26992 17980 27056 17984
rect 26992 17924 26996 17980
rect 26996 17924 27052 17980
rect 27052 17924 27056 17980
rect 26992 17920 27056 17924
rect 27072 17980 27136 17984
rect 27072 17924 27076 17980
rect 27076 17924 27132 17980
rect 27132 17924 27136 17980
rect 27072 17920 27136 17924
rect 27152 17980 27216 17984
rect 27152 17924 27156 17980
rect 27156 17924 27212 17980
rect 27212 17924 27216 17980
rect 27152 17920 27216 17924
rect 27232 17980 27296 17984
rect 27232 17924 27236 17980
rect 27236 17924 27292 17980
rect 27292 17924 27296 17980
rect 27232 17920 27296 17924
rect 3652 17436 3716 17440
rect 3652 17380 3656 17436
rect 3656 17380 3712 17436
rect 3712 17380 3716 17436
rect 3652 17376 3716 17380
rect 3732 17436 3796 17440
rect 3732 17380 3736 17436
rect 3736 17380 3792 17436
rect 3792 17380 3796 17436
rect 3732 17376 3796 17380
rect 3812 17436 3876 17440
rect 3812 17380 3816 17436
rect 3816 17380 3872 17436
rect 3872 17380 3876 17436
rect 3812 17376 3876 17380
rect 3892 17436 3956 17440
rect 3892 17380 3896 17436
rect 3896 17380 3952 17436
rect 3952 17380 3956 17436
rect 3892 17376 3956 17380
rect 3972 17436 4036 17440
rect 3972 17380 3976 17436
rect 3976 17380 4032 17436
rect 4032 17380 4036 17436
rect 3972 17376 4036 17380
rect 11652 17436 11716 17440
rect 11652 17380 11656 17436
rect 11656 17380 11712 17436
rect 11712 17380 11716 17436
rect 11652 17376 11716 17380
rect 11732 17436 11796 17440
rect 11732 17380 11736 17436
rect 11736 17380 11792 17436
rect 11792 17380 11796 17436
rect 11732 17376 11796 17380
rect 11812 17436 11876 17440
rect 11812 17380 11816 17436
rect 11816 17380 11872 17436
rect 11872 17380 11876 17436
rect 11812 17376 11876 17380
rect 11892 17436 11956 17440
rect 11892 17380 11896 17436
rect 11896 17380 11952 17436
rect 11952 17380 11956 17436
rect 11892 17376 11956 17380
rect 11972 17436 12036 17440
rect 11972 17380 11976 17436
rect 11976 17380 12032 17436
rect 12032 17380 12036 17436
rect 11972 17376 12036 17380
rect 19652 17436 19716 17440
rect 19652 17380 19656 17436
rect 19656 17380 19712 17436
rect 19712 17380 19716 17436
rect 19652 17376 19716 17380
rect 19732 17436 19796 17440
rect 19732 17380 19736 17436
rect 19736 17380 19792 17436
rect 19792 17380 19796 17436
rect 19732 17376 19796 17380
rect 19812 17436 19876 17440
rect 19812 17380 19816 17436
rect 19816 17380 19872 17436
rect 19872 17380 19876 17436
rect 19812 17376 19876 17380
rect 19892 17436 19956 17440
rect 19892 17380 19896 17436
rect 19896 17380 19952 17436
rect 19952 17380 19956 17436
rect 19892 17376 19956 17380
rect 19972 17436 20036 17440
rect 19972 17380 19976 17436
rect 19976 17380 20032 17436
rect 20032 17380 20036 17436
rect 19972 17376 20036 17380
rect 27652 17436 27716 17440
rect 27652 17380 27656 17436
rect 27656 17380 27712 17436
rect 27712 17380 27716 17436
rect 27652 17376 27716 17380
rect 27732 17436 27796 17440
rect 27732 17380 27736 17436
rect 27736 17380 27792 17436
rect 27792 17380 27796 17436
rect 27732 17376 27796 17380
rect 27812 17436 27876 17440
rect 27812 17380 27816 17436
rect 27816 17380 27872 17436
rect 27872 17380 27876 17436
rect 27812 17376 27876 17380
rect 27892 17436 27956 17440
rect 27892 17380 27896 17436
rect 27896 17380 27952 17436
rect 27952 17380 27956 17436
rect 27892 17376 27956 17380
rect 27972 17436 28036 17440
rect 27972 17380 27976 17436
rect 27976 17380 28032 17436
rect 28032 17380 28036 17436
rect 27972 17376 28036 17380
rect 2912 16892 2976 16896
rect 2912 16836 2916 16892
rect 2916 16836 2972 16892
rect 2972 16836 2976 16892
rect 2912 16832 2976 16836
rect 2992 16892 3056 16896
rect 2992 16836 2996 16892
rect 2996 16836 3052 16892
rect 3052 16836 3056 16892
rect 2992 16832 3056 16836
rect 3072 16892 3136 16896
rect 3072 16836 3076 16892
rect 3076 16836 3132 16892
rect 3132 16836 3136 16892
rect 3072 16832 3136 16836
rect 3152 16892 3216 16896
rect 3152 16836 3156 16892
rect 3156 16836 3212 16892
rect 3212 16836 3216 16892
rect 3152 16832 3216 16836
rect 3232 16892 3296 16896
rect 3232 16836 3236 16892
rect 3236 16836 3292 16892
rect 3292 16836 3296 16892
rect 3232 16832 3296 16836
rect 10912 16892 10976 16896
rect 10912 16836 10916 16892
rect 10916 16836 10972 16892
rect 10972 16836 10976 16892
rect 10912 16832 10976 16836
rect 10992 16892 11056 16896
rect 10992 16836 10996 16892
rect 10996 16836 11052 16892
rect 11052 16836 11056 16892
rect 10992 16832 11056 16836
rect 11072 16892 11136 16896
rect 11072 16836 11076 16892
rect 11076 16836 11132 16892
rect 11132 16836 11136 16892
rect 11072 16832 11136 16836
rect 11152 16892 11216 16896
rect 11152 16836 11156 16892
rect 11156 16836 11212 16892
rect 11212 16836 11216 16892
rect 11152 16832 11216 16836
rect 11232 16892 11296 16896
rect 11232 16836 11236 16892
rect 11236 16836 11292 16892
rect 11292 16836 11296 16892
rect 11232 16832 11296 16836
rect 18912 16892 18976 16896
rect 18912 16836 18916 16892
rect 18916 16836 18972 16892
rect 18972 16836 18976 16892
rect 18912 16832 18976 16836
rect 18992 16892 19056 16896
rect 18992 16836 18996 16892
rect 18996 16836 19052 16892
rect 19052 16836 19056 16892
rect 18992 16832 19056 16836
rect 19072 16892 19136 16896
rect 19072 16836 19076 16892
rect 19076 16836 19132 16892
rect 19132 16836 19136 16892
rect 19072 16832 19136 16836
rect 19152 16892 19216 16896
rect 19152 16836 19156 16892
rect 19156 16836 19212 16892
rect 19212 16836 19216 16892
rect 19152 16832 19216 16836
rect 19232 16892 19296 16896
rect 19232 16836 19236 16892
rect 19236 16836 19292 16892
rect 19292 16836 19296 16892
rect 19232 16832 19296 16836
rect 26912 16892 26976 16896
rect 26912 16836 26916 16892
rect 26916 16836 26972 16892
rect 26972 16836 26976 16892
rect 26912 16832 26976 16836
rect 26992 16892 27056 16896
rect 26992 16836 26996 16892
rect 26996 16836 27052 16892
rect 27052 16836 27056 16892
rect 26992 16832 27056 16836
rect 27072 16892 27136 16896
rect 27072 16836 27076 16892
rect 27076 16836 27132 16892
rect 27132 16836 27136 16892
rect 27072 16832 27136 16836
rect 27152 16892 27216 16896
rect 27152 16836 27156 16892
rect 27156 16836 27212 16892
rect 27212 16836 27216 16892
rect 27152 16832 27216 16836
rect 27232 16892 27296 16896
rect 27232 16836 27236 16892
rect 27236 16836 27292 16892
rect 27292 16836 27296 16892
rect 27232 16832 27296 16836
rect 3652 16348 3716 16352
rect 3652 16292 3656 16348
rect 3656 16292 3712 16348
rect 3712 16292 3716 16348
rect 3652 16288 3716 16292
rect 3732 16348 3796 16352
rect 3732 16292 3736 16348
rect 3736 16292 3792 16348
rect 3792 16292 3796 16348
rect 3732 16288 3796 16292
rect 3812 16348 3876 16352
rect 3812 16292 3816 16348
rect 3816 16292 3872 16348
rect 3872 16292 3876 16348
rect 3812 16288 3876 16292
rect 3892 16348 3956 16352
rect 3892 16292 3896 16348
rect 3896 16292 3952 16348
rect 3952 16292 3956 16348
rect 3892 16288 3956 16292
rect 3972 16348 4036 16352
rect 3972 16292 3976 16348
rect 3976 16292 4032 16348
rect 4032 16292 4036 16348
rect 3972 16288 4036 16292
rect 11652 16348 11716 16352
rect 11652 16292 11656 16348
rect 11656 16292 11712 16348
rect 11712 16292 11716 16348
rect 11652 16288 11716 16292
rect 11732 16348 11796 16352
rect 11732 16292 11736 16348
rect 11736 16292 11792 16348
rect 11792 16292 11796 16348
rect 11732 16288 11796 16292
rect 11812 16348 11876 16352
rect 11812 16292 11816 16348
rect 11816 16292 11872 16348
rect 11872 16292 11876 16348
rect 11812 16288 11876 16292
rect 11892 16348 11956 16352
rect 11892 16292 11896 16348
rect 11896 16292 11952 16348
rect 11952 16292 11956 16348
rect 11892 16288 11956 16292
rect 11972 16348 12036 16352
rect 11972 16292 11976 16348
rect 11976 16292 12032 16348
rect 12032 16292 12036 16348
rect 11972 16288 12036 16292
rect 19652 16348 19716 16352
rect 19652 16292 19656 16348
rect 19656 16292 19712 16348
rect 19712 16292 19716 16348
rect 19652 16288 19716 16292
rect 19732 16348 19796 16352
rect 19732 16292 19736 16348
rect 19736 16292 19792 16348
rect 19792 16292 19796 16348
rect 19732 16288 19796 16292
rect 19812 16348 19876 16352
rect 19812 16292 19816 16348
rect 19816 16292 19872 16348
rect 19872 16292 19876 16348
rect 19812 16288 19876 16292
rect 19892 16348 19956 16352
rect 19892 16292 19896 16348
rect 19896 16292 19952 16348
rect 19952 16292 19956 16348
rect 19892 16288 19956 16292
rect 19972 16348 20036 16352
rect 19972 16292 19976 16348
rect 19976 16292 20032 16348
rect 20032 16292 20036 16348
rect 19972 16288 20036 16292
rect 27652 16348 27716 16352
rect 27652 16292 27656 16348
rect 27656 16292 27712 16348
rect 27712 16292 27716 16348
rect 27652 16288 27716 16292
rect 27732 16348 27796 16352
rect 27732 16292 27736 16348
rect 27736 16292 27792 16348
rect 27792 16292 27796 16348
rect 27732 16288 27796 16292
rect 27812 16348 27876 16352
rect 27812 16292 27816 16348
rect 27816 16292 27872 16348
rect 27872 16292 27876 16348
rect 27812 16288 27876 16292
rect 27892 16348 27956 16352
rect 27892 16292 27896 16348
rect 27896 16292 27952 16348
rect 27952 16292 27956 16348
rect 27892 16288 27956 16292
rect 27972 16348 28036 16352
rect 27972 16292 27976 16348
rect 27976 16292 28032 16348
rect 28032 16292 28036 16348
rect 27972 16288 28036 16292
rect 2912 15804 2976 15808
rect 2912 15748 2916 15804
rect 2916 15748 2972 15804
rect 2972 15748 2976 15804
rect 2912 15744 2976 15748
rect 2992 15804 3056 15808
rect 2992 15748 2996 15804
rect 2996 15748 3052 15804
rect 3052 15748 3056 15804
rect 2992 15744 3056 15748
rect 3072 15804 3136 15808
rect 3072 15748 3076 15804
rect 3076 15748 3132 15804
rect 3132 15748 3136 15804
rect 3072 15744 3136 15748
rect 3152 15804 3216 15808
rect 3152 15748 3156 15804
rect 3156 15748 3212 15804
rect 3212 15748 3216 15804
rect 3152 15744 3216 15748
rect 3232 15804 3296 15808
rect 3232 15748 3236 15804
rect 3236 15748 3292 15804
rect 3292 15748 3296 15804
rect 3232 15744 3296 15748
rect 10912 15804 10976 15808
rect 10912 15748 10916 15804
rect 10916 15748 10972 15804
rect 10972 15748 10976 15804
rect 10912 15744 10976 15748
rect 10992 15804 11056 15808
rect 10992 15748 10996 15804
rect 10996 15748 11052 15804
rect 11052 15748 11056 15804
rect 10992 15744 11056 15748
rect 11072 15804 11136 15808
rect 11072 15748 11076 15804
rect 11076 15748 11132 15804
rect 11132 15748 11136 15804
rect 11072 15744 11136 15748
rect 11152 15804 11216 15808
rect 11152 15748 11156 15804
rect 11156 15748 11212 15804
rect 11212 15748 11216 15804
rect 11152 15744 11216 15748
rect 11232 15804 11296 15808
rect 11232 15748 11236 15804
rect 11236 15748 11292 15804
rect 11292 15748 11296 15804
rect 11232 15744 11296 15748
rect 18912 15804 18976 15808
rect 18912 15748 18916 15804
rect 18916 15748 18972 15804
rect 18972 15748 18976 15804
rect 18912 15744 18976 15748
rect 18992 15804 19056 15808
rect 18992 15748 18996 15804
rect 18996 15748 19052 15804
rect 19052 15748 19056 15804
rect 18992 15744 19056 15748
rect 19072 15804 19136 15808
rect 19072 15748 19076 15804
rect 19076 15748 19132 15804
rect 19132 15748 19136 15804
rect 19072 15744 19136 15748
rect 19152 15804 19216 15808
rect 19152 15748 19156 15804
rect 19156 15748 19212 15804
rect 19212 15748 19216 15804
rect 19152 15744 19216 15748
rect 19232 15804 19296 15808
rect 19232 15748 19236 15804
rect 19236 15748 19292 15804
rect 19292 15748 19296 15804
rect 19232 15744 19296 15748
rect 26912 15804 26976 15808
rect 26912 15748 26916 15804
rect 26916 15748 26972 15804
rect 26972 15748 26976 15804
rect 26912 15744 26976 15748
rect 26992 15804 27056 15808
rect 26992 15748 26996 15804
rect 26996 15748 27052 15804
rect 27052 15748 27056 15804
rect 26992 15744 27056 15748
rect 27072 15804 27136 15808
rect 27072 15748 27076 15804
rect 27076 15748 27132 15804
rect 27132 15748 27136 15804
rect 27072 15744 27136 15748
rect 27152 15804 27216 15808
rect 27152 15748 27156 15804
rect 27156 15748 27212 15804
rect 27212 15748 27216 15804
rect 27152 15744 27216 15748
rect 27232 15804 27296 15808
rect 27232 15748 27236 15804
rect 27236 15748 27292 15804
rect 27292 15748 27296 15804
rect 27232 15744 27296 15748
rect 11468 15404 11532 15468
rect 3652 15260 3716 15264
rect 3652 15204 3656 15260
rect 3656 15204 3712 15260
rect 3712 15204 3716 15260
rect 3652 15200 3716 15204
rect 3732 15260 3796 15264
rect 3732 15204 3736 15260
rect 3736 15204 3792 15260
rect 3792 15204 3796 15260
rect 3732 15200 3796 15204
rect 3812 15260 3876 15264
rect 3812 15204 3816 15260
rect 3816 15204 3872 15260
rect 3872 15204 3876 15260
rect 3812 15200 3876 15204
rect 3892 15260 3956 15264
rect 3892 15204 3896 15260
rect 3896 15204 3952 15260
rect 3952 15204 3956 15260
rect 3892 15200 3956 15204
rect 3972 15260 4036 15264
rect 3972 15204 3976 15260
rect 3976 15204 4032 15260
rect 4032 15204 4036 15260
rect 3972 15200 4036 15204
rect 11652 15260 11716 15264
rect 11652 15204 11656 15260
rect 11656 15204 11712 15260
rect 11712 15204 11716 15260
rect 11652 15200 11716 15204
rect 11732 15260 11796 15264
rect 11732 15204 11736 15260
rect 11736 15204 11792 15260
rect 11792 15204 11796 15260
rect 11732 15200 11796 15204
rect 11812 15260 11876 15264
rect 11812 15204 11816 15260
rect 11816 15204 11872 15260
rect 11872 15204 11876 15260
rect 11812 15200 11876 15204
rect 11892 15260 11956 15264
rect 11892 15204 11896 15260
rect 11896 15204 11952 15260
rect 11952 15204 11956 15260
rect 11892 15200 11956 15204
rect 11972 15260 12036 15264
rect 11972 15204 11976 15260
rect 11976 15204 12032 15260
rect 12032 15204 12036 15260
rect 11972 15200 12036 15204
rect 19652 15260 19716 15264
rect 19652 15204 19656 15260
rect 19656 15204 19712 15260
rect 19712 15204 19716 15260
rect 19652 15200 19716 15204
rect 19732 15260 19796 15264
rect 19732 15204 19736 15260
rect 19736 15204 19792 15260
rect 19792 15204 19796 15260
rect 19732 15200 19796 15204
rect 19812 15260 19876 15264
rect 19812 15204 19816 15260
rect 19816 15204 19872 15260
rect 19872 15204 19876 15260
rect 19812 15200 19876 15204
rect 19892 15260 19956 15264
rect 19892 15204 19896 15260
rect 19896 15204 19952 15260
rect 19952 15204 19956 15260
rect 19892 15200 19956 15204
rect 19972 15260 20036 15264
rect 19972 15204 19976 15260
rect 19976 15204 20032 15260
rect 20032 15204 20036 15260
rect 19972 15200 20036 15204
rect 27652 15260 27716 15264
rect 27652 15204 27656 15260
rect 27656 15204 27712 15260
rect 27712 15204 27716 15260
rect 27652 15200 27716 15204
rect 27732 15260 27796 15264
rect 27732 15204 27736 15260
rect 27736 15204 27792 15260
rect 27792 15204 27796 15260
rect 27732 15200 27796 15204
rect 27812 15260 27876 15264
rect 27812 15204 27816 15260
rect 27816 15204 27872 15260
rect 27872 15204 27876 15260
rect 27812 15200 27876 15204
rect 27892 15260 27956 15264
rect 27892 15204 27896 15260
rect 27896 15204 27952 15260
rect 27952 15204 27956 15260
rect 27892 15200 27956 15204
rect 27972 15260 28036 15264
rect 27972 15204 27976 15260
rect 27976 15204 28032 15260
rect 28032 15204 28036 15260
rect 27972 15200 28036 15204
rect 2912 14716 2976 14720
rect 2912 14660 2916 14716
rect 2916 14660 2972 14716
rect 2972 14660 2976 14716
rect 2912 14656 2976 14660
rect 2992 14716 3056 14720
rect 2992 14660 2996 14716
rect 2996 14660 3052 14716
rect 3052 14660 3056 14716
rect 2992 14656 3056 14660
rect 3072 14716 3136 14720
rect 3072 14660 3076 14716
rect 3076 14660 3132 14716
rect 3132 14660 3136 14716
rect 3072 14656 3136 14660
rect 3152 14716 3216 14720
rect 3152 14660 3156 14716
rect 3156 14660 3212 14716
rect 3212 14660 3216 14716
rect 3152 14656 3216 14660
rect 3232 14716 3296 14720
rect 3232 14660 3236 14716
rect 3236 14660 3292 14716
rect 3292 14660 3296 14716
rect 3232 14656 3296 14660
rect 10912 14716 10976 14720
rect 10912 14660 10916 14716
rect 10916 14660 10972 14716
rect 10972 14660 10976 14716
rect 10912 14656 10976 14660
rect 10992 14716 11056 14720
rect 10992 14660 10996 14716
rect 10996 14660 11052 14716
rect 11052 14660 11056 14716
rect 10992 14656 11056 14660
rect 11072 14716 11136 14720
rect 11072 14660 11076 14716
rect 11076 14660 11132 14716
rect 11132 14660 11136 14716
rect 11072 14656 11136 14660
rect 11152 14716 11216 14720
rect 11152 14660 11156 14716
rect 11156 14660 11212 14716
rect 11212 14660 11216 14716
rect 11152 14656 11216 14660
rect 11232 14716 11296 14720
rect 11232 14660 11236 14716
rect 11236 14660 11292 14716
rect 11292 14660 11296 14716
rect 11232 14656 11296 14660
rect 18912 14716 18976 14720
rect 18912 14660 18916 14716
rect 18916 14660 18972 14716
rect 18972 14660 18976 14716
rect 18912 14656 18976 14660
rect 18992 14716 19056 14720
rect 18992 14660 18996 14716
rect 18996 14660 19052 14716
rect 19052 14660 19056 14716
rect 18992 14656 19056 14660
rect 19072 14716 19136 14720
rect 19072 14660 19076 14716
rect 19076 14660 19132 14716
rect 19132 14660 19136 14716
rect 19072 14656 19136 14660
rect 19152 14716 19216 14720
rect 19152 14660 19156 14716
rect 19156 14660 19212 14716
rect 19212 14660 19216 14716
rect 19152 14656 19216 14660
rect 19232 14716 19296 14720
rect 19232 14660 19236 14716
rect 19236 14660 19292 14716
rect 19292 14660 19296 14716
rect 19232 14656 19296 14660
rect 26912 14716 26976 14720
rect 26912 14660 26916 14716
rect 26916 14660 26972 14716
rect 26972 14660 26976 14716
rect 26912 14656 26976 14660
rect 26992 14716 27056 14720
rect 26992 14660 26996 14716
rect 26996 14660 27052 14716
rect 27052 14660 27056 14716
rect 26992 14656 27056 14660
rect 27072 14716 27136 14720
rect 27072 14660 27076 14716
rect 27076 14660 27132 14716
rect 27132 14660 27136 14716
rect 27072 14656 27136 14660
rect 27152 14716 27216 14720
rect 27152 14660 27156 14716
rect 27156 14660 27212 14716
rect 27212 14660 27216 14716
rect 27152 14656 27216 14660
rect 27232 14716 27296 14720
rect 27232 14660 27236 14716
rect 27236 14660 27292 14716
rect 27292 14660 27296 14716
rect 27232 14656 27296 14660
rect 3652 14172 3716 14176
rect 3652 14116 3656 14172
rect 3656 14116 3712 14172
rect 3712 14116 3716 14172
rect 3652 14112 3716 14116
rect 3732 14172 3796 14176
rect 3732 14116 3736 14172
rect 3736 14116 3792 14172
rect 3792 14116 3796 14172
rect 3732 14112 3796 14116
rect 3812 14172 3876 14176
rect 3812 14116 3816 14172
rect 3816 14116 3872 14172
rect 3872 14116 3876 14172
rect 3812 14112 3876 14116
rect 3892 14172 3956 14176
rect 3892 14116 3896 14172
rect 3896 14116 3952 14172
rect 3952 14116 3956 14172
rect 3892 14112 3956 14116
rect 3972 14172 4036 14176
rect 3972 14116 3976 14172
rect 3976 14116 4032 14172
rect 4032 14116 4036 14172
rect 3972 14112 4036 14116
rect 11652 14172 11716 14176
rect 11652 14116 11656 14172
rect 11656 14116 11712 14172
rect 11712 14116 11716 14172
rect 11652 14112 11716 14116
rect 11732 14172 11796 14176
rect 11732 14116 11736 14172
rect 11736 14116 11792 14172
rect 11792 14116 11796 14172
rect 11732 14112 11796 14116
rect 11812 14172 11876 14176
rect 11812 14116 11816 14172
rect 11816 14116 11872 14172
rect 11872 14116 11876 14172
rect 11812 14112 11876 14116
rect 11892 14172 11956 14176
rect 11892 14116 11896 14172
rect 11896 14116 11952 14172
rect 11952 14116 11956 14172
rect 11892 14112 11956 14116
rect 11972 14172 12036 14176
rect 11972 14116 11976 14172
rect 11976 14116 12032 14172
rect 12032 14116 12036 14172
rect 11972 14112 12036 14116
rect 19652 14172 19716 14176
rect 19652 14116 19656 14172
rect 19656 14116 19712 14172
rect 19712 14116 19716 14172
rect 19652 14112 19716 14116
rect 19732 14172 19796 14176
rect 19732 14116 19736 14172
rect 19736 14116 19792 14172
rect 19792 14116 19796 14172
rect 19732 14112 19796 14116
rect 19812 14172 19876 14176
rect 19812 14116 19816 14172
rect 19816 14116 19872 14172
rect 19872 14116 19876 14172
rect 19812 14112 19876 14116
rect 19892 14172 19956 14176
rect 19892 14116 19896 14172
rect 19896 14116 19952 14172
rect 19952 14116 19956 14172
rect 19892 14112 19956 14116
rect 19972 14172 20036 14176
rect 19972 14116 19976 14172
rect 19976 14116 20032 14172
rect 20032 14116 20036 14172
rect 19972 14112 20036 14116
rect 27652 14172 27716 14176
rect 27652 14116 27656 14172
rect 27656 14116 27712 14172
rect 27712 14116 27716 14172
rect 27652 14112 27716 14116
rect 27732 14172 27796 14176
rect 27732 14116 27736 14172
rect 27736 14116 27792 14172
rect 27792 14116 27796 14172
rect 27732 14112 27796 14116
rect 27812 14172 27876 14176
rect 27812 14116 27816 14172
rect 27816 14116 27872 14172
rect 27872 14116 27876 14172
rect 27812 14112 27876 14116
rect 27892 14172 27956 14176
rect 27892 14116 27896 14172
rect 27896 14116 27952 14172
rect 27952 14116 27956 14172
rect 27892 14112 27956 14116
rect 27972 14172 28036 14176
rect 27972 14116 27976 14172
rect 27976 14116 28032 14172
rect 28032 14116 28036 14172
rect 27972 14112 28036 14116
rect 2912 13628 2976 13632
rect 2912 13572 2916 13628
rect 2916 13572 2972 13628
rect 2972 13572 2976 13628
rect 2912 13568 2976 13572
rect 2992 13628 3056 13632
rect 2992 13572 2996 13628
rect 2996 13572 3052 13628
rect 3052 13572 3056 13628
rect 2992 13568 3056 13572
rect 3072 13628 3136 13632
rect 3072 13572 3076 13628
rect 3076 13572 3132 13628
rect 3132 13572 3136 13628
rect 3072 13568 3136 13572
rect 3152 13628 3216 13632
rect 3152 13572 3156 13628
rect 3156 13572 3212 13628
rect 3212 13572 3216 13628
rect 3152 13568 3216 13572
rect 3232 13628 3296 13632
rect 3232 13572 3236 13628
rect 3236 13572 3292 13628
rect 3292 13572 3296 13628
rect 3232 13568 3296 13572
rect 10912 13628 10976 13632
rect 10912 13572 10916 13628
rect 10916 13572 10972 13628
rect 10972 13572 10976 13628
rect 10912 13568 10976 13572
rect 10992 13628 11056 13632
rect 10992 13572 10996 13628
rect 10996 13572 11052 13628
rect 11052 13572 11056 13628
rect 10992 13568 11056 13572
rect 11072 13628 11136 13632
rect 11072 13572 11076 13628
rect 11076 13572 11132 13628
rect 11132 13572 11136 13628
rect 11072 13568 11136 13572
rect 11152 13628 11216 13632
rect 11152 13572 11156 13628
rect 11156 13572 11212 13628
rect 11212 13572 11216 13628
rect 11152 13568 11216 13572
rect 11232 13628 11296 13632
rect 11232 13572 11236 13628
rect 11236 13572 11292 13628
rect 11292 13572 11296 13628
rect 11232 13568 11296 13572
rect 18912 13628 18976 13632
rect 18912 13572 18916 13628
rect 18916 13572 18972 13628
rect 18972 13572 18976 13628
rect 18912 13568 18976 13572
rect 18992 13628 19056 13632
rect 18992 13572 18996 13628
rect 18996 13572 19052 13628
rect 19052 13572 19056 13628
rect 18992 13568 19056 13572
rect 19072 13628 19136 13632
rect 19072 13572 19076 13628
rect 19076 13572 19132 13628
rect 19132 13572 19136 13628
rect 19072 13568 19136 13572
rect 19152 13628 19216 13632
rect 19152 13572 19156 13628
rect 19156 13572 19212 13628
rect 19212 13572 19216 13628
rect 19152 13568 19216 13572
rect 19232 13628 19296 13632
rect 19232 13572 19236 13628
rect 19236 13572 19292 13628
rect 19292 13572 19296 13628
rect 19232 13568 19296 13572
rect 26912 13628 26976 13632
rect 26912 13572 26916 13628
rect 26916 13572 26972 13628
rect 26972 13572 26976 13628
rect 26912 13568 26976 13572
rect 26992 13628 27056 13632
rect 26992 13572 26996 13628
rect 26996 13572 27052 13628
rect 27052 13572 27056 13628
rect 26992 13568 27056 13572
rect 27072 13628 27136 13632
rect 27072 13572 27076 13628
rect 27076 13572 27132 13628
rect 27132 13572 27136 13628
rect 27072 13568 27136 13572
rect 27152 13628 27216 13632
rect 27152 13572 27156 13628
rect 27156 13572 27212 13628
rect 27212 13572 27216 13628
rect 27152 13568 27216 13572
rect 27232 13628 27296 13632
rect 27232 13572 27236 13628
rect 27236 13572 27292 13628
rect 27292 13572 27296 13628
rect 27232 13568 27296 13572
rect 3652 13084 3716 13088
rect 3652 13028 3656 13084
rect 3656 13028 3712 13084
rect 3712 13028 3716 13084
rect 3652 13024 3716 13028
rect 3732 13084 3796 13088
rect 3732 13028 3736 13084
rect 3736 13028 3792 13084
rect 3792 13028 3796 13084
rect 3732 13024 3796 13028
rect 3812 13084 3876 13088
rect 3812 13028 3816 13084
rect 3816 13028 3872 13084
rect 3872 13028 3876 13084
rect 3812 13024 3876 13028
rect 3892 13084 3956 13088
rect 3892 13028 3896 13084
rect 3896 13028 3952 13084
rect 3952 13028 3956 13084
rect 3892 13024 3956 13028
rect 3972 13084 4036 13088
rect 3972 13028 3976 13084
rect 3976 13028 4032 13084
rect 4032 13028 4036 13084
rect 3972 13024 4036 13028
rect 11652 13084 11716 13088
rect 11652 13028 11656 13084
rect 11656 13028 11712 13084
rect 11712 13028 11716 13084
rect 11652 13024 11716 13028
rect 11732 13084 11796 13088
rect 11732 13028 11736 13084
rect 11736 13028 11792 13084
rect 11792 13028 11796 13084
rect 11732 13024 11796 13028
rect 11812 13084 11876 13088
rect 11812 13028 11816 13084
rect 11816 13028 11872 13084
rect 11872 13028 11876 13084
rect 11812 13024 11876 13028
rect 11892 13084 11956 13088
rect 11892 13028 11896 13084
rect 11896 13028 11952 13084
rect 11952 13028 11956 13084
rect 11892 13024 11956 13028
rect 11972 13084 12036 13088
rect 11972 13028 11976 13084
rect 11976 13028 12032 13084
rect 12032 13028 12036 13084
rect 11972 13024 12036 13028
rect 19652 13084 19716 13088
rect 19652 13028 19656 13084
rect 19656 13028 19712 13084
rect 19712 13028 19716 13084
rect 19652 13024 19716 13028
rect 19732 13084 19796 13088
rect 19732 13028 19736 13084
rect 19736 13028 19792 13084
rect 19792 13028 19796 13084
rect 19732 13024 19796 13028
rect 19812 13084 19876 13088
rect 19812 13028 19816 13084
rect 19816 13028 19872 13084
rect 19872 13028 19876 13084
rect 19812 13024 19876 13028
rect 19892 13084 19956 13088
rect 19892 13028 19896 13084
rect 19896 13028 19952 13084
rect 19952 13028 19956 13084
rect 19892 13024 19956 13028
rect 19972 13084 20036 13088
rect 19972 13028 19976 13084
rect 19976 13028 20032 13084
rect 20032 13028 20036 13084
rect 19972 13024 20036 13028
rect 27652 13084 27716 13088
rect 27652 13028 27656 13084
rect 27656 13028 27712 13084
rect 27712 13028 27716 13084
rect 27652 13024 27716 13028
rect 27732 13084 27796 13088
rect 27732 13028 27736 13084
rect 27736 13028 27792 13084
rect 27792 13028 27796 13084
rect 27732 13024 27796 13028
rect 27812 13084 27876 13088
rect 27812 13028 27816 13084
rect 27816 13028 27872 13084
rect 27872 13028 27876 13084
rect 27812 13024 27876 13028
rect 27892 13084 27956 13088
rect 27892 13028 27896 13084
rect 27896 13028 27952 13084
rect 27952 13028 27956 13084
rect 27892 13024 27956 13028
rect 27972 13084 28036 13088
rect 27972 13028 27976 13084
rect 27976 13028 28032 13084
rect 28032 13028 28036 13084
rect 27972 13024 28036 13028
rect 2912 12540 2976 12544
rect 2912 12484 2916 12540
rect 2916 12484 2972 12540
rect 2972 12484 2976 12540
rect 2912 12480 2976 12484
rect 2992 12540 3056 12544
rect 2992 12484 2996 12540
rect 2996 12484 3052 12540
rect 3052 12484 3056 12540
rect 2992 12480 3056 12484
rect 3072 12540 3136 12544
rect 3072 12484 3076 12540
rect 3076 12484 3132 12540
rect 3132 12484 3136 12540
rect 3072 12480 3136 12484
rect 3152 12540 3216 12544
rect 3152 12484 3156 12540
rect 3156 12484 3212 12540
rect 3212 12484 3216 12540
rect 3152 12480 3216 12484
rect 3232 12540 3296 12544
rect 3232 12484 3236 12540
rect 3236 12484 3292 12540
rect 3292 12484 3296 12540
rect 3232 12480 3296 12484
rect 10912 12540 10976 12544
rect 10912 12484 10916 12540
rect 10916 12484 10972 12540
rect 10972 12484 10976 12540
rect 10912 12480 10976 12484
rect 10992 12540 11056 12544
rect 10992 12484 10996 12540
rect 10996 12484 11052 12540
rect 11052 12484 11056 12540
rect 10992 12480 11056 12484
rect 11072 12540 11136 12544
rect 11072 12484 11076 12540
rect 11076 12484 11132 12540
rect 11132 12484 11136 12540
rect 11072 12480 11136 12484
rect 11152 12540 11216 12544
rect 11152 12484 11156 12540
rect 11156 12484 11212 12540
rect 11212 12484 11216 12540
rect 11152 12480 11216 12484
rect 11232 12540 11296 12544
rect 11232 12484 11236 12540
rect 11236 12484 11292 12540
rect 11292 12484 11296 12540
rect 11232 12480 11296 12484
rect 18912 12540 18976 12544
rect 18912 12484 18916 12540
rect 18916 12484 18972 12540
rect 18972 12484 18976 12540
rect 18912 12480 18976 12484
rect 18992 12540 19056 12544
rect 18992 12484 18996 12540
rect 18996 12484 19052 12540
rect 19052 12484 19056 12540
rect 18992 12480 19056 12484
rect 19072 12540 19136 12544
rect 19072 12484 19076 12540
rect 19076 12484 19132 12540
rect 19132 12484 19136 12540
rect 19072 12480 19136 12484
rect 19152 12540 19216 12544
rect 19152 12484 19156 12540
rect 19156 12484 19212 12540
rect 19212 12484 19216 12540
rect 19152 12480 19216 12484
rect 19232 12540 19296 12544
rect 19232 12484 19236 12540
rect 19236 12484 19292 12540
rect 19292 12484 19296 12540
rect 19232 12480 19296 12484
rect 26912 12540 26976 12544
rect 26912 12484 26916 12540
rect 26916 12484 26972 12540
rect 26972 12484 26976 12540
rect 26912 12480 26976 12484
rect 26992 12540 27056 12544
rect 26992 12484 26996 12540
rect 26996 12484 27052 12540
rect 27052 12484 27056 12540
rect 26992 12480 27056 12484
rect 27072 12540 27136 12544
rect 27072 12484 27076 12540
rect 27076 12484 27132 12540
rect 27132 12484 27136 12540
rect 27072 12480 27136 12484
rect 27152 12540 27216 12544
rect 27152 12484 27156 12540
rect 27156 12484 27212 12540
rect 27212 12484 27216 12540
rect 27152 12480 27216 12484
rect 27232 12540 27296 12544
rect 27232 12484 27236 12540
rect 27236 12484 27292 12540
rect 27292 12484 27296 12540
rect 27232 12480 27296 12484
rect 3652 11996 3716 12000
rect 3652 11940 3656 11996
rect 3656 11940 3712 11996
rect 3712 11940 3716 11996
rect 3652 11936 3716 11940
rect 3732 11996 3796 12000
rect 3732 11940 3736 11996
rect 3736 11940 3792 11996
rect 3792 11940 3796 11996
rect 3732 11936 3796 11940
rect 3812 11996 3876 12000
rect 3812 11940 3816 11996
rect 3816 11940 3872 11996
rect 3872 11940 3876 11996
rect 3812 11936 3876 11940
rect 3892 11996 3956 12000
rect 3892 11940 3896 11996
rect 3896 11940 3952 11996
rect 3952 11940 3956 11996
rect 3892 11936 3956 11940
rect 3972 11996 4036 12000
rect 3972 11940 3976 11996
rect 3976 11940 4032 11996
rect 4032 11940 4036 11996
rect 3972 11936 4036 11940
rect 11652 11996 11716 12000
rect 11652 11940 11656 11996
rect 11656 11940 11712 11996
rect 11712 11940 11716 11996
rect 11652 11936 11716 11940
rect 11732 11996 11796 12000
rect 11732 11940 11736 11996
rect 11736 11940 11792 11996
rect 11792 11940 11796 11996
rect 11732 11936 11796 11940
rect 11812 11996 11876 12000
rect 11812 11940 11816 11996
rect 11816 11940 11872 11996
rect 11872 11940 11876 11996
rect 11812 11936 11876 11940
rect 11892 11996 11956 12000
rect 11892 11940 11896 11996
rect 11896 11940 11952 11996
rect 11952 11940 11956 11996
rect 11892 11936 11956 11940
rect 11972 11996 12036 12000
rect 11972 11940 11976 11996
rect 11976 11940 12032 11996
rect 12032 11940 12036 11996
rect 11972 11936 12036 11940
rect 19652 11996 19716 12000
rect 19652 11940 19656 11996
rect 19656 11940 19712 11996
rect 19712 11940 19716 11996
rect 19652 11936 19716 11940
rect 19732 11996 19796 12000
rect 19732 11940 19736 11996
rect 19736 11940 19792 11996
rect 19792 11940 19796 11996
rect 19732 11936 19796 11940
rect 19812 11996 19876 12000
rect 19812 11940 19816 11996
rect 19816 11940 19872 11996
rect 19872 11940 19876 11996
rect 19812 11936 19876 11940
rect 19892 11996 19956 12000
rect 19892 11940 19896 11996
rect 19896 11940 19952 11996
rect 19952 11940 19956 11996
rect 19892 11936 19956 11940
rect 19972 11996 20036 12000
rect 19972 11940 19976 11996
rect 19976 11940 20032 11996
rect 20032 11940 20036 11996
rect 19972 11936 20036 11940
rect 27652 11996 27716 12000
rect 27652 11940 27656 11996
rect 27656 11940 27712 11996
rect 27712 11940 27716 11996
rect 27652 11936 27716 11940
rect 27732 11996 27796 12000
rect 27732 11940 27736 11996
rect 27736 11940 27792 11996
rect 27792 11940 27796 11996
rect 27732 11936 27796 11940
rect 27812 11996 27876 12000
rect 27812 11940 27816 11996
rect 27816 11940 27872 11996
rect 27872 11940 27876 11996
rect 27812 11936 27876 11940
rect 27892 11996 27956 12000
rect 27892 11940 27896 11996
rect 27896 11940 27952 11996
rect 27952 11940 27956 11996
rect 27892 11936 27956 11940
rect 27972 11996 28036 12000
rect 27972 11940 27976 11996
rect 27976 11940 28032 11996
rect 28032 11940 28036 11996
rect 27972 11936 28036 11940
rect 2912 11452 2976 11456
rect 2912 11396 2916 11452
rect 2916 11396 2972 11452
rect 2972 11396 2976 11452
rect 2912 11392 2976 11396
rect 2992 11452 3056 11456
rect 2992 11396 2996 11452
rect 2996 11396 3052 11452
rect 3052 11396 3056 11452
rect 2992 11392 3056 11396
rect 3072 11452 3136 11456
rect 3072 11396 3076 11452
rect 3076 11396 3132 11452
rect 3132 11396 3136 11452
rect 3072 11392 3136 11396
rect 3152 11452 3216 11456
rect 3152 11396 3156 11452
rect 3156 11396 3212 11452
rect 3212 11396 3216 11452
rect 3152 11392 3216 11396
rect 3232 11452 3296 11456
rect 3232 11396 3236 11452
rect 3236 11396 3292 11452
rect 3292 11396 3296 11452
rect 3232 11392 3296 11396
rect 10912 11452 10976 11456
rect 10912 11396 10916 11452
rect 10916 11396 10972 11452
rect 10972 11396 10976 11452
rect 10912 11392 10976 11396
rect 10992 11452 11056 11456
rect 10992 11396 10996 11452
rect 10996 11396 11052 11452
rect 11052 11396 11056 11452
rect 10992 11392 11056 11396
rect 11072 11452 11136 11456
rect 11072 11396 11076 11452
rect 11076 11396 11132 11452
rect 11132 11396 11136 11452
rect 11072 11392 11136 11396
rect 11152 11452 11216 11456
rect 11152 11396 11156 11452
rect 11156 11396 11212 11452
rect 11212 11396 11216 11452
rect 11152 11392 11216 11396
rect 11232 11452 11296 11456
rect 11232 11396 11236 11452
rect 11236 11396 11292 11452
rect 11292 11396 11296 11452
rect 11232 11392 11296 11396
rect 18912 11452 18976 11456
rect 18912 11396 18916 11452
rect 18916 11396 18972 11452
rect 18972 11396 18976 11452
rect 18912 11392 18976 11396
rect 18992 11452 19056 11456
rect 18992 11396 18996 11452
rect 18996 11396 19052 11452
rect 19052 11396 19056 11452
rect 18992 11392 19056 11396
rect 19072 11452 19136 11456
rect 19072 11396 19076 11452
rect 19076 11396 19132 11452
rect 19132 11396 19136 11452
rect 19072 11392 19136 11396
rect 19152 11452 19216 11456
rect 19152 11396 19156 11452
rect 19156 11396 19212 11452
rect 19212 11396 19216 11452
rect 19152 11392 19216 11396
rect 19232 11452 19296 11456
rect 19232 11396 19236 11452
rect 19236 11396 19292 11452
rect 19292 11396 19296 11452
rect 19232 11392 19296 11396
rect 26912 11452 26976 11456
rect 26912 11396 26916 11452
rect 26916 11396 26972 11452
rect 26972 11396 26976 11452
rect 26912 11392 26976 11396
rect 26992 11452 27056 11456
rect 26992 11396 26996 11452
rect 26996 11396 27052 11452
rect 27052 11396 27056 11452
rect 26992 11392 27056 11396
rect 27072 11452 27136 11456
rect 27072 11396 27076 11452
rect 27076 11396 27132 11452
rect 27132 11396 27136 11452
rect 27072 11392 27136 11396
rect 27152 11452 27216 11456
rect 27152 11396 27156 11452
rect 27156 11396 27212 11452
rect 27212 11396 27216 11452
rect 27152 11392 27216 11396
rect 27232 11452 27296 11456
rect 27232 11396 27236 11452
rect 27236 11396 27292 11452
rect 27292 11396 27296 11452
rect 27232 11392 27296 11396
rect 3652 10908 3716 10912
rect 3652 10852 3656 10908
rect 3656 10852 3712 10908
rect 3712 10852 3716 10908
rect 3652 10848 3716 10852
rect 3732 10908 3796 10912
rect 3732 10852 3736 10908
rect 3736 10852 3792 10908
rect 3792 10852 3796 10908
rect 3732 10848 3796 10852
rect 3812 10908 3876 10912
rect 3812 10852 3816 10908
rect 3816 10852 3872 10908
rect 3872 10852 3876 10908
rect 3812 10848 3876 10852
rect 3892 10908 3956 10912
rect 3892 10852 3896 10908
rect 3896 10852 3952 10908
rect 3952 10852 3956 10908
rect 3892 10848 3956 10852
rect 3972 10908 4036 10912
rect 3972 10852 3976 10908
rect 3976 10852 4032 10908
rect 4032 10852 4036 10908
rect 3972 10848 4036 10852
rect 11652 10908 11716 10912
rect 11652 10852 11656 10908
rect 11656 10852 11712 10908
rect 11712 10852 11716 10908
rect 11652 10848 11716 10852
rect 11732 10908 11796 10912
rect 11732 10852 11736 10908
rect 11736 10852 11792 10908
rect 11792 10852 11796 10908
rect 11732 10848 11796 10852
rect 11812 10908 11876 10912
rect 11812 10852 11816 10908
rect 11816 10852 11872 10908
rect 11872 10852 11876 10908
rect 11812 10848 11876 10852
rect 11892 10908 11956 10912
rect 11892 10852 11896 10908
rect 11896 10852 11952 10908
rect 11952 10852 11956 10908
rect 11892 10848 11956 10852
rect 11972 10908 12036 10912
rect 11972 10852 11976 10908
rect 11976 10852 12032 10908
rect 12032 10852 12036 10908
rect 11972 10848 12036 10852
rect 19652 10908 19716 10912
rect 19652 10852 19656 10908
rect 19656 10852 19712 10908
rect 19712 10852 19716 10908
rect 19652 10848 19716 10852
rect 19732 10908 19796 10912
rect 19732 10852 19736 10908
rect 19736 10852 19792 10908
rect 19792 10852 19796 10908
rect 19732 10848 19796 10852
rect 19812 10908 19876 10912
rect 19812 10852 19816 10908
rect 19816 10852 19872 10908
rect 19872 10852 19876 10908
rect 19812 10848 19876 10852
rect 19892 10908 19956 10912
rect 19892 10852 19896 10908
rect 19896 10852 19952 10908
rect 19952 10852 19956 10908
rect 19892 10848 19956 10852
rect 19972 10908 20036 10912
rect 19972 10852 19976 10908
rect 19976 10852 20032 10908
rect 20032 10852 20036 10908
rect 19972 10848 20036 10852
rect 27652 10908 27716 10912
rect 27652 10852 27656 10908
rect 27656 10852 27712 10908
rect 27712 10852 27716 10908
rect 27652 10848 27716 10852
rect 27732 10908 27796 10912
rect 27732 10852 27736 10908
rect 27736 10852 27792 10908
rect 27792 10852 27796 10908
rect 27732 10848 27796 10852
rect 27812 10908 27876 10912
rect 27812 10852 27816 10908
rect 27816 10852 27872 10908
rect 27872 10852 27876 10908
rect 27812 10848 27876 10852
rect 27892 10908 27956 10912
rect 27892 10852 27896 10908
rect 27896 10852 27952 10908
rect 27952 10852 27956 10908
rect 27892 10848 27956 10852
rect 27972 10908 28036 10912
rect 27972 10852 27976 10908
rect 27976 10852 28032 10908
rect 28032 10852 28036 10908
rect 27972 10848 28036 10852
rect 11468 10432 11532 10436
rect 11468 10376 11518 10432
rect 11518 10376 11532 10432
rect 11468 10372 11532 10376
rect 2912 10364 2976 10368
rect 2912 10308 2916 10364
rect 2916 10308 2972 10364
rect 2972 10308 2976 10364
rect 2912 10304 2976 10308
rect 2992 10364 3056 10368
rect 2992 10308 2996 10364
rect 2996 10308 3052 10364
rect 3052 10308 3056 10364
rect 2992 10304 3056 10308
rect 3072 10364 3136 10368
rect 3072 10308 3076 10364
rect 3076 10308 3132 10364
rect 3132 10308 3136 10364
rect 3072 10304 3136 10308
rect 3152 10364 3216 10368
rect 3152 10308 3156 10364
rect 3156 10308 3212 10364
rect 3212 10308 3216 10364
rect 3152 10304 3216 10308
rect 3232 10364 3296 10368
rect 3232 10308 3236 10364
rect 3236 10308 3292 10364
rect 3292 10308 3296 10364
rect 3232 10304 3296 10308
rect 10912 10364 10976 10368
rect 10912 10308 10916 10364
rect 10916 10308 10972 10364
rect 10972 10308 10976 10364
rect 10912 10304 10976 10308
rect 10992 10364 11056 10368
rect 10992 10308 10996 10364
rect 10996 10308 11052 10364
rect 11052 10308 11056 10364
rect 10992 10304 11056 10308
rect 11072 10364 11136 10368
rect 11072 10308 11076 10364
rect 11076 10308 11132 10364
rect 11132 10308 11136 10364
rect 11072 10304 11136 10308
rect 11152 10364 11216 10368
rect 11152 10308 11156 10364
rect 11156 10308 11212 10364
rect 11212 10308 11216 10364
rect 11152 10304 11216 10308
rect 11232 10364 11296 10368
rect 11232 10308 11236 10364
rect 11236 10308 11292 10364
rect 11292 10308 11296 10364
rect 11232 10304 11296 10308
rect 18912 10364 18976 10368
rect 18912 10308 18916 10364
rect 18916 10308 18972 10364
rect 18972 10308 18976 10364
rect 18912 10304 18976 10308
rect 18992 10364 19056 10368
rect 18992 10308 18996 10364
rect 18996 10308 19052 10364
rect 19052 10308 19056 10364
rect 18992 10304 19056 10308
rect 19072 10364 19136 10368
rect 19072 10308 19076 10364
rect 19076 10308 19132 10364
rect 19132 10308 19136 10364
rect 19072 10304 19136 10308
rect 19152 10364 19216 10368
rect 19152 10308 19156 10364
rect 19156 10308 19212 10364
rect 19212 10308 19216 10364
rect 19152 10304 19216 10308
rect 19232 10364 19296 10368
rect 19232 10308 19236 10364
rect 19236 10308 19292 10364
rect 19292 10308 19296 10364
rect 19232 10304 19296 10308
rect 26912 10364 26976 10368
rect 26912 10308 26916 10364
rect 26916 10308 26972 10364
rect 26972 10308 26976 10364
rect 26912 10304 26976 10308
rect 26992 10364 27056 10368
rect 26992 10308 26996 10364
rect 26996 10308 27052 10364
rect 27052 10308 27056 10364
rect 26992 10304 27056 10308
rect 27072 10364 27136 10368
rect 27072 10308 27076 10364
rect 27076 10308 27132 10364
rect 27132 10308 27136 10364
rect 27072 10304 27136 10308
rect 27152 10364 27216 10368
rect 27152 10308 27156 10364
rect 27156 10308 27212 10364
rect 27212 10308 27216 10364
rect 27152 10304 27216 10308
rect 27232 10364 27296 10368
rect 27232 10308 27236 10364
rect 27236 10308 27292 10364
rect 27292 10308 27296 10364
rect 27232 10304 27296 10308
rect 3652 9820 3716 9824
rect 3652 9764 3656 9820
rect 3656 9764 3712 9820
rect 3712 9764 3716 9820
rect 3652 9760 3716 9764
rect 3732 9820 3796 9824
rect 3732 9764 3736 9820
rect 3736 9764 3792 9820
rect 3792 9764 3796 9820
rect 3732 9760 3796 9764
rect 3812 9820 3876 9824
rect 3812 9764 3816 9820
rect 3816 9764 3872 9820
rect 3872 9764 3876 9820
rect 3812 9760 3876 9764
rect 3892 9820 3956 9824
rect 3892 9764 3896 9820
rect 3896 9764 3952 9820
rect 3952 9764 3956 9820
rect 3892 9760 3956 9764
rect 3972 9820 4036 9824
rect 3972 9764 3976 9820
rect 3976 9764 4032 9820
rect 4032 9764 4036 9820
rect 3972 9760 4036 9764
rect 11652 9820 11716 9824
rect 11652 9764 11656 9820
rect 11656 9764 11712 9820
rect 11712 9764 11716 9820
rect 11652 9760 11716 9764
rect 11732 9820 11796 9824
rect 11732 9764 11736 9820
rect 11736 9764 11792 9820
rect 11792 9764 11796 9820
rect 11732 9760 11796 9764
rect 11812 9820 11876 9824
rect 11812 9764 11816 9820
rect 11816 9764 11872 9820
rect 11872 9764 11876 9820
rect 11812 9760 11876 9764
rect 11892 9820 11956 9824
rect 11892 9764 11896 9820
rect 11896 9764 11952 9820
rect 11952 9764 11956 9820
rect 11892 9760 11956 9764
rect 11972 9820 12036 9824
rect 11972 9764 11976 9820
rect 11976 9764 12032 9820
rect 12032 9764 12036 9820
rect 11972 9760 12036 9764
rect 19652 9820 19716 9824
rect 19652 9764 19656 9820
rect 19656 9764 19712 9820
rect 19712 9764 19716 9820
rect 19652 9760 19716 9764
rect 19732 9820 19796 9824
rect 19732 9764 19736 9820
rect 19736 9764 19792 9820
rect 19792 9764 19796 9820
rect 19732 9760 19796 9764
rect 19812 9820 19876 9824
rect 19812 9764 19816 9820
rect 19816 9764 19872 9820
rect 19872 9764 19876 9820
rect 19812 9760 19876 9764
rect 19892 9820 19956 9824
rect 19892 9764 19896 9820
rect 19896 9764 19952 9820
rect 19952 9764 19956 9820
rect 19892 9760 19956 9764
rect 19972 9820 20036 9824
rect 19972 9764 19976 9820
rect 19976 9764 20032 9820
rect 20032 9764 20036 9820
rect 19972 9760 20036 9764
rect 27652 9820 27716 9824
rect 27652 9764 27656 9820
rect 27656 9764 27712 9820
rect 27712 9764 27716 9820
rect 27652 9760 27716 9764
rect 27732 9820 27796 9824
rect 27732 9764 27736 9820
rect 27736 9764 27792 9820
rect 27792 9764 27796 9820
rect 27732 9760 27796 9764
rect 27812 9820 27876 9824
rect 27812 9764 27816 9820
rect 27816 9764 27872 9820
rect 27872 9764 27876 9820
rect 27812 9760 27876 9764
rect 27892 9820 27956 9824
rect 27892 9764 27896 9820
rect 27896 9764 27952 9820
rect 27952 9764 27956 9820
rect 27892 9760 27956 9764
rect 27972 9820 28036 9824
rect 27972 9764 27976 9820
rect 27976 9764 28032 9820
rect 28032 9764 28036 9820
rect 27972 9760 28036 9764
rect 2912 9276 2976 9280
rect 2912 9220 2916 9276
rect 2916 9220 2972 9276
rect 2972 9220 2976 9276
rect 2912 9216 2976 9220
rect 2992 9276 3056 9280
rect 2992 9220 2996 9276
rect 2996 9220 3052 9276
rect 3052 9220 3056 9276
rect 2992 9216 3056 9220
rect 3072 9276 3136 9280
rect 3072 9220 3076 9276
rect 3076 9220 3132 9276
rect 3132 9220 3136 9276
rect 3072 9216 3136 9220
rect 3152 9276 3216 9280
rect 3152 9220 3156 9276
rect 3156 9220 3212 9276
rect 3212 9220 3216 9276
rect 3152 9216 3216 9220
rect 3232 9276 3296 9280
rect 3232 9220 3236 9276
rect 3236 9220 3292 9276
rect 3292 9220 3296 9276
rect 3232 9216 3296 9220
rect 10912 9276 10976 9280
rect 10912 9220 10916 9276
rect 10916 9220 10972 9276
rect 10972 9220 10976 9276
rect 10912 9216 10976 9220
rect 10992 9276 11056 9280
rect 10992 9220 10996 9276
rect 10996 9220 11052 9276
rect 11052 9220 11056 9276
rect 10992 9216 11056 9220
rect 11072 9276 11136 9280
rect 11072 9220 11076 9276
rect 11076 9220 11132 9276
rect 11132 9220 11136 9276
rect 11072 9216 11136 9220
rect 11152 9276 11216 9280
rect 11152 9220 11156 9276
rect 11156 9220 11212 9276
rect 11212 9220 11216 9276
rect 11152 9216 11216 9220
rect 11232 9276 11296 9280
rect 11232 9220 11236 9276
rect 11236 9220 11292 9276
rect 11292 9220 11296 9276
rect 11232 9216 11296 9220
rect 18912 9276 18976 9280
rect 18912 9220 18916 9276
rect 18916 9220 18972 9276
rect 18972 9220 18976 9276
rect 18912 9216 18976 9220
rect 18992 9276 19056 9280
rect 18992 9220 18996 9276
rect 18996 9220 19052 9276
rect 19052 9220 19056 9276
rect 18992 9216 19056 9220
rect 19072 9276 19136 9280
rect 19072 9220 19076 9276
rect 19076 9220 19132 9276
rect 19132 9220 19136 9276
rect 19072 9216 19136 9220
rect 19152 9276 19216 9280
rect 19152 9220 19156 9276
rect 19156 9220 19212 9276
rect 19212 9220 19216 9276
rect 19152 9216 19216 9220
rect 19232 9276 19296 9280
rect 19232 9220 19236 9276
rect 19236 9220 19292 9276
rect 19292 9220 19296 9276
rect 19232 9216 19296 9220
rect 26912 9276 26976 9280
rect 26912 9220 26916 9276
rect 26916 9220 26972 9276
rect 26972 9220 26976 9276
rect 26912 9216 26976 9220
rect 26992 9276 27056 9280
rect 26992 9220 26996 9276
rect 26996 9220 27052 9276
rect 27052 9220 27056 9276
rect 26992 9216 27056 9220
rect 27072 9276 27136 9280
rect 27072 9220 27076 9276
rect 27076 9220 27132 9276
rect 27132 9220 27136 9276
rect 27072 9216 27136 9220
rect 27152 9276 27216 9280
rect 27152 9220 27156 9276
rect 27156 9220 27212 9276
rect 27212 9220 27216 9276
rect 27152 9216 27216 9220
rect 27232 9276 27296 9280
rect 27232 9220 27236 9276
rect 27236 9220 27292 9276
rect 27292 9220 27296 9276
rect 27232 9216 27296 9220
rect 3652 8732 3716 8736
rect 3652 8676 3656 8732
rect 3656 8676 3712 8732
rect 3712 8676 3716 8732
rect 3652 8672 3716 8676
rect 3732 8732 3796 8736
rect 3732 8676 3736 8732
rect 3736 8676 3792 8732
rect 3792 8676 3796 8732
rect 3732 8672 3796 8676
rect 3812 8732 3876 8736
rect 3812 8676 3816 8732
rect 3816 8676 3872 8732
rect 3872 8676 3876 8732
rect 3812 8672 3876 8676
rect 3892 8732 3956 8736
rect 3892 8676 3896 8732
rect 3896 8676 3952 8732
rect 3952 8676 3956 8732
rect 3892 8672 3956 8676
rect 3972 8732 4036 8736
rect 3972 8676 3976 8732
rect 3976 8676 4032 8732
rect 4032 8676 4036 8732
rect 3972 8672 4036 8676
rect 11652 8732 11716 8736
rect 11652 8676 11656 8732
rect 11656 8676 11712 8732
rect 11712 8676 11716 8732
rect 11652 8672 11716 8676
rect 11732 8732 11796 8736
rect 11732 8676 11736 8732
rect 11736 8676 11792 8732
rect 11792 8676 11796 8732
rect 11732 8672 11796 8676
rect 11812 8732 11876 8736
rect 11812 8676 11816 8732
rect 11816 8676 11872 8732
rect 11872 8676 11876 8732
rect 11812 8672 11876 8676
rect 11892 8732 11956 8736
rect 11892 8676 11896 8732
rect 11896 8676 11952 8732
rect 11952 8676 11956 8732
rect 11892 8672 11956 8676
rect 11972 8732 12036 8736
rect 11972 8676 11976 8732
rect 11976 8676 12032 8732
rect 12032 8676 12036 8732
rect 11972 8672 12036 8676
rect 19652 8732 19716 8736
rect 19652 8676 19656 8732
rect 19656 8676 19712 8732
rect 19712 8676 19716 8732
rect 19652 8672 19716 8676
rect 19732 8732 19796 8736
rect 19732 8676 19736 8732
rect 19736 8676 19792 8732
rect 19792 8676 19796 8732
rect 19732 8672 19796 8676
rect 19812 8732 19876 8736
rect 19812 8676 19816 8732
rect 19816 8676 19872 8732
rect 19872 8676 19876 8732
rect 19812 8672 19876 8676
rect 19892 8732 19956 8736
rect 19892 8676 19896 8732
rect 19896 8676 19952 8732
rect 19952 8676 19956 8732
rect 19892 8672 19956 8676
rect 19972 8732 20036 8736
rect 19972 8676 19976 8732
rect 19976 8676 20032 8732
rect 20032 8676 20036 8732
rect 19972 8672 20036 8676
rect 27652 8732 27716 8736
rect 27652 8676 27656 8732
rect 27656 8676 27712 8732
rect 27712 8676 27716 8732
rect 27652 8672 27716 8676
rect 27732 8732 27796 8736
rect 27732 8676 27736 8732
rect 27736 8676 27792 8732
rect 27792 8676 27796 8732
rect 27732 8672 27796 8676
rect 27812 8732 27876 8736
rect 27812 8676 27816 8732
rect 27816 8676 27872 8732
rect 27872 8676 27876 8732
rect 27812 8672 27876 8676
rect 27892 8732 27956 8736
rect 27892 8676 27896 8732
rect 27896 8676 27952 8732
rect 27952 8676 27956 8732
rect 27892 8672 27956 8676
rect 27972 8732 28036 8736
rect 27972 8676 27976 8732
rect 27976 8676 28032 8732
rect 28032 8676 28036 8732
rect 27972 8672 28036 8676
rect 2912 8188 2976 8192
rect 2912 8132 2916 8188
rect 2916 8132 2972 8188
rect 2972 8132 2976 8188
rect 2912 8128 2976 8132
rect 2992 8188 3056 8192
rect 2992 8132 2996 8188
rect 2996 8132 3052 8188
rect 3052 8132 3056 8188
rect 2992 8128 3056 8132
rect 3072 8188 3136 8192
rect 3072 8132 3076 8188
rect 3076 8132 3132 8188
rect 3132 8132 3136 8188
rect 3072 8128 3136 8132
rect 3152 8188 3216 8192
rect 3152 8132 3156 8188
rect 3156 8132 3212 8188
rect 3212 8132 3216 8188
rect 3152 8128 3216 8132
rect 3232 8188 3296 8192
rect 3232 8132 3236 8188
rect 3236 8132 3292 8188
rect 3292 8132 3296 8188
rect 3232 8128 3296 8132
rect 10912 8188 10976 8192
rect 10912 8132 10916 8188
rect 10916 8132 10972 8188
rect 10972 8132 10976 8188
rect 10912 8128 10976 8132
rect 10992 8188 11056 8192
rect 10992 8132 10996 8188
rect 10996 8132 11052 8188
rect 11052 8132 11056 8188
rect 10992 8128 11056 8132
rect 11072 8188 11136 8192
rect 11072 8132 11076 8188
rect 11076 8132 11132 8188
rect 11132 8132 11136 8188
rect 11072 8128 11136 8132
rect 11152 8188 11216 8192
rect 11152 8132 11156 8188
rect 11156 8132 11212 8188
rect 11212 8132 11216 8188
rect 11152 8128 11216 8132
rect 11232 8188 11296 8192
rect 11232 8132 11236 8188
rect 11236 8132 11292 8188
rect 11292 8132 11296 8188
rect 11232 8128 11296 8132
rect 18912 8188 18976 8192
rect 18912 8132 18916 8188
rect 18916 8132 18972 8188
rect 18972 8132 18976 8188
rect 18912 8128 18976 8132
rect 18992 8188 19056 8192
rect 18992 8132 18996 8188
rect 18996 8132 19052 8188
rect 19052 8132 19056 8188
rect 18992 8128 19056 8132
rect 19072 8188 19136 8192
rect 19072 8132 19076 8188
rect 19076 8132 19132 8188
rect 19132 8132 19136 8188
rect 19072 8128 19136 8132
rect 19152 8188 19216 8192
rect 19152 8132 19156 8188
rect 19156 8132 19212 8188
rect 19212 8132 19216 8188
rect 19152 8128 19216 8132
rect 19232 8188 19296 8192
rect 19232 8132 19236 8188
rect 19236 8132 19292 8188
rect 19292 8132 19296 8188
rect 19232 8128 19296 8132
rect 26912 8188 26976 8192
rect 26912 8132 26916 8188
rect 26916 8132 26972 8188
rect 26972 8132 26976 8188
rect 26912 8128 26976 8132
rect 26992 8188 27056 8192
rect 26992 8132 26996 8188
rect 26996 8132 27052 8188
rect 27052 8132 27056 8188
rect 26992 8128 27056 8132
rect 27072 8188 27136 8192
rect 27072 8132 27076 8188
rect 27076 8132 27132 8188
rect 27132 8132 27136 8188
rect 27072 8128 27136 8132
rect 27152 8188 27216 8192
rect 27152 8132 27156 8188
rect 27156 8132 27212 8188
rect 27212 8132 27216 8188
rect 27152 8128 27216 8132
rect 27232 8188 27296 8192
rect 27232 8132 27236 8188
rect 27236 8132 27292 8188
rect 27292 8132 27296 8188
rect 27232 8128 27296 8132
rect 3652 7644 3716 7648
rect 3652 7588 3656 7644
rect 3656 7588 3712 7644
rect 3712 7588 3716 7644
rect 3652 7584 3716 7588
rect 3732 7644 3796 7648
rect 3732 7588 3736 7644
rect 3736 7588 3792 7644
rect 3792 7588 3796 7644
rect 3732 7584 3796 7588
rect 3812 7644 3876 7648
rect 3812 7588 3816 7644
rect 3816 7588 3872 7644
rect 3872 7588 3876 7644
rect 3812 7584 3876 7588
rect 3892 7644 3956 7648
rect 3892 7588 3896 7644
rect 3896 7588 3952 7644
rect 3952 7588 3956 7644
rect 3892 7584 3956 7588
rect 3972 7644 4036 7648
rect 3972 7588 3976 7644
rect 3976 7588 4032 7644
rect 4032 7588 4036 7644
rect 3972 7584 4036 7588
rect 11652 7644 11716 7648
rect 11652 7588 11656 7644
rect 11656 7588 11712 7644
rect 11712 7588 11716 7644
rect 11652 7584 11716 7588
rect 11732 7644 11796 7648
rect 11732 7588 11736 7644
rect 11736 7588 11792 7644
rect 11792 7588 11796 7644
rect 11732 7584 11796 7588
rect 11812 7644 11876 7648
rect 11812 7588 11816 7644
rect 11816 7588 11872 7644
rect 11872 7588 11876 7644
rect 11812 7584 11876 7588
rect 11892 7644 11956 7648
rect 11892 7588 11896 7644
rect 11896 7588 11952 7644
rect 11952 7588 11956 7644
rect 11892 7584 11956 7588
rect 11972 7644 12036 7648
rect 11972 7588 11976 7644
rect 11976 7588 12032 7644
rect 12032 7588 12036 7644
rect 11972 7584 12036 7588
rect 19652 7644 19716 7648
rect 19652 7588 19656 7644
rect 19656 7588 19712 7644
rect 19712 7588 19716 7644
rect 19652 7584 19716 7588
rect 19732 7644 19796 7648
rect 19732 7588 19736 7644
rect 19736 7588 19792 7644
rect 19792 7588 19796 7644
rect 19732 7584 19796 7588
rect 19812 7644 19876 7648
rect 19812 7588 19816 7644
rect 19816 7588 19872 7644
rect 19872 7588 19876 7644
rect 19812 7584 19876 7588
rect 19892 7644 19956 7648
rect 19892 7588 19896 7644
rect 19896 7588 19952 7644
rect 19952 7588 19956 7644
rect 19892 7584 19956 7588
rect 19972 7644 20036 7648
rect 19972 7588 19976 7644
rect 19976 7588 20032 7644
rect 20032 7588 20036 7644
rect 19972 7584 20036 7588
rect 27652 7644 27716 7648
rect 27652 7588 27656 7644
rect 27656 7588 27712 7644
rect 27712 7588 27716 7644
rect 27652 7584 27716 7588
rect 27732 7644 27796 7648
rect 27732 7588 27736 7644
rect 27736 7588 27792 7644
rect 27792 7588 27796 7644
rect 27732 7584 27796 7588
rect 27812 7644 27876 7648
rect 27812 7588 27816 7644
rect 27816 7588 27872 7644
rect 27872 7588 27876 7644
rect 27812 7584 27876 7588
rect 27892 7644 27956 7648
rect 27892 7588 27896 7644
rect 27896 7588 27952 7644
rect 27952 7588 27956 7644
rect 27892 7584 27956 7588
rect 27972 7644 28036 7648
rect 27972 7588 27976 7644
rect 27976 7588 28032 7644
rect 28032 7588 28036 7644
rect 27972 7584 28036 7588
rect 2912 7100 2976 7104
rect 2912 7044 2916 7100
rect 2916 7044 2972 7100
rect 2972 7044 2976 7100
rect 2912 7040 2976 7044
rect 2992 7100 3056 7104
rect 2992 7044 2996 7100
rect 2996 7044 3052 7100
rect 3052 7044 3056 7100
rect 2992 7040 3056 7044
rect 3072 7100 3136 7104
rect 3072 7044 3076 7100
rect 3076 7044 3132 7100
rect 3132 7044 3136 7100
rect 3072 7040 3136 7044
rect 3152 7100 3216 7104
rect 3152 7044 3156 7100
rect 3156 7044 3212 7100
rect 3212 7044 3216 7100
rect 3152 7040 3216 7044
rect 3232 7100 3296 7104
rect 3232 7044 3236 7100
rect 3236 7044 3292 7100
rect 3292 7044 3296 7100
rect 3232 7040 3296 7044
rect 10912 7100 10976 7104
rect 10912 7044 10916 7100
rect 10916 7044 10972 7100
rect 10972 7044 10976 7100
rect 10912 7040 10976 7044
rect 10992 7100 11056 7104
rect 10992 7044 10996 7100
rect 10996 7044 11052 7100
rect 11052 7044 11056 7100
rect 10992 7040 11056 7044
rect 11072 7100 11136 7104
rect 11072 7044 11076 7100
rect 11076 7044 11132 7100
rect 11132 7044 11136 7100
rect 11072 7040 11136 7044
rect 11152 7100 11216 7104
rect 11152 7044 11156 7100
rect 11156 7044 11212 7100
rect 11212 7044 11216 7100
rect 11152 7040 11216 7044
rect 11232 7100 11296 7104
rect 11232 7044 11236 7100
rect 11236 7044 11292 7100
rect 11292 7044 11296 7100
rect 11232 7040 11296 7044
rect 18912 7100 18976 7104
rect 18912 7044 18916 7100
rect 18916 7044 18972 7100
rect 18972 7044 18976 7100
rect 18912 7040 18976 7044
rect 18992 7100 19056 7104
rect 18992 7044 18996 7100
rect 18996 7044 19052 7100
rect 19052 7044 19056 7100
rect 18992 7040 19056 7044
rect 19072 7100 19136 7104
rect 19072 7044 19076 7100
rect 19076 7044 19132 7100
rect 19132 7044 19136 7100
rect 19072 7040 19136 7044
rect 19152 7100 19216 7104
rect 19152 7044 19156 7100
rect 19156 7044 19212 7100
rect 19212 7044 19216 7100
rect 19152 7040 19216 7044
rect 19232 7100 19296 7104
rect 19232 7044 19236 7100
rect 19236 7044 19292 7100
rect 19292 7044 19296 7100
rect 19232 7040 19296 7044
rect 26912 7100 26976 7104
rect 26912 7044 26916 7100
rect 26916 7044 26972 7100
rect 26972 7044 26976 7100
rect 26912 7040 26976 7044
rect 26992 7100 27056 7104
rect 26992 7044 26996 7100
rect 26996 7044 27052 7100
rect 27052 7044 27056 7100
rect 26992 7040 27056 7044
rect 27072 7100 27136 7104
rect 27072 7044 27076 7100
rect 27076 7044 27132 7100
rect 27132 7044 27136 7100
rect 27072 7040 27136 7044
rect 27152 7100 27216 7104
rect 27152 7044 27156 7100
rect 27156 7044 27212 7100
rect 27212 7044 27216 7100
rect 27152 7040 27216 7044
rect 27232 7100 27296 7104
rect 27232 7044 27236 7100
rect 27236 7044 27292 7100
rect 27292 7044 27296 7100
rect 27232 7040 27296 7044
rect 3652 6556 3716 6560
rect 3652 6500 3656 6556
rect 3656 6500 3712 6556
rect 3712 6500 3716 6556
rect 3652 6496 3716 6500
rect 3732 6556 3796 6560
rect 3732 6500 3736 6556
rect 3736 6500 3792 6556
rect 3792 6500 3796 6556
rect 3732 6496 3796 6500
rect 3812 6556 3876 6560
rect 3812 6500 3816 6556
rect 3816 6500 3872 6556
rect 3872 6500 3876 6556
rect 3812 6496 3876 6500
rect 3892 6556 3956 6560
rect 3892 6500 3896 6556
rect 3896 6500 3952 6556
rect 3952 6500 3956 6556
rect 3892 6496 3956 6500
rect 3972 6556 4036 6560
rect 3972 6500 3976 6556
rect 3976 6500 4032 6556
rect 4032 6500 4036 6556
rect 3972 6496 4036 6500
rect 11652 6556 11716 6560
rect 11652 6500 11656 6556
rect 11656 6500 11712 6556
rect 11712 6500 11716 6556
rect 11652 6496 11716 6500
rect 11732 6556 11796 6560
rect 11732 6500 11736 6556
rect 11736 6500 11792 6556
rect 11792 6500 11796 6556
rect 11732 6496 11796 6500
rect 11812 6556 11876 6560
rect 11812 6500 11816 6556
rect 11816 6500 11872 6556
rect 11872 6500 11876 6556
rect 11812 6496 11876 6500
rect 11892 6556 11956 6560
rect 11892 6500 11896 6556
rect 11896 6500 11952 6556
rect 11952 6500 11956 6556
rect 11892 6496 11956 6500
rect 11972 6556 12036 6560
rect 11972 6500 11976 6556
rect 11976 6500 12032 6556
rect 12032 6500 12036 6556
rect 11972 6496 12036 6500
rect 19652 6556 19716 6560
rect 19652 6500 19656 6556
rect 19656 6500 19712 6556
rect 19712 6500 19716 6556
rect 19652 6496 19716 6500
rect 19732 6556 19796 6560
rect 19732 6500 19736 6556
rect 19736 6500 19792 6556
rect 19792 6500 19796 6556
rect 19732 6496 19796 6500
rect 19812 6556 19876 6560
rect 19812 6500 19816 6556
rect 19816 6500 19872 6556
rect 19872 6500 19876 6556
rect 19812 6496 19876 6500
rect 19892 6556 19956 6560
rect 19892 6500 19896 6556
rect 19896 6500 19952 6556
rect 19952 6500 19956 6556
rect 19892 6496 19956 6500
rect 19972 6556 20036 6560
rect 19972 6500 19976 6556
rect 19976 6500 20032 6556
rect 20032 6500 20036 6556
rect 19972 6496 20036 6500
rect 27652 6556 27716 6560
rect 27652 6500 27656 6556
rect 27656 6500 27712 6556
rect 27712 6500 27716 6556
rect 27652 6496 27716 6500
rect 27732 6556 27796 6560
rect 27732 6500 27736 6556
rect 27736 6500 27792 6556
rect 27792 6500 27796 6556
rect 27732 6496 27796 6500
rect 27812 6556 27876 6560
rect 27812 6500 27816 6556
rect 27816 6500 27872 6556
rect 27872 6500 27876 6556
rect 27812 6496 27876 6500
rect 27892 6556 27956 6560
rect 27892 6500 27896 6556
rect 27896 6500 27952 6556
rect 27952 6500 27956 6556
rect 27892 6496 27956 6500
rect 27972 6556 28036 6560
rect 27972 6500 27976 6556
rect 27976 6500 28032 6556
rect 28032 6500 28036 6556
rect 27972 6496 28036 6500
rect 2912 6012 2976 6016
rect 2912 5956 2916 6012
rect 2916 5956 2972 6012
rect 2972 5956 2976 6012
rect 2912 5952 2976 5956
rect 2992 6012 3056 6016
rect 2992 5956 2996 6012
rect 2996 5956 3052 6012
rect 3052 5956 3056 6012
rect 2992 5952 3056 5956
rect 3072 6012 3136 6016
rect 3072 5956 3076 6012
rect 3076 5956 3132 6012
rect 3132 5956 3136 6012
rect 3072 5952 3136 5956
rect 3152 6012 3216 6016
rect 3152 5956 3156 6012
rect 3156 5956 3212 6012
rect 3212 5956 3216 6012
rect 3152 5952 3216 5956
rect 3232 6012 3296 6016
rect 3232 5956 3236 6012
rect 3236 5956 3292 6012
rect 3292 5956 3296 6012
rect 3232 5952 3296 5956
rect 10912 6012 10976 6016
rect 10912 5956 10916 6012
rect 10916 5956 10972 6012
rect 10972 5956 10976 6012
rect 10912 5952 10976 5956
rect 10992 6012 11056 6016
rect 10992 5956 10996 6012
rect 10996 5956 11052 6012
rect 11052 5956 11056 6012
rect 10992 5952 11056 5956
rect 11072 6012 11136 6016
rect 11072 5956 11076 6012
rect 11076 5956 11132 6012
rect 11132 5956 11136 6012
rect 11072 5952 11136 5956
rect 11152 6012 11216 6016
rect 11152 5956 11156 6012
rect 11156 5956 11212 6012
rect 11212 5956 11216 6012
rect 11152 5952 11216 5956
rect 11232 6012 11296 6016
rect 11232 5956 11236 6012
rect 11236 5956 11292 6012
rect 11292 5956 11296 6012
rect 11232 5952 11296 5956
rect 18912 6012 18976 6016
rect 18912 5956 18916 6012
rect 18916 5956 18972 6012
rect 18972 5956 18976 6012
rect 18912 5952 18976 5956
rect 18992 6012 19056 6016
rect 18992 5956 18996 6012
rect 18996 5956 19052 6012
rect 19052 5956 19056 6012
rect 18992 5952 19056 5956
rect 19072 6012 19136 6016
rect 19072 5956 19076 6012
rect 19076 5956 19132 6012
rect 19132 5956 19136 6012
rect 19072 5952 19136 5956
rect 19152 6012 19216 6016
rect 19152 5956 19156 6012
rect 19156 5956 19212 6012
rect 19212 5956 19216 6012
rect 19152 5952 19216 5956
rect 19232 6012 19296 6016
rect 19232 5956 19236 6012
rect 19236 5956 19292 6012
rect 19292 5956 19296 6012
rect 19232 5952 19296 5956
rect 26912 6012 26976 6016
rect 26912 5956 26916 6012
rect 26916 5956 26972 6012
rect 26972 5956 26976 6012
rect 26912 5952 26976 5956
rect 26992 6012 27056 6016
rect 26992 5956 26996 6012
rect 26996 5956 27052 6012
rect 27052 5956 27056 6012
rect 26992 5952 27056 5956
rect 27072 6012 27136 6016
rect 27072 5956 27076 6012
rect 27076 5956 27132 6012
rect 27132 5956 27136 6012
rect 27072 5952 27136 5956
rect 27152 6012 27216 6016
rect 27152 5956 27156 6012
rect 27156 5956 27212 6012
rect 27212 5956 27216 6012
rect 27152 5952 27216 5956
rect 27232 6012 27296 6016
rect 27232 5956 27236 6012
rect 27236 5956 27292 6012
rect 27292 5956 27296 6012
rect 27232 5952 27296 5956
rect 3652 5468 3716 5472
rect 3652 5412 3656 5468
rect 3656 5412 3712 5468
rect 3712 5412 3716 5468
rect 3652 5408 3716 5412
rect 3732 5468 3796 5472
rect 3732 5412 3736 5468
rect 3736 5412 3792 5468
rect 3792 5412 3796 5468
rect 3732 5408 3796 5412
rect 3812 5468 3876 5472
rect 3812 5412 3816 5468
rect 3816 5412 3872 5468
rect 3872 5412 3876 5468
rect 3812 5408 3876 5412
rect 3892 5468 3956 5472
rect 3892 5412 3896 5468
rect 3896 5412 3952 5468
rect 3952 5412 3956 5468
rect 3892 5408 3956 5412
rect 3972 5468 4036 5472
rect 3972 5412 3976 5468
rect 3976 5412 4032 5468
rect 4032 5412 4036 5468
rect 3972 5408 4036 5412
rect 11652 5468 11716 5472
rect 11652 5412 11656 5468
rect 11656 5412 11712 5468
rect 11712 5412 11716 5468
rect 11652 5408 11716 5412
rect 11732 5468 11796 5472
rect 11732 5412 11736 5468
rect 11736 5412 11792 5468
rect 11792 5412 11796 5468
rect 11732 5408 11796 5412
rect 11812 5468 11876 5472
rect 11812 5412 11816 5468
rect 11816 5412 11872 5468
rect 11872 5412 11876 5468
rect 11812 5408 11876 5412
rect 11892 5468 11956 5472
rect 11892 5412 11896 5468
rect 11896 5412 11952 5468
rect 11952 5412 11956 5468
rect 11892 5408 11956 5412
rect 11972 5468 12036 5472
rect 11972 5412 11976 5468
rect 11976 5412 12032 5468
rect 12032 5412 12036 5468
rect 11972 5408 12036 5412
rect 19652 5468 19716 5472
rect 19652 5412 19656 5468
rect 19656 5412 19712 5468
rect 19712 5412 19716 5468
rect 19652 5408 19716 5412
rect 19732 5468 19796 5472
rect 19732 5412 19736 5468
rect 19736 5412 19792 5468
rect 19792 5412 19796 5468
rect 19732 5408 19796 5412
rect 19812 5468 19876 5472
rect 19812 5412 19816 5468
rect 19816 5412 19872 5468
rect 19872 5412 19876 5468
rect 19812 5408 19876 5412
rect 19892 5468 19956 5472
rect 19892 5412 19896 5468
rect 19896 5412 19952 5468
rect 19952 5412 19956 5468
rect 19892 5408 19956 5412
rect 19972 5468 20036 5472
rect 19972 5412 19976 5468
rect 19976 5412 20032 5468
rect 20032 5412 20036 5468
rect 19972 5408 20036 5412
rect 27652 5468 27716 5472
rect 27652 5412 27656 5468
rect 27656 5412 27712 5468
rect 27712 5412 27716 5468
rect 27652 5408 27716 5412
rect 27732 5468 27796 5472
rect 27732 5412 27736 5468
rect 27736 5412 27792 5468
rect 27792 5412 27796 5468
rect 27732 5408 27796 5412
rect 27812 5468 27876 5472
rect 27812 5412 27816 5468
rect 27816 5412 27872 5468
rect 27872 5412 27876 5468
rect 27812 5408 27876 5412
rect 27892 5468 27956 5472
rect 27892 5412 27896 5468
rect 27896 5412 27952 5468
rect 27952 5412 27956 5468
rect 27892 5408 27956 5412
rect 27972 5468 28036 5472
rect 27972 5412 27976 5468
rect 27976 5412 28032 5468
rect 28032 5412 28036 5468
rect 27972 5408 28036 5412
rect 796 5204 860 5268
rect 796 4932 860 4996
rect 2912 4924 2976 4928
rect 2912 4868 2916 4924
rect 2916 4868 2972 4924
rect 2972 4868 2976 4924
rect 2912 4864 2976 4868
rect 2992 4924 3056 4928
rect 2992 4868 2996 4924
rect 2996 4868 3052 4924
rect 3052 4868 3056 4924
rect 2992 4864 3056 4868
rect 3072 4924 3136 4928
rect 3072 4868 3076 4924
rect 3076 4868 3132 4924
rect 3132 4868 3136 4924
rect 3072 4864 3136 4868
rect 3152 4924 3216 4928
rect 3152 4868 3156 4924
rect 3156 4868 3212 4924
rect 3212 4868 3216 4924
rect 3152 4864 3216 4868
rect 3232 4924 3296 4928
rect 3232 4868 3236 4924
rect 3236 4868 3292 4924
rect 3292 4868 3296 4924
rect 3232 4864 3296 4868
rect 10912 4924 10976 4928
rect 10912 4868 10916 4924
rect 10916 4868 10972 4924
rect 10972 4868 10976 4924
rect 10912 4864 10976 4868
rect 10992 4924 11056 4928
rect 10992 4868 10996 4924
rect 10996 4868 11052 4924
rect 11052 4868 11056 4924
rect 10992 4864 11056 4868
rect 11072 4924 11136 4928
rect 11072 4868 11076 4924
rect 11076 4868 11132 4924
rect 11132 4868 11136 4924
rect 11072 4864 11136 4868
rect 11152 4924 11216 4928
rect 11152 4868 11156 4924
rect 11156 4868 11212 4924
rect 11212 4868 11216 4924
rect 11152 4864 11216 4868
rect 11232 4924 11296 4928
rect 11232 4868 11236 4924
rect 11236 4868 11292 4924
rect 11292 4868 11296 4924
rect 11232 4864 11296 4868
rect 18912 4924 18976 4928
rect 18912 4868 18916 4924
rect 18916 4868 18972 4924
rect 18972 4868 18976 4924
rect 18912 4864 18976 4868
rect 18992 4924 19056 4928
rect 18992 4868 18996 4924
rect 18996 4868 19052 4924
rect 19052 4868 19056 4924
rect 18992 4864 19056 4868
rect 19072 4924 19136 4928
rect 19072 4868 19076 4924
rect 19076 4868 19132 4924
rect 19132 4868 19136 4924
rect 19072 4864 19136 4868
rect 19152 4924 19216 4928
rect 19152 4868 19156 4924
rect 19156 4868 19212 4924
rect 19212 4868 19216 4924
rect 19152 4864 19216 4868
rect 19232 4924 19296 4928
rect 19232 4868 19236 4924
rect 19236 4868 19292 4924
rect 19292 4868 19296 4924
rect 19232 4864 19296 4868
rect 26912 4924 26976 4928
rect 26912 4868 26916 4924
rect 26916 4868 26972 4924
rect 26972 4868 26976 4924
rect 26912 4864 26976 4868
rect 26992 4924 27056 4928
rect 26992 4868 26996 4924
rect 26996 4868 27052 4924
rect 27052 4868 27056 4924
rect 26992 4864 27056 4868
rect 27072 4924 27136 4928
rect 27072 4868 27076 4924
rect 27076 4868 27132 4924
rect 27132 4868 27136 4924
rect 27072 4864 27136 4868
rect 27152 4924 27216 4928
rect 27152 4868 27156 4924
rect 27156 4868 27212 4924
rect 27212 4868 27216 4924
rect 27152 4864 27216 4868
rect 27232 4924 27296 4928
rect 27232 4868 27236 4924
rect 27236 4868 27292 4924
rect 27292 4868 27296 4924
rect 27232 4864 27296 4868
rect 3652 4380 3716 4384
rect 3652 4324 3656 4380
rect 3656 4324 3712 4380
rect 3712 4324 3716 4380
rect 3652 4320 3716 4324
rect 3732 4380 3796 4384
rect 3732 4324 3736 4380
rect 3736 4324 3792 4380
rect 3792 4324 3796 4380
rect 3732 4320 3796 4324
rect 3812 4380 3876 4384
rect 3812 4324 3816 4380
rect 3816 4324 3872 4380
rect 3872 4324 3876 4380
rect 3812 4320 3876 4324
rect 3892 4380 3956 4384
rect 3892 4324 3896 4380
rect 3896 4324 3952 4380
rect 3952 4324 3956 4380
rect 3892 4320 3956 4324
rect 3972 4380 4036 4384
rect 3972 4324 3976 4380
rect 3976 4324 4032 4380
rect 4032 4324 4036 4380
rect 3972 4320 4036 4324
rect 11652 4380 11716 4384
rect 11652 4324 11656 4380
rect 11656 4324 11712 4380
rect 11712 4324 11716 4380
rect 11652 4320 11716 4324
rect 11732 4380 11796 4384
rect 11732 4324 11736 4380
rect 11736 4324 11792 4380
rect 11792 4324 11796 4380
rect 11732 4320 11796 4324
rect 11812 4380 11876 4384
rect 11812 4324 11816 4380
rect 11816 4324 11872 4380
rect 11872 4324 11876 4380
rect 11812 4320 11876 4324
rect 11892 4380 11956 4384
rect 11892 4324 11896 4380
rect 11896 4324 11952 4380
rect 11952 4324 11956 4380
rect 11892 4320 11956 4324
rect 11972 4380 12036 4384
rect 11972 4324 11976 4380
rect 11976 4324 12032 4380
rect 12032 4324 12036 4380
rect 11972 4320 12036 4324
rect 19652 4380 19716 4384
rect 19652 4324 19656 4380
rect 19656 4324 19712 4380
rect 19712 4324 19716 4380
rect 19652 4320 19716 4324
rect 19732 4380 19796 4384
rect 19732 4324 19736 4380
rect 19736 4324 19792 4380
rect 19792 4324 19796 4380
rect 19732 4320 19796 4324
rect 19812 4380 19876 4384
rect 19812 4324 19816 4380
rect 19816 4324 19872 4380
rect 19872 4324 19876 4380
rect 19812 4320 19876 4324
rect 19892 4380 19956 4384
rect 19892 4324 19896 4380
rect 19896 4324 19952 4380
rect 19952 4324 19956 4380
rect 19892 4320 19956 4324
rect 19972 4380 20036 4384
rect 19972 4324 19976 4380
rect 19976 4324 20032 4380
rect 20032 4324 20036 4380
rect 19972 4320 20036 4324
rect 27652 4380 27716 4384
rect 27652 4324 27656 4380
rect 27656 4324 27712 4380
rect 27712 4324 27716 4380
rect 27652 4320 27716 4324
rect 27732 4380 27796 4384
rect 27732 4324 27736 4380
rect 27736 4324 27792 4380
rect 27792 4324 27796 4380
rect 27732 4320 27796 4324
rect 27812 4380 27876 4384
rect 27812 4324 27816 4380
rect 27816 4324 27872 4380
rect 27872 4324 27876 4380
rect 27812 4320 27876 4324
rect 27892 4380 27956 4384
rect 27892 4324 27896 4380
rect 27896 4324 27952 4380
rect 27952 4324 27956 4380
rect 27892 4320 27956 4324
rect 27972 4380 28036 4384
rect 27972 4324 27976 4380
rect 27976 4324 28032 4380
rect 28032 4324 28036 4380
rect 27972 4320 28036 4324
rect 2912 3836 2976 3840
rect 2912 3780 2916 3836
rect 2916 3780 2972 3836
rect 2972 3780 2976 3836
rect 2912 3776 2976 3780
rect 2992 3836 3056 3840
rect 2992 3780 2996 3836
rect 2996 3780 3052 3836
rect 3052 3780 3056 3836
rect 2992 3776 3056 3780
rect 3072 3836 3136 3840
rect 3072 3780 3076 3836
rect 3076 3780 3132 3836
rect 3132 3780 3136 3836
rect 3072 3776 3136 3780
rect 3152 3836 3216 3840
rect 3152 3780 3156 3836
rect 3156 3780 3212 3836
rect 3212 3780 3216 3836
rect 3152 3776 3216 3780
rect 3232 3836 3296 3840
rect 3232 3780 3236 3836
rect 3236 3780 3292 3836
rect 3292 3780 3296 3836
rect 3232 3776 3296 3780
rect 10912 3836 10976 3840
rect 10912 3780 10916 3836
rect 10916 3780 10972 3836
rect 10972 3780 10976 3836
rect 10912 3776 10976 3780
rect 10992 3836 11056 3840
rect 10992 3780 10996 3836
rect 10996 3780 11052 3836
rect 11052 3780 11056 3836
rect 10992 3776 11056 3780
rect 11072 3836 11136 3840
rect 11072 3780 11076 3836
rect 11076 3780 11132 3836
rect 11132 3780 11136 3836
rect 11072 3776 11136 3780
rect 11152 3836 11216 3840
rect 11152 3780 11156 3836
rect 11156 3780 11212 3836
rect 11212 3780 11216 3836
rect 11152 3776 11216 3780
rect 11232 3836 11296 3840
rect 11232 3780 11236 3836
rect 11236 3780 11292 3836
rect 11292 3780 11296 3836
rect 11232 3776 11296 3780
rect 18912 3836 18976 3840
rect 18912 3780 18916 3836
rect 18916 3780 18972 3836
rect 18972 3780 18976 3836
rect 18912 3776 18976 3780
rect 18992 3836 19056 3840
rect 18992 3780 18996 3836
rect 18996 3780 19052 3836
rect 19052 3780 19056 3836
rect 18992 3776 19056 3780
rect 19072 3836 19136 3840
rect 19072 3780 19076 3836
rect 19076 3780 19132 3836
rect 19132 3780 19136 3836
rect 19072 3776 19136 3780
rect 19152 3836 19216 3840
rect 19152 3780 19156 3836
rect 19156 3780 19212 3836
rect 19212 3780 19216 3836
rect 19152 3776 19216 3780
rect 19232 3836 19296 3840
rect 19232 3780 19236 3836
rect 19236 3780 19292 3836
rect 19292 3780 19296 3836
rect 19232 3776 19296 3780
rect 26912 3836 26976 3840
rect 26912 3780 26916 3836
rect 26916 3780 26972 3836
rect 26972 3780 26976 3836
rect 26912 3776 26976 3780
rect 26992 3836 27056 3840
rect 26992 3780 26996 3836
rect 26996 3780 27052 3836
rect 27052 3780 27056 3836
rect 26992 3776 27056 3780
rect 27072 3836 27136 3840
rect 27072 3780 27076 3836
rect 27076 3780 27132 3836
rect 27132 3780 27136 3836
rect 27072 3776 27136 3780
rect 27152 3836 27216 3840
rect 27152 3780 27156 3836
rect 27156 3780 27212 3836
rect 27212 3780 27216 3836
rect 27152 3776 27216 3780
rect 27232 3836 27296 3840
rect 27232 3780 27236 3836
rect 27236 3780 27292 3836
rect 27292 3780 27296 3836
rect 27232 3776 27296 3780
rect 3652 3292 3716 3296
rect 3652 3236 3656 3292
rect 3656 3236 3712 3292
rect 3712 3236 3716 3292
rect 3652 3232 3716 3236
rect 3732 3292 3796 3296
rect 3732 3236 3736 3292
rect 3736 3236 3792 3292
rect 3792 3236 3796 3292
rect 3732 3232 3796 3236
rect 3812 3292 3876 3296
rect 3812 3236 3816 3292
rect 3816 3236 3872 3292
rect 3872 3236 3876 3292
rect 3812 3232 3876 3236
rect 3892 3292 3956 3296
rect 3892 3236 3896 3292
rect 3896 3236 3952 3292
rect 3952 3236 3956 3292
rect 3892 3232 3956 3236
rect 3972 3292 4036 3296
rect 3972 3236 3976 3292
rect 3976 3236 4032 3292
rect 4032 3236 4036 3292
rect 3972 3232 4036 3236
rect 11652 3292 11716 3296
rect 11652 3236 11656 3292
rect 11656 3236 11712 3292
rect 11712 3236 11716 3292
rect 11652 3232 11716 3236
rect 11732 3292 11796 3296
rect 11732 3236 11736 3292
rect 11736 3236 11792 3292
rect 11792 3236 11796 3292
rect 11732 3232 11796 3236
rect 11812 3292 11876 3296
rect 11812 3236 11816 3292
rect 11816 3236 11872 3292
rect 11872 3236 11876 3292
rect 11812 3232 11876 3236
rect 11892 3292 11956 3296
rect 11892 3236 11896 3292
rect 11896 3236 11952 3292
rect 11952 3236 11956 3292
rect 11892 3232 11956 3236
rect 11972 3292 12036 3296
rect 11972 3236 11976 3292
rect 11976 3236 12032 3292
rect 12032 3236 12036 3292
rect 11972 3232 12036 3236
rect 19652 3292 19716 3296
rect 19652 3236 19656 3292
rect 19656 3236 19712 3292
rect 19712 3236 19716 3292
rect 19652 3232 19716 3236
rect 19732 3292 19796 3296
rect 19732 3236 19736 3292
rect 19736 3236 19792 3292
rect 19792 3236 19796 3292
rect 19732 3232 19796 3236
rect 19812 3292 19876 3296
rect 19812 3236 19816 3292
rect 19816 3236 19872 3292
rect 19872 3236 19876 3292
rect 19812 3232 19876 3236
rect 19892 3292 19956 3296
rect 19892 3236 19896 3292
rect 19896 3236 19952 3292
rect 19952 3236 19956 3292
rect 19892 3232 19956 3236
rect 19972 3292 20036 3296
rect 19972 3236 19976 3292
rect 19976 3236 20032 3292
rect 20032 3236 20036 3292
rect 19972 3232 20036 3236
rect 27652 3292 27716 3296
rect 27652 3236 27656 3292
rect 27656 3236 27712 3292
rect 27712 3236 27716 3292
rect 27652 3232 27716 3236
rect 27732 3292 27796 3296
rect 27732 3236 27736 3292
rect 27736 3236 27792 3292
rect 27792 3236 27796 3292
rect 27732 3232 27796 3236
rect 27812 3292 27876 3296
rect 27812 3236 27816 3292
rect 27816 3236 27872 3292
rect 27872 3236 27876 3292
rect 27812 3232 27876 3236
rect 27892 3292 27956 3296
rect 27892 3236 27896 3292
rect 27896 3236 27952 3292
rect 27952 3236 27956 3292
rect 27892 3232 27956 3236
rect 27972 3292 28036 3296
rect 27972 3236 27976 3292
rect 27976 3236 28032 3292
rect 28032 3236 28036 3292
rect 27972 3232 28036 3236
rect 2912 2748 2976 2752
rect 2912 2692 2916 2748
rect 2916 2692 2972 2748
rect 2972 2692 2976 2748
rect 2912 2688 2976 2692
rect 2992 2748 3056 2752
rect 2992 2692 2996 2748
rect 2996 2692 3052 2748
rect 3052 2692 3056 2748
rect 2992 2688 3056 2692
rect 3072 2748 3136 2752
rect 3072 2692 3076 2748
rect 3076 2692 3132 2748
rect 3132 2692 3136 2748
rect 3072 2688 3136 2692
rect 3152 2748 3216 2752
rect 3152 2692 3156 2748
rect 3156 2692 3212 2748
rect 3212 2692 3216 2748
rect 3152 2688 3216 2692
rect 3232 2748 3296 2752
rect 3232 2692 3236 2748
rect 3236 2692 3292 2748
rect 3292 2692 3296 2748
rect 3232 2688 3296 2692
rect 10912 2748 10976 2752
rect 10912 2692 10916 2748
rect 10916 2692 10972 2748
rect 10972 2692 10976 2748
rect 10912 2688 10976 2692
rect 10992 2748 11056 2752
rect 10992 2692 10996 2748
rect 10996 2692 11052 2748
rect 11052 2692 11056 2748
rect 10992 2688 11056 2692
rect 11072 2748 11136 2752
rect 11072 2692 11076 2748
rect 11076 2692 11132 2748
rect 11132 2692 11136 2748
rect 11072 2688 11136 2692
rect 11152 2748 11216 2752
rect 11152 2692 11156 2748
rect 11156 2692 11212 2748
rect 11212 2692 11216 2748
rect 11152 2688 11216 2692
rect 11232 2748 11296 2752
rect 11232 2692 11236 2748
rect 11236 2692 11292 2748
rect 11292 2692 11296 2748
rect 11232 2688 11296 2692
rect 18912 2748 18976 2752
rect 18912 2692 18916 2748
rect 18916 2692 18972 2748
rect 18972 2692 18976 2748
rect 18912 2688 18976 2692
rect 18992 2748 19056 2752
rect 18992 2692 18996 2748
rect 18996 2692 19052 2748
rect 19052 2692 19056 2748
rect 18992 2688 19056 2692
rect 19072 2748 19136 2752
rect 19072 2692 19076 2748
rect 19076 2692 19132 2748
rect 19132 2692 19136 2748
rect 19072 2688 19136 2692
rect 19152 2748 19216 2752
rect 19152 2692 19156 2748
rect 19156 2692 19212 2748
rect 19212 2692 19216 2748
rect 19152 2688 19216 2692
rect 19232 2748 19296 2752
rect 19232 2692 19236 2748
rect 19236 2692 19292 2748
rect 19292 2692 19296 2748
rect 19232 2688 19296 2692
rect 26912 2748 26976 2752
rect 26912 2692 26916 2748
rect 26916 2692 26972 2748
rect 26972 2692 26976 2748
rect 26912 2688 26976 2692
rect 26992 2748 27056 2752
rect 26992 2692 26996 2748
rect 26996 2692 27052 2748
rect 27052 2692 27056 2748
rect 26992 2688 27056 2692
rect 27072 2748 27136 2752
rect 27072 2692 27076 2748
rect 27076 2692 27132 2748
rect 27132 2692 27136 2748
rect 27072 2688 27136 2692
rect 27152 2748 27216 2752
rect 27152 2692 27156 2748
rect 27156 2692 27212 2748
rect 27212 2692 27216 2748
rect 27152 2688 27216 2692
rect 27232 2748 27296 2752
rect 27232 2692 27236 2748
rect 27236 2692 27292 2748
rect 27292 2692 27296 2748
rect 27232 2688 27296 2692
rect 3652 2204 3716 2208
rect 3652 2148 3656 2204
rect 3656 2148 3712 2204
rect 3712 2148 3716 2204
rect 3652 2144 3716 2148
rect 3732 2204 3796 2208
rect 3732 2148 3736 2204
rect 3736 2148 3792 2204
rect 3792 2148 3796 2204
rect 3732 2144 3796 2148
rect 3812 2204 3876 2208
rect 3812 2148 3816 2204
rect 3816 2148 3872 2204
rect 3872 2148 3876 2204
rect 3812 2144 3876 2148
rect 3892 2204 3956 2208
rect 3892 2148 3896 2204
rect 3896 2148 3952 2204
rect 3952 2148 3956 2204
rect 3892 2144 3956 2148
rect 3972 2204 4036 2208
rect 3972 2148 3976 2204
rect 3976 2148 4032 2204
rect 4032 2148 4036 2204
rect 3972 2144 4036 2148
rect 11652 2204 11716 2208
rect 11652 2148 11656 2204
rect 11656 2148 11712 2204
rect 11712 2148 11716 2204
rect 11652 2144 11716 2148
rect 11732 2204 11796 2208
rect 11732 2148 11736 2204
rect 11736 2148 11792 2204
rect 11792 2148 11796 2204
rect 11732 2144 11796 2148
rect 11812 2204 11876 2208
rect 11812 2148 11816 2204
rect 11816 2148 11872 2204
rect 11872 2148 11876 2204
rect 11812 2144 11876 2148
rect 11892 2204 11956 2208
rect 11892 2148 11896 2204
rect 11896 2148 11952 2204
rect 11952 2148 11956 2204
rect 11892 2144 11956 2148
rect 11972 2204 12036 2208
rect 11972 2148 11976 2204
rect 11976 2148 12032 2204
rect 12032 2148 12036 2204
rect 11972 2144 12036 2148
rect 19652 2204 19716 2208
rect 19652 2148 19656 2204
rect 19656 2148 19712 2204
rect 19712 2148 19716 2204
rect 19652 2144 19716 2148
rect 19732 2204 19796 2208
rect 19732 2148 19736 2204
rect 19736 2148 19792 2204
rect 19792 2148 19796 2204
rect 19732 2144 19796 2148
rect 19812 2204 19876 2208
rect 19812 2148 19816 2204
rect 19816 2148 19872 2204
rect 19872 2148 19876 2204
rect 19812 2144 19876 2148
rect 19892 2204 19956 2208
rect 19892 2148 19896 2204
rect 19896 2148 19952 2204
rect 19952 2148 19956 2204
rect 19892 2144 19956 2148
rect 19972 2204 20036 2208
rect 19972 2148 19976 2204
rect 19976 2148 20032 2204
rect 20032 2148 20036 2204
rect 19972 2144 20036 2148
rect 27652 2204 27716 2208
rect 27652 2148 27656 2204
rect 27656 2148 27712 2204
rect 27712 2148 27716 2204
rect 27652 2144 27716 2148
rect 27732 2204 27796 2208
rect 27732 2148 27736 2204
rect 27736 2148 27792 2204
rect 27792 2148 27796 2204
rect 27732 2144 27796 2148
rect 27812 2204 27876 2208
rect 27812 2148 27816 2204
rect 27816 2148 27872 2204
rect 27872 2148 27876 2204
rect 27812 2144 27876 2148
rect 27892 2204 27956 2208
rect 27892 2148 27896 2204
rect 27896 2148 27952 2204
rect 27952 2148 27956 2204
rect 27892 2144 27956 2148
rect 27972 2204 28036 2208
rect 27972 2148 27976 2204
rect 27976 2148 28032 2204
rect 28032 2148 28036 2204
rect 27972 2144 28036 2148
<< metal4 >>
rect 2904 27776 3304 27792
rect 2904 27712 2912 27776
rect 2976 27712 2992 27776
rect 3056 27712 3072 27776
rect 3136 27712 3152 27776
rect 3216 27712 3232 27776
rect 3296 27712 3304 27776
rect 2904 26688 3304 27712
rect 2904 26624 2912 26688
rect 2976 26624 2992 26688
rect 3056 26624 3072 26688
rect 3136 26624 3152 26688
rect 3216 26624 3232 26688
rect 3296 26624 3304 26688
rect 2904 25600 3304 26624
rect 2904 25536 2912 25600
rect 2976 25536 2992 25600
rect 3056 25536 3072 25600
rect 3136 25536 3152 25600
rect 3216 25536 3232 25600
rect 3296 25536 3304 25600
rect 2904 24512 3304 25536
rect 2904 24448 2912 24512
rect 2976 24448 2992 24512
rect 3056 24448 3072 24512
rect 3136 24448 3152 24512
rect 3216 24448 3232 24512
rect 3296 24448 3304 24512
rect 2904 23424 3304 24448
rect 2904 23360 2912 23424
rect 2976 23360 2992 23424
rect 3056 23360 3072 23424
rect 3136 23360 3152 23424
rect 3216 23360 3232 23424
rect 3296 23360 3304 23424
rect 2904 22336 3304 23360
rect 2904 22272 2912 22336
rect 2976 22272 2992 22336
rect 3056 22272 3072 22336
rect 3136 22272 3152 22336
rect 3216 22272 3232 22336
rect 3296 22272 3304 22336
rect 2904 21248 3304 22272
rect 2904 21184 2912 21248
rect 2976 21184 2992 21248
rect 3056 21184 3072 21248
rect 3136 21184 3152 21248
rect 3216 21184 3232 21248
rect 3296 21184 3304 21248
rect 2904 20160 3304 21184
rect 2904 20096 2912 20160
rect 2976 20096 2992 20160
rect 3056 20096 3072 20160
rect 3136 20096 3152 20160
rect 3216 20096 3232 20160
rect 3296 20096 3304 20160
rect 2904 19072 3304 20096
rect 2904 19008 2912 19072
rect 2976 19008 2992 19072
rect 3056 19008 3072 19072
rect 3136 19008 3152 19072
rect 3216 19008 3232 19072
rect 3296 19008 3304 19072
rect 2904 17984 3304 19008
rect 2904 17920 2912 17984
rect 2976 17920 2992 17984
rect 3056 17920 3072 17984
rect 3136 17920 3152 17984
rect 3216 17920 3232 17984
rect 3296 17920 3304 17984
rect 2904 16896 3304 17920
rect 2904 16832 2912 16896
rect 2976 16832 2992 16896
rect 3056 16832 3072 16896
rect 3136 16832 3152 16896
rect 3216 16832 3232 16896
rect 3296 16832 3304 16896
rect 2904 15808 3304 16832
rect 2904 15744 2912 15808
rect 2976 15744 2992 15808
rect 3056 15744 3072 15808
rect 3136 15744 3152 15808
rect 3216 15744 3232 15808
rect 3296 15744 3304 15808
rect 2904 14720 3304 15744
rect 2904 14656 2912 14720
rect 2976 14656 2992 14720
rect 3056 14656 3072 14720
rect 3136 14656 3152 14720
rect 3216 14656 3232 14720
rect 3296 14656 3304 14720
rect 2904 13632 3304 14656
rect 2904 13568 2912 13632
rect 2976 13568 2992 13632
rect 3056 13568 3072 13632
rect 3136 13568 3152 13632
rect 3216 13568 3232 13632
rect 3296 13568 3304 13632
rect 2904 12544 3304 13568
rect 2904 12480 2912 12544
rect 2976 12480 2992 12544
rect 3056 12480 3072 12544
rect 3136 12480 3152 12544
rect 3216 12480 3232 12544
rect 3296 12480 3304 12544
rect 2904 11456 3304 12480
rect 2904 11392 2912 11456
rect 2976 11392 2992 11456
rect 3056 11392 3072 11456
rect 3136 11392 3152 11456
rect 3216 11392 3232 11456
rect 3296 11392 3304 11456
rect 2904 10368 3304 11392
rect 2904 10304 2912 10368
rect 2976 10304 2992 10368
rect 3056 10304 3072 10368
rect 3136 10304 3152 10368
rect 3216 10304 3232 10368
rect 3296 10304 3304 10368
rect 2904 9280 3304 10304
rect 2904 9216 2912 9280
rect 2976 9216 2992 9280
rect 3056 9216 3072 9280
rect 3136 9216 3152 9280
rect 3216 9216 3232 9280
rect 3296 9216 3304 9280
rect 2904 8192 3304 9216
rect 2904 8128 2912 8192
rect 2976 8128 2992 8192
rect 3056 8128 3072 8192
rect 3136 8128 3152 8192
rect 3216 8128 3232 8192
rect 3296 8128 3304 8192
rect 2904 7104 3304 8128
rect 2904 7040 2912 7104
rect 2976 7040 2992 7104
rect 3056 7040 3072 7104
rect 3136 7040 3152 7104
rect 3216 7040 3232 7104
rect 3296 7040 3304 7104
rect 2904 6016 3304 7040
rect 2904 5952 2912 6016
rect 2976 5952 2992 6016
rect 3056 5952 3072 6016
rect 3136 5952 3152 6016
rect 3216 5952 3232 6016
rect 3296 5952 3304 6016
rect 795 5268 861 5269
rect 795 5204 796 5268
rect 860 5204 861 5268
rect 795 5203 861 5204
rect 798 4997 858 5203
rect 795 4996 861 4997
rect 795 4932 796 4996
rect 860 4932 861 4996
rect 795 4931 861 4932
rect 2904 4928 3304 5952
rect 2904 4864 2912 4928
rect 2976 4864 2992 4928
rect 3056 4864 3072 4928
rect 3136 4864 3152 4928
rect 3216 4864 3232 4928
rect 3296 4864 3304 4928
rect 2904 3840 3304 4864
rect 2904 3776 2912 3840
rect 2976 3776 2992 3840
rect 3056 3776 3072 3840
rect 3136 3776 3152 3840
rect 3216 3776 3232 3840
rect 3296 3776 3304 3840
rect 2904 2752 3304 3776
rect 2904 2688 2912 2752
rect 2976 2688 2992 2752
rect 3056 2688 3072 2752
rect 3136 2688 3152 2752
rect 3216 2688 3232 2752
rect 3296 2688 3304 2752
rect 2904 2128 3304 2688
rect 3644 27232 4044 27792
rect 3644 27168 3652 27232
rect 3716 27168 3732 27232
rect 3796 27168 3812 27232
rect 3876 27168 3892 27232
rect 3956 27168 3972 27232
rect 4036 27168 4044 27232
rect 3644 26144 4044 27168
rect 3644 26080 3652 26144
rect 3716 26080 3732 26144
rect 3796 26080 3812 26144
rect 3876 26080 3892 26144
rect 3956 26080 3972 26144
rect 4036 26080 4044 26144
rect 3644 25056 4044 26080
rect 3644 24992 3652 25056
rect 3716 24992 3732 25056
rect 3796 24992 3812 25056
rect 3876 24992 3892 25056
rect 3956 24992 3972 25056
rect 4036 24992 4044 25056
rect 3644 23968 4044 24992
rect 3644 23904 3652 23968
rect 3716 23904 3732 23968
rect 3796 23904 3812 23968
rect 3876 23904 3892 23968
rect 3956 23904 3972 23968
rect 4036 23904 4044 23968
rect 3644 22880 4044 23904
rect 3644 22816 3652 22880
rect 3716 22816 3732 22880
rect 3796 22816 3812 22880
rect 3876 22816 3892 22880
rect 3956 22816 3972 22880
rect 4036 22816 4044 22880
rect 3644 21792 4044 22816
rect 3644 21728 3652 21792
rect 3716 21728 3732 21792
rect 3796 21728 3812 21792
rect 3876 21728 3892 21792
rect 3956 21728 3972 21792
rect 4036 21728 4044 21792
rect 3644 20704 4044 21728
rect 3644 20640 3652 20704
rect 3716 20640 3732 20704
rect 3796 20640 3812 20704
rect 3876 20640 3892 20704
rect 3956 20640 3972 20704
rect 4036 20640 4044 20704
rect 3644 19616 4044 20640
rect 3644 19552 3652 19616
rect 3716 19552 3732 19616
rect 3796 19552 3812 19616
rect 3876 19552 3892 19616
rect 3956 19552 3972 19616
rect 4036 19552 4044 19616
rect 3644 18528 4044 19552
rect 3644 18464 3652 18528
rect 3716 18464 3732 18528
rect 3796 18464 3812 18528
rect 3876 18464 3892 18528
rect 3956 18464 3972 18528
rect 4036 18464 4044 18528
rect 3644 17440 4044 18464
rect 3644 17376 3652 17440
rect 3716 17376 3732 17440
rect 3796 17376 3812 17440
rect 3876 17376 3892 17440
rect 3956 17376 3972 17440
rect 4036 17376 4044 17440
rect 3644 16352 4044 17376
rect 3644 16288 3652 16352
rect 3716 16288 3732 16352
rect 3796 16288 3812 16352
rect 3876 16288 3892 16352
rect 3956 16288 3972 16352
rect 4036 16288 4044 16352
rect 3644 15264 4044 16288
rect 3644 15200 3652 15264
rect 3716 15200 3732 15264
rect 3796 15200 3812 15264
rect 3876 15200 3892 15264
rect 3956 15200 3972 15264
rect 4036 15200 4044 15264
rect 3644 14176 4044 15200
rect 3644 14112 3652 14176
rect 3716 14112 3732 14176
rect 3796 14112 3812 14176
rect 3876 14112 3892 14176
rect 3956 14112 3972 14176
rect 4036 14112 4044 14176
rect 3644 13088 4044 14112
rect 3644 13024 3652 13088
rect 3716 13024 3732 13088
rect 3796 13024 3812 13088
rect 3876 13024 3892 13088
rect 3956 13024 3972 13088
rect 4036 13024 4044 13088
rect 3644 12000 4044 13024
rect 3644 11936 3652 12000
rect 3716 11936 3732 12000
rect 3796 11936 3812 12000
rect 3876 11936 3892 12000
rect 3956 11936 3972 12000
rect 4036 11936 4044 12000
rect 3644 10912 4044 11936
rect 3644 10848 3652 10912
rect 3716 10848 3732 10912
rect 3796 10848 3812 10912
rect 3876 10848 3892 10912
rect 3956 10848 3972 10912
rect 4036 10848 4044 10912
rect 3644 9824 4044 10848
rect 3644 9760 3652 9824
rect 3716 9760 3732 9824
rect 3796 9760 3812 9824
rect 3876 9760 3892 9824
rect 3956 9760 3972 9824
rect 4036 9760 4044 9824
rect 3644 8736 4044 9760
rect 3644 8672 3652 8736
rect 3716 8672 3732 8736
rect 3796 8672 3812 8736
rect 3876 8672 3892 8736
rect 3956 8672 3972 8736
rect 4036 8672 4044 8736
rect 3644 7648 4044 8672
rect 3644 7584 3652 7648
rect 3716 7584 3732 7648
rect 3796 7584 3812 7648
rect 3876 7584 3892 7648
rect 3956 7584 3972 7648
rect 4036 7584 4044 7648
rect 3644 6560 4044 7584
rect 3644 6496 3652 6560
rect 3716 6496 3732 6560
rect 3796 6496 3812 6560
rect 3876 6496 3892 6560
rect 3956 6496 3972 6560
rect 4036 6496 4044 6560
rect 3644 5472 4044 6496
rect 3644 5408 3652 5472
rect 3716 5408 3732 5472
rect 3796 5408 3812 5472
rect 3876 5408 3892 5472
rect 3956 5408 3972 5472
rect 4036 5408 4044 5472
rect 3644 4384 4044 5408
rect 3644 4320 3652 4384
rect 3716 4320 3732 4384
rect 3796 4320 3812 4384
rect 3876 4320 3892 4384
rect 3956 4320 3972 4384
rect 4036 4320 4044 4384
rect 3644 3296 4044 4320
rect 3644 3232 3652 3296
rect 3716 3232 3732 3296
rect 3796 3232 3812 3296
rect 3876 3232 3892 3296
rect 3956 3232 3972 3296
rect 4036 3232 4044 3296
rect 3644 2208 4044 3232
rect 3644 2144 3652 2208
rect 3716 2144 3732 2208
rect 3796 2144 3812 2208
rect 3876 2144 3892 2208
rect 3956 2144 3972 2208
rect 4036 2144 4044 2208
rect 3644 2128 4044 2144
rect 10904 27776 11304 27792
rect 10904 27712 10912 27776
rect 10976 27712 10992 27776
rect 11056 27712 11072 27776
rect 11136 27712 11152 27776
rect 11216 27712 11232 27776
rect 11296 27712 11304 27776
rect 10904 26688 11304 27712
rect 10904 26624 10912 26688
rect 10976 26624 10992 26688
rect 11056 26624 11072 26688
rect 11136 26624 11152 26688
rect 11216 26624 11232 26688
rect 11296 26624 11304 26688
rect 10904 25600 11304 26624
rect 10904 25536 10912 25600
rect 10976 25536 10992 25600
rect 11056 25536 11072 25600
rect 11136 25536 11152 25600
rect 11216 25536 11232 25600
rect 11296 25536 11304 25600
rect 10904 24512 11304 25536
rect 10904 24448 10912 24512
rect 10976 24448 10992 24512
rect 11056 24448 11072 24512
rect 11136 24448 11152 24512
rect 11216 24448 11232 24512
rect 11296 24448 11304 24512
rect 10904 23424 11304 24448
rect 10904 23360 10912 23424
rect 10976 23360 10992 23424
rect 11056 23360 11072 23424
rect 11136 23360 11152 23424
rect 11216 23360 11232 23424
rect 11296 23360 11304 23424
rect 10904 22336 11304 23360
rect 10904 22272 10912 22336
rect 10976 22272 10992 22336
rect 11056 22272 11072 22336
rect 11136 22272 11152 22336
rect 11216 22272 11232 22336
rect 11296 22272 11304 22336
rect 10904 21248 11304 22272
rect 10904 21184 10912 21248
rect 10976 21184 10992 21248
rect 11056 21184 11072 21248
rect 11136 21184 11152 21248
rect 11216 21184 11232 21248
rect 11296 21184 11304 21248
rect 10904 20160 11304 21184
rect 10904 20096 10912 20160
rect 10976 20096 10992 20160
rect 11056 20096 11072 20160
rect 11136 20096 11152 20160
rect 11216 20096 11232 20160
rect 11296 20096 11304 20160
rect 10904 19072 11304 20096
rect 10904 19008 10912 19072
rect 10976 19008 10992 19072
rect 11056 19008 11072 19072
rect 11136 19008 11152 19072
rect 11216 19008 11232 19072
rect 11296 19008 11304 19072
rect 10904 17984 11304 19008
rect 10904 17920 10912 17984
rect 10976 17920 10992 17984
rect 11056 17920 11072 17984
rect 11136 17920 11152 17984
rect 11216 17920 11232 17984
rect 11296 17920 11304 17984
rect 10904 16896 11304 17920
rect 10904 16832 10912 16896
rect 10976 16832 10992 16896
rect 11056 16832 11072 16896
rect 11136 16832 11152 16896
rect 11216 16832 11232 16896
rect 11296 16832 11304 16896
rect 10904 15808 11304 16832
rect 10904 15744 10912 15808
rect 10976 15744 10992 15808
rect 11056 15744 11072 15808
rect 11136 15744 11152 15808
rect 11216 15744 11232 15808
rect 11296 15744 11304 15808
rect 10904 14720 11304 15744
rect 11644 27232 12044 27792
rect 11644 27168 11652 27232
rect 11716 27168 11732 27232
rect 11796 27168 11812 27232
rect 11876 27168 11892 27232
rect 11956 27168 11972 27232
rect 12036 27168 12044 27232
rect 11644 26144 12044 27168
rect 11644 26080 11652 26144
rect 11716 26080 11732 26144
rect 11796 26080 11812 26144
rect 11876 26080 11892 26144
rect 11956 26080 11972 26144
rect 12036 26080 12044 26144
rect 11644 25056 12044 26080
rect 11644 24992 11652 25056
rect 11716 24992 11732 25056
rect 11796 24992 11812 25056
rect 11876 24992 11892 25056
rect 11956 24992 11972 25056
rect 12036 24992 12044 25056
rect 11644 23968 12044 24992
rect 11644 23904 11652 23968
rect 11716 23904 11732 23968
rect 11796 23904 11812 23968
rect 11876 23904 11892 23968
rect 11956 23904 11972 23968
rect 12036 23904 12044 23968
rect 11644 22880 12044 23904
rect 11644 22816 11652 22880
rect 11716 22816 11732 22880
rect 11796 22816 11812 22880
rect 11876 22816 11892 22880
rect 11956 22816 11972 22880
rect 12036 22816 12044 22880
rect 11644 21792 12044 22816
rect 11644 21728 11652 21792
rect 11716 21728 11732 21792
rect 11796 21728 11812 21792
rect 11876 21728 11892 21792
rect 11956 21728 11972 21792
rect 12036 21728 12044 21792
rect 11644 20704 12044 21728
rect 11644 20640 11652 20704
rect 11716 20640 11732 20704
rect 11796 20640 11812 20704
rect 11876 20640 11892 20704
rect 11956 20640 11972 20704
rect 12036 20640 12044 20704
rect 11644 19616 12044 20640
rect 11644 19552 11652 19616
rect 11716 19552 11732 19616
rect 11796 19552 11812 19616
rect 11876 19552 11892 19616
rect 11956 19552 11972 19616
rect 12036 19552 12044 19616
rect 11644 18528 12044 19552
rect 11644 18464 11652 18528
rect 11716 18464 11732 18528
rect 11796 18464 11812 18528
rect 11876 18464 11892 18528
rect 11956 18464 11972 18528
rect 12036 18464 12044 18528
rect 11644 17440 12044 18464
rect 11644 17376 11652 17440
rect 11716 17376 11732 17440
rect 11796 17376 11812 17440
rect 11876 17376 11892 17440
rect 11956 17376 11972 17440
rect 12036 17376 12044 17440
rect 11644 16352 12044 17376
rect 11644 16288 11652 16352
rect 11716 16288 11732 16352
rect 11796 16288 11812 16352
rect 11876 16288 11892 16352
rect 11956 16288 11972 16352
rect 12036 16288 12044 16352
rect 11467 15468 11533 15469
rect 11467 15404 11468 15468
rect 11532 15404 11533 15468
rect 11467 15403 11533 15404
rect 10904 14656 10912 14720
rect 10976 14656 10992 14720
rect 11056 14656 11072 14720
rect 11136 14656 11152 14720
rect 11216 14656 11232 14720
rect 11296 14656 11304 14720
rect 10904 13632 11304 14656
rect 10904 13568 10912 13632
rect 10976 13568 10992 13632
rect 11056 13568 11072 13632
rect 11136 13568 11152 13632
rect 11216 13568 11232 13632
rect 11296 13568 11304 13632
rect 10904 12544 11304 13568
rect 10904 12480 10912 12544
rect 10976 12480 10992 12544
rect 11056 12480 11072 12544
rect 11136 12480 11152 12544
rect 11216 12480 11232 12544
rect 11296 12480 11304 12544
rect 10904 11456 11304 12480
rect 10904 11392 10912 11456
rect 10976 11392 10992 11456
rect 11056 11392 11072 11456
rect 11136 11392 11152 11456
rect 11216 11392 11232 11456
rect 11296 11392 11304 11456
rect 10904 10368 11304 11392
rect 11470 10437 11530 15403
rect 11644 15264 12044 16288
rect 11644 15200 11652 15264
rect 11716 15200 11732 15264
rect 11796 15200 11812 15264
rect 11876 15200 11892 15264
rect 11956 15200 11972 15264
rect 12036 15200 12044 15264
rect 11644 14176 12044 15200
rect 11644 14112 11652 14176
rect 11716 14112 11732 14176
rect 11796 14112 11812 14176
rect 11876 14112 11892 14176
rect 11956 14112 11972 14176
rect 12036 14112 12044 14176
rect 11644 13088 12044 14112
rect 11644 13024 11652 13088
rect 11716 13024 11732 13088
rect 11796 13024 11812 13088
rect 11876 13024 11892 13088
rect 11956 13024 11972 13088
rect 12036 13024 12044 13088
rect 11644 12000 12044 13024
rect 11644 11936 11652 12000
rect 11716 11936 11732 12000
rect 11796 11936 11812 12000
rect 11876 11936 11892 12000
rect 11956 11936 11972 12000
rect 12036 11936 12044 12000
rect 11644 10912 12044 11936
rect 11644 10848 11652 10912
rect 11716 10848 11732 10912
rect 11796 10848 11812 10912
rect 11876 10848 11892 10912
rect 11956 10848 11972 10912
rect 12036 10848 12044 10912
rect 11467 10436 11533 10437
rect 11467 10372 11468 10436
rect 11532 10372 11533 10436
rect 11467 10371 11533 10372
rect 10904 10304 10912 10368
rect 10976 10304 10992 10368
rect 11056 10304 11072 10368
rect 11136 10304 11152 10368
rect 11216 10304 11232 10368
rect 11296 10304 11304 10368
rect 10904 9280 11304 10304
rect 10904 9216 10912 9280
rect 10976 9216 10992 9280
rect 11056 9216 11072 9280
rect 11136 9216 11152 9280
rect 11216 9216 11232 9280
rect 11296 9216 11304 9280
rect 10904 8192 11304 9216
rect 10904 8128 10912 8192
rect 10976 8128 10992 8192
rect 11056 8128 11072 8192
rect 11136 8128 11152 8192
rect 11216 8128 11232 8192
rect 11296 8128 11304 8192
rect 10904 7104 11304 8128
rect 10904 7040 10912 7104
rect 10976 7040 10992 7104
rect 11056 7040 11072 7104
rect 11136 7040 11152 7104
rect 11216 7040 11232 7104
rect 11296 7040 11304 7104
rect 10904 6016 11304 7040
rect 10904 5952 10912 6016
rect 10976 5952 10992 6016
rect 11056 5952 11072 6016
rect 11136 5952 11152 6016
rect 11216 5952 11232 6016
rect 11296 5952 11304 6016
rect 10904 4928 11304 5952
rect 10904 4864 10912 4928
rect 10976 4864 10992 4928
rect 11056 4864 11072 4928
rect 11136 4864 11152 4928
rect 11216 4864 11232 4928
rect 11296 4864 11304 4928
rect 10904 3840 11304 4864
rect 10904 3776 10912 3840
rect 10976 3776 10992 3840
rect 11056 3776 11072 3840
rect 11136 3776 11152 3840
rect 11216 3776 11232 3840
rect 11296 3776 11304 3840
rect 10904 2752 11304 3776
rect 10904 2688 10912 2752
rect 10976 2688 10992 2752
rect 11056 2688 11072 2752
rect 11136 2688 11152 2752
rect 11216 2688 11232 2752
rect 11296 2688 11304 2752
rect 10904 2128 11304 2688
rect 11644 9824 12044 10848
rect 11644 9760 11652 9824
rect 11716 9760 11732 9824
rect 11796 9760 11812 9824
rect 11876 9760 11892 9824
rect 11956 9760 11972 9824
rect 12036 9760 12044 9824
rect 11644 8736 12044 9760
rect 11644 8672 11652 8736
rect 11716 8672 11732 8736
rect 11796 8672 11812 8736
rect 11876 8672 11892 8736
rect 11956 8672 11972 8736
rect 12036 8672 12044 8736
rect 11644 7648 12044 8672
rect 11644 7584 11652 7648
rect 11716 7584 11732 7648
rect 11796 7584 11812 7648
rect 11876 7584 11892 7648
rect 11956 7584 11972 7648
rect 12036 7584 12044 7648
rect 11644 6560 12044 7584
rect 11644 6496 11652 6560
rect 11716 6496 11732 6560
rect 11796 6496 11812 6560
rect 11876 6496 11892 6560
rect 11956 6496 11972 6560
rect 12036 6496 12044 6560
rect 11644 5472 12044 6496
rect 11644 5408 11652 5472
rect 11716 5408 11732 5472
rect 11796 5408 11812 5472
rect 11876 5408 11892 5472
rect 11956 5408 11972 5472
rect 12036 5408 12044 5472
rect 11644 4384 12044 5408
rect 11644 4320 11652 4384
rect 11716 4320 11732 4384
rect 11796 4320 11812 4384
rect 11876 4320 11892 4384
rect 11956 4320 11972 4384
rect 12036 4320 12044 4384
rect 11644 3296 12044 4320
rect 11644 3232 11652 3296
rect 11716 3232 11732 3296
rect 11796 3232 11812 3296
rect 11876 3232 11892 3296
rect 11956 3232 11972 3296
rect 12036 3232 12044 3296
rect 11644 2208 12044 3232
rect 11644 2144 11652 2208
rect 11716 2144 11732 2208
rect 11796 2144 11812 2208
rect 11876 2144 11892 2208
rect 11956 2144 11972 2208
rect 12036 2144 12044 2208
rect 11644 2128 12044 2144
rect 18904 27776 19304 27792
rect 18904 27712 18912 27776
rect 18976 27712 18992 27776
rect 19056 27712 19072 27776
rect 19136 27712 19152 27776
rect 19216 27712 19232 27776
rect 19296 27712 19304 27776
rect 18904 26688 19304 27712
rect 18904 26624 18912 26688
rect 18976 26624 18992 26688
rect 19056 26624 19072 26688
rect 19136 26624 19152 26688
rect 19216 26624 19232 26688
rect 19296 26624 19304 26688
rect 18904 25600 19304 26624
rect 18904 25536 18912 25600
rect 18976 25536 18992 25600
rect 19056 25536 19072 25600
rect 19136 25536 19152 25600
rect 19216 25536 19232 25600
rect 19296 25536 19304 25600
rect 18904 24512 19304 25536
rect 18904 24448 18912 24512
rect 18976 24448 18992 24512
rect 19056 24448 19072 24512
rect 19136 24448 19152 24512
rect 19216 24448 19232 24512
rect 19296 24448 19304 24512
rect 18904 23424 19304 24448
rect 18904 23360 18912 23424
rect 18976 23360 18992 23424
rect 19056 23360 19072 23424
rect 19136 23360 19152 23424
rect 19216 23360 19232 23424
rect 19296 23360 19304 23424
rect 18904 22336 19304 23360
rect 18904 22272 18912 22336
rect 18976 22272 18992 22336
rect 19056 22272 19072 22336
rect 19136 22272 19152 22336
rect 19216 22272 19232 22336
rect 19296 22272 19304 22336
rect 18904 21248 19304 22272
rect 18904 21184 18912 21248
rect 18976 21184 18992 21248
rect 19056 21184 19072 21248
rect 19136 21184 19152 21248
rect 19216 21184 19232 21248
rect 19296 21184 19304 21248
rect 18904 20160 19304 21184
rect 18904 20096 18912 20160
rect 18976 20096 18992 20160
rect 19056 20096 19072 20160
rect 19136 20096 19152 20160
rect 19216 20096 19232 20160
rect 19296 20096 19304 20160
rect 18904 19072 19304 20096
rect 18904 19008 18912 19072
rect 18976 19008 18992 19072
rect 19056 19008 19072 19072
rect 19136 19008 19152 19072
rect 19216 19008 19232 19072
rect 19296 19008 19304 19072
rect 18904 17984 19304 19008
rect 18904 17920 18912 17984
rect 18976 17920 18992 17984
rect 19056 17920 19072 17984
rect 19136 17920 19152 17984
rect 19216 17920 19232 17984
rect 19296 17920 19304 17984
rect 18904 16896 19304 17920
rect 18904 16832 18912 16896
rect 18976 16832 18992 16896
rect 19056 16832 19072 16896
rect 19136 16832 19152 16896
rect 19216 16832 19232 16896
rect 19296 16832 19304 16896
rect 18904 15808 19304 16832
rect 18904 15744 18912 15808
rect 18976 15744 18992 15808
rect 19056 15744 19072 15808
rect 19136 15744 19152 15808
rect 19216 15744 19232 15808
rect 19296 15744 19304 15808
rect 18904 14720 19304 15744
rect 18904 14656 18912 14720
rect 18976 14656 18992 14720
rect 19056 14656 19072 14720
rect 19136 14656 19152 14720
rect 19216 14656 19232 14720
rect 19296 14656 19304 14720
rect 18904 13632 19304 14656
rect 18904 13568 18912 13632
rect 18976 13568 18992 13632
rect 19056 13568 19072 13632
rect 19136 13568 19152 13632
rect 19216 13568 19232 13632
rect 19296 13568 19304 13632
rect 18904 12544 19304 13568
rect 18904 12480 18912 12544
rect 18976 12480 18992 12544
rect 19056 12480 19072 12544
rect 19136 12480 19152 12544
rect 19216 12480 19232 12544
rect 19296 12480 19304 12544
rect 18904 11456 19304 12480
rect 18904 11392 18912 11456
rect 18976 11392 18992 11456
rect 19056 11392 19072 11456
rect 19136 11392 19152 11456
rect 19216 11392 19232 11456
rect 19296 11392 19304 11456
rect 18904 10368 19304 11392
rect 18904 10304 18912 10368
rect 18976 10304 18992 10368
rect 19056 10304 19072 10368
rect 19136 10304 19152 10368
rect 19216 10304 19232 10368
rect 19296 10304 19304 10368
rect 18904 9280 19304 10304
rect 18904 9216 18912 9280
rect 18976 9216 18992 9280
rect 19056 9216 19072 9280
rect 19136 9216 19152 9280
rect 19216 9216 19232 9280
rect 19296 9216 19304 9280
rect 18904 8192 19304 9216
rect 18904 8128 18912 8192
rect 18976 8128 18992 8192
rect 19056 8128 19072 8192
rect 19136 8128 19152 8192
rect 19216 8128 19232 8192
rect 19296 8128 19304 8192
rect 18904 7104 19304 8128
rect 18904 7040 18912 7104
rect 18976 7040 18992 7104
rect 19056 7040 19072 7104
rect 19136 7040 19152 7104
rect 19216 7040 19232 7104
rect 19296 7040 19304 7104
rect 18904 6016 19304 7040
rect 18904 5952 18912 6016
rect 18976 5952 18992 6016
rect 19056 5952 19072 6016
rect 19136 5952 19152 6016
rect 19216 5952 19232 6016
rect 19296 5952 19304 6016
rect 18904 4928 19304 5952
rect 18904 4864 18912 4928
rect 18976 4864 18992 4928
rect 19056 4864 19072 4928
rect 19136 4864 19152 4928
rect 19216 4864 19232 4928
rect 19296 4864 19304 4928
rect 18904 3840 19304 4864
rect 18904 3776 18912 3840
rect 18976 3776 18992 3840
rect 19056 3776 19072 3840
rect 19136 3776 19152 3840
rect 19216 3776 19232 3840
rect 19296 3776 19304 3840
rect 18904 2752 19304 3776
rect 18904 2688 18912 2752
rect 18976 2688 18992 2752
rect 19056 2688 19072 2752
rect 19136 2688 19152 2752
rect 19216 2688 19232 2752
rect 19296 2688 19304 2752
rect 18904 2128 19304 2688
rect 19644 27232 20044 27792
rect 19644 27168 19652 27232
rect 19716 27168 19732 27232
rect 19796 27168 19812 27232
rect 19876 27168 19892 27232
rect 19956 27168 19972 27232
rect 20036 27168 20044 27232
rect 19644 26144 20044 27168
rect 19644 26080 19652 26144
rect 19716 26080 19732 26144
rect 19796 26080 19812 26144
rect 19876 26080 19892 26144
rect 19956 26080 19972 26144
rect 20036 26080 20044 26144
rect 19644 25056 20044 26080
rect 19644 24992 19652 25056
rect 19716 24992 19732 25056
rect 19796 24992 19812 25056
rect 19876 24992 19892 25056
rect 19956 24992 19972 25056
rect 20036 24992 20044 25056
rect 19644 23968 20044 24992
rect 19644 23904 19652 23968
rect 19716 23904 19732 23968
rect 19796 23904 19812 23968
rect 19876 23904 19892 23968
rect 19956 23904 19972 23968
rect 20036 23904 20044 23968
rect 19644 22880 20044 23904
rect 19644 22816 19652 22880
rect 19716 22816 19732 22880
rect 19796 22816 19812 22880
rect 19876 22816 19892 22880
rect 19956 22816 19972 22880
rect 20036 22816 20044 22880
rect 19644 21792 20044 22816
rect 19644 21728 19652 21792
rect 19716 21728 19732 21792
rect 19796 21728 19812 21792
rect 19876 21728 19892 21792
rect 19956 21728 19972 21792
rect 20036 21728 20044 21792
rect 19644 20704 20044 21728
rect 19644 20640 19652 20704
rect 19716 20640 19732 20704
rect 19796 20640 19812 20704
rect 19876 20640 19892 20704
rect 19956 20640 19972 20704
rect 20036 20640 20044 20704
rect 19644 19616 20044 20640
rect 19644 19552 19652 19616
rect 19716 19552 19732 19616
rect 19796 19552 19812 19616
rect 19876 19552 19892 19616
rect 19956 19552 19972 19616
rect 20036 19552 20044 19616
rect 19644 18528 20044 19552
rect 19644 18464 19652 18528
rect 19716 18464 19732 18528
rect 19796 18464 19812 18528
rect 19876 18464 19892 18528
rect 19956 18464 19972 18528
rect 20036 18464 20044 18528
rect 19644 17440 20044 18464
rect 19644 17376 19652 17440
rect 19716 17376 19732 17440
rect 19796 17376 19812 17440
rect 19876 17376 19892 17440
rect 19956 17376 19972 17440
rect 20036 17376 20044 17440
rect 19644 16352 20044 17376
rect 19644 16288 19652 16352
rect 19716 16288 19732 16352
rect 19796 16288 19812 16352
rect 19876 16288 19892 16352
rect 19956 16288 19972 16352
rect 20036 16288 20044 16352
rect 19644 15264 20044 16288
rect 19644 15200 19652 15264
rect 19716 15200 19732 15264
rect 19796 15200 19812 15264
rect 19876 15200 19892 15264
rect 19956 15200 19972 15264
rect 20036 15200 20044 15264
rect 19644 14176 20044 15200
rect 19644 14112 19652 14176
rect 19716 14112 19732 14176
rect 19796 14112 19812 14176
rect 19876 14112 19892 14176
rect 19956 14112 19972 14176
rect 20036 14112 20044 14176
rect 19644 13088 20044 14112
rect 19644 13024 19652 13088
rect 19716 13024 19732 13088
rect 19796 13024 19812 13088
rect 19876 13024 19892 13088
rect 19956 13024 19972 13088
rect 20036 13024 20044 13088
rect 19644 12000 20044 13024
rect 19644 11936 19652 12000
rect 19716 11936 19732 12000
rect 19796 11936 19812 12000
rect 19876 11936 19892 12000
rect 19956 11936 19972 12000
rect 20036 11936 20044 12000
rect 19644 10912 20044 11936
rect 19644 10848 19652 10912
rect 19716 10848 19732 10912
rect 19796 10848 19812 10912
rect 19876 10848 19892 10912
rect 19956 10848 19972 10912
rect 20036 10848 20044 10912
rect 19644 9824 20044 10848
rect 19644 9760 19652 9824
rect 19716 9760 19732 9824
rect 19796 9760 19812 9824
rect 19876 9760 19892 9824
rect 19956 9760 19972 9824
rect 20036 9760 20044 9824
rect 19644 8736 20044 9760
rect 19644 8672 19652 8736
rect 19716 8672 19732 8736
rect 19796 8672 19812 8736
rect 19876 8672 19892 8736
rect 19956 8672 19972 8736
rect 20036 8672 20044 8736
rect 19644 7648 20044 8672
rect 19644 7584 19652 7648
rect 19716 7584 19732 7648
rect 19796 7584 19812 7648
rect 19876 7584 19892 7648
rect 19956 7584 19972 7648
rect 20036 7584 20044 7648
rect 19644 6560 20044 7584
rect 19644 6496 19652 6560
rect 19716 6496 19732 6560
rect 19796 6496 19812 6560
rect 19876 6496 19892 6560
rect 19956 6496 19972 6560
rect 20036 6496 20044 6560
rect 19644 5472 20044 6496
rect 19644 5408 19652 5472
rect 19716 5408 19732 5472
rect 19796 5408 19812 5472
rect 19876 5408 19892 5472
rect 19956 5408 19972 5472
rect 20036 5408 20044 5472
rect 19644 4384 20044 5408
rect 19644 4320 19652 4384
rect 19716 4320 19732 4384
rect 19796 4320 19812 4384
rect 19876 4320 19892 4384
rect 19956 4320 19972 4384
rect 20036 4320 20044 4384
rect 19644 3296 20044 4320
rect 19644 3232 19652 3296
rect 19716 3232 19732 3296
rect 19796 3232 19812 3296
rect 19876 3232 19892 3296
rect 19956 3232 19972 3296
rect 20036 3232 20044 3296
rect 19644 2208 20044 3232
rect 19644 2144 19652 2208
rect 19716 2144 19732 2208
rect 19796 2144 19812 2208
rect 19876 2144 19892 2208
rect 19956 2144 19972 2208
rect 20036 2144 20044 2208
rect 19644 2128 20044 2144
rect 26904 27776 27304 27792
rect 26904 27712 26912 27776
rect 26976 27712 26992 27776
rect 27056 27712 27072 27776
rect 27136 27712 27152 27776
rect 27216 27712 27232 27776
rect 27296 27712 27304 27776
rect 26904 26688 27304 27712
rect 26904 26624 26912 26688
rect 26976 26624 26992 26688
rect 27056 26624 27072 26688
rect 27136 26624 27152 26688
rect 27216 26624 27232 26688
rect 27296 26624 27304 26688
rect 26904 25600 27304 26624
rect 26904 25536 26912 25600
rect 26976 25536 26992 25600
rect 27056 25536 27072 25600
rect 27136 25536 27152 25600
rect 27216 25536 27232 25600
rect 27296 25536 27304 25600
rect 26904 24512 27304 25536
rect 26904 24448 26912 24512
rect 26976 24448 26992 24512
rect 27056 24448 27072 24512
rect 27136 24448 27152 24512
rect 27216 24448 27232 24512
rect 27296 24448 27304 24512
rect 26904 23424 27304 24448
rect 26904 23360 26912 23424
rect 26976 23360 26992 23424
rect 27056 23360 27072 23424
rect 27136 23360 27152 23424
rect 27216 23360 27232 23424
rect 27296 23360 27304 23424
rect 26904 22336 27304 23360
rect 26904 22272 26912 22336
rect 26976 22272 26992 22336
rect 27056 22272 27072 22336
rect 27136 22272 27152 22336
rect 27216 22272 27232 22336
rect 27296 22272 27304 22336
rect 26904 21248 27304 22272
rect 26904 21184 26912 21248
rect 26976 21184 26992 21248
rect 27056 21184 27072 21248
rect 27136 21184 27152 21248
rect 27216 21184 27232 21248
rect 27296 21184 27304 21248
rect 26904 20160 27304 21184
rect 26904 20096 26912 20160
rect 26976 20096 26992 20160
rect 27056 20096 27072 20160
rect 27136 20096 27152 20160
rect 27216 20096 27232 20160
rect 27296 20096 27304 20160
rect 26904 19072 27304 20096
rect 26904 19008 26912 19072
rect 26976 19008 26992 19072
rect 27056 19008 27072 19072
rect 27136 19008 27152 19072
rect 27216 19008 27232 19072
rect 27296 19008 27304 19072
rect 26904 17984 27304 19008
rect 26904 17920 26912 17984
rect 26976 17920 26992 17984
rect 27056 17920 27072 17984
rect 27136 17920 27152 17984
rect 27216 17920 27232 17984
rect 27296 17920 27304 17984
rect 26904 16896 27304 17920
rect 26904 16832 26912 16896
rect 26976 16832 26992 16896
rect 27056 16832 27072 16896
rect 27136 16832 27152 16896
rect 27216 16832 27232 16896
rect 27296 16832 27304 16896
rect 26904 15808 27304 16832
rect 26904 15744 26912 15808
rect 26976 15744 26992 15808
rect 27056 15744 27072 15808
rect 27136 15744 27152 15808
rect 27216 15744 27232 15808
rect 27296 15744 27304 15808
rect 26904 14720 27304 15744
rect 26904 14656 26912 14720
rect 26976 14656 26992 14720
rect 27056 14656 27072 14720
rect 27136 14656 27152 14720
rect 27216 14656 27232 14720
rect 27296 14656 27304 14720
rect 26904 13632 27304 14656
rect 26904 13568 26912 13632
rect 26976 13568 26992 13632
rect 27056 13568 27072 13632
rect 27136 13568 27152 13632
rect 27216 13568 27232 13632
rect 27296 13568 27304 13632
rect 26904 12544 27304 13568
rect 26904 12480 26912 12544
rect 26976 12480 26992 12544
rect 27056 12480 27072 12544
rect 27136 12480 27152 12544
rect 27216 12480 27232 12544
rect 27296 12480 27304 12544
rect 26904 11456 27304 12480
rect 26904 11392 26912 11456
rect 26976 11392 26992 11456
rect 27056 11392 27072 11456
rect 27136 11392 27152 11456
rect 27216 11392 27232 11456
rect 27296 11392 27304 11456
rect 26904 10368 27304 11392
rect 26904 10304 26912 10368
rect 26976 10304 26992 10368
rect 27056 10304 27072 10368
rect 27136 10304 27152 10368
rect 27216 10304 27232 10368
rect 27296 10304 27304 10368
rect 26904 9280 27304 10304
rect 26904 9216 26912 9280
rect 26976 9216 26992 9280
rect 27056 9216 27072 9280
rect 27136 9216 27152 9280
rect 27216 9216 27232 9280
rect 27296 9216 27304 9280
rect 26904 8192 27304 9216
rect 26904 8128 26912 8192
rect 26976 8128 26992 8192
rect 27056 8128 27072 8192
rect 27136 8128 27152 8192
rect 27216 8128 27232 8192
rect 27296 8128 27304 8192
rect 26904 7104 27304 8128
rect 26904 7040 26912 7104
rect 26976 7040 26992 7104
rect 27056 7040 27072 7104
rect 27136 7040 27152 7104
rect 27216 7040 27232 7104
rect 27296 7040 27304 7104
rect 26904 6016 27304 7040
rect 26904 5952 26912 6016
rect 26976 5952 26992 6016
rect 27056 5952 27072 6016
rect 27136 5952 27152 6016
rect 27216 5952 27232 6016
rect 27296 5952 27304 6016
rect 26904 4928 27304 5952
rect 26904 4864 26912 4928
rect 26976 4864 26992 4928
rect 27056 4864 27072 4928
rect 27136 4864 27152 4928
rect 27216 4864 27232 4928
rect 27296 4864 27304 4928
rect 26904 3840 27304 4864
rect 26904 3776 26912 3840
rect 26976 3776 26992 3840
rect 27056 3776 27072 3840
rect 27136 3776 27152 3840
rect 27216 3776 27232 3840
rect 27296 3776 27304 3840
rect 26904 2752 27304 3776
rect 26904 2688 26912 2752
rect 26976 2688 26992 2752
rect 27056 2688 27072 2752
rect 27136 2688 27152 2752
rect 27216 2688 27232 2752
rect 27296 2688 27304 2752
rect 26904 2128 27304 2688
rect 27644 27232 28044 27792
rect 27644 27168 27652 27232
rect 27716 27168 27732 27232
rect 27796 27168 27812 27232
rect 27876 27168 27892 27232
rect 27956 27168 27972 27232
rect 28036 27168 28044 27232
rect 27644 26144 28044 27168
rect 27644 26080 27652 26144
rect 27716 26080 27732 26144
rect 27796 26080 27812 26144
rect 27876 26080 27892 26144
rect 27956 26080 27972 26144
rect 28036 26080 28044 26144
rect 27644 25056 28044 26080
rect 27644 24992 27652 25056
rect 27716 24992 27732 25056
rect 27796 24992 27812 25056
rect 27876 24992 27892 25056
rect 27956 24992 27972 25056
rect 28036 24992 28044 25056
rect 27644 23968 28044 24992
rect 27644 23904 27652 23968
rect 27716 23904 27732 23968
rect 27796 23904 27812 23968
rect 27876 23904 27892 23968
rect 27956 23904 27972 23968
rect 28036 23904 28044 23968
rect 27644 22880 28044 23904
rect 27644 22816 27652 22880
rect 27716 22816 27732 22880
rect 27796 22816 27812 22880
rect 27876 22816 27892 22880
rect 27956 22816 27972 22880
rect 28036 22816 28044 22880
rect 27644 21792 28044 22816
rect 27644 21728 27652 21792
rect 27716 21728 27732 21792
rect 27796 21728 27812 21792
rect 27876 21728 27892 21792
rect 27956 21728 27972 21792
rect 28036 21728 28044 21792
rect 27644 20704 28044 21728
rect 27644 20640 27652 20704
rect 27716 20640 27732 20704
rect 27796 20640 27812 20704
rect 27876 20640 27892 20704
rect 27956 20640 27972 20704
rect 28036 20640 28044 20704
rect 27644 19616 28044 20640
rect 27644 19552 27652 19616
rect 27716 19552 27732 19616
rect 27796 19552 27812 19616
rect 27876 19552 27892 19616
rect 27956 19552 27972 19616
rect 28036 19552 28044 19616
rect 27644 18528 28044 19552
rect 27644 18464 27652 18528
rect 27716 18464 27732 18528
rect 27796 18464 27812 18528
rect 27876 18464 27892 18528
rect 27956 18464 27972 18528
rect 28036 18464 28044 18528
rect 27644 17440 28044 18464
rect 27644 17376 27652 17440
rect 27716 17376 27732 17440
rect 27796 17376 27812 17440
rect 27876 17376 27892 17440
rect 27956 17376 27972 17440
rect 28036 17376 28044 17440
rect 27644 16352 28044 17376
rect 27644 16288 27652 16352
rect 27716 16288 27732 16352
rect 27796 16288 27812 16352
rect 27876 16288 27892 16352
rect 27956 16288 27972 16352
rect 28036 16288 28044 16352
rect 27644 15264 28044 16288
rect 27644 15200 27652 15264
rect 27716 15200 27732 15264
rect 27796 15200 27812 15264
rect 27876 15200 27892 15264
rect 27956 15200 27972 15264
rect 28036 15200 28044 15264
rect 27644 14176 28044 15200
rect 27644 14112 27652 14176
rect 27716 14112 27732 14176
rect 27796 14112 27812 14176
rect 27876 14112 27892 14176
rect 27956 14112 27972 14176
rect 28036 14112 28044 14176
rect 27644 13088 28044 14112
rect 27644 13024 27652 13088
rect 27716 13024 27732 13088
rect 27796 13024 27812 13088
rect 27876 13024 27892 13088
rect 27956 13024 27972 13088
rect 28036 13024 28044 13088
rect 27644 12000 28044 13024
rect 27644 11936 27652 12000
rect 27716 11936 27732 12000
rect 27796 11936 27812 12000
rect 27876 11936 27892 12000
rect 27956 11936 27972 12000
rect 28036 11936 28044 12000
rect 27644 10912 28044 11936
rect 27644 10848 27652 10912
rect 27716 10848 27732 10912
rect 27796 10848 27812 10912
rect 27876 10848 27892 10912
rect 27956 10848 27972 10912
rect 28036 10848 28044 10912
rect 27644 9824 28044 10848
rect 27644 9760 27652 9824
rect 27716 9760 27732 9824
rect 27796 9760 27812 9824
rect 27876 9760 27892 9824
rect 27956 9760 27972 9824
rect 28036 9760 28044 9824
rect 27644 8736 28044 9760
rect 27644 8672 27652 8736
rect 27716 8672 27732 8736
rect 27796 8672 27812 8736
rect 27876 8672 27892 8736
rect 27956 8672 27972 8736
rect 28036 8672 28044 8736
rect 27644 7648 28044 8672
rect 27644 7584 27652 7648
rect 27716 7584 27732 7648
rect 27796 7584 27812 7648
rect 27876 7584 27892 7648
rect 27956 7584 27972 7648
rect 28036 7584 28044 7648
rect 27644 6560 28044 7584
rect 27644 6496 27652 6560
rect 27716 6496 27732 6560
rect 27796 6496 27812 6560
rect 27876 6496 27892 6560
rect 27956 6496 27972 6560
rect 28036 6496 28044 6560
rect 27644 5472 28044 6496
rect 27644 5408 27652 5472
rect 27716 5408 27732 5472
rect 27796 5408 27812 5472
rect 27876 5408 27892 5472
rect 27956 5408 27972 5472
rect 28036 5408 28044 5472
rect 27644 4384 28044 5408
rect 27644 4320 27652 4384
rect 27716 4320 27732 4384
rect 27796 4320 27812 4384
rect 27876 4320 27892 4384
rect 27956 4320 27972 4384
rect 28036 4320 28044 4384
rect 27644 3296 28044 4320
rect 27644 3232 27652 3296
rect 27716 3232 27732 3296
rect 27796 3232 27812 3296
rect 27876 3232 27892 3296
rect 27956 3232 27972 3296
rect 28036 3232 28044 3296
rect 27644 2208 28044 3232
rect 27644 2144 27652 2208
rect 27716 2144 27732 2208
rect 27796 2144 27812 2208
rect 27876 2144 27892 2208
rect 27956 2144 27972 2208
rect 28036 2144 28044 2208
rect 27644 2128 28044 2144
use sky130_fd_sc_hd__mux2_1  _32_
timestamp -25199
transform -1 0 11408 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _33_
timestamp -25199
transform 1 0 12420 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _34_
timestamp -25199
transform 1 0 12420 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _35_
timestamp -25199
transform 1 0 11500 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _36_
timestamp -25199
transform -1 0 10580 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _37_
timestamp -25199
transform -1 0 11408 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _38_
timestamp -25199
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _39_
timestamp -25199
transform -1 0 11408 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _40_
timestamp -25199
transform -1 0 11408 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _41_
timestamp -25199
transform 1 0 12604 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _42_
timestamp -25199
transform 1 0 11500 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _43_
timestamp -25199
transform -1 0 11408 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _44_
timestamp -25199
transform -1 0 11408 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _45_
timestamp -25199
transform 1 0 12512 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _46_
timestamp -25199
transform 1 0 11500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _47_
timestamp -25199
transform 1 0 10580 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _48_
timestamp -25199
transform 1 0 11500 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _49_
timestamp -25199
transform 1 0 14076 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _50_
timestamp -25199
transform 1 0 11500 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _51_
timestamp -25199
transform 1 0 12972 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _52_
timestamp -25199
transform -1 0 11408 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _53_
timestamp -25199
transform 1 0 12972 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _54_
timestamp -25199
transform 1 0 11500 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _55_
timestamp -25199
transform 1 0 10580 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _56_
timestamp -25199
transform -1 0 11408 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _57_
timestamp -25199
transform 1 0 12052 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _58_
timestamp -25199
transform 1 0 14076 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _59_
timestamp -25199
transform 1 0 14076 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _60_
timestamp -25199
transform 1 0 13156 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _61_
timestamp -25199
transform 1 0 11500 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _62_
timestamp -25199
transform 1 0 14076 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _63_
timestamp -25199
transform 1 0 14076 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _64_
timestamp -25199
transform 1 0 11500 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _65_
timestamp -25199
transform 1 0 10580 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _66_
timestamp -25199
transform 1 0 11500 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _67_
timestamp -25199
transform 1 0 10580 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _68_
timestamp -25199
transform 1 0 10672 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _69_
timestamp -25199
transform 1 0 11500 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _70_
timestamp -25199
transform 1 0 10672 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _71_
timestamp -25199
transform 1 0 11500 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _72_
timestamp -25199
transform 1 0 11500 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _73_
timestamp -25199
transform 1 0 10672 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _74_
timestamp -25199
transform 1 0 10672 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _75_
timestamp -25199
transform 1 0 11500 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _76_
timestamp -25199
transform 1 0 10672 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _77_
timestamp -25199
transform 1 0 11500 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _78_
timestamp -25199
transform 1 0 10580 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _79_
timestamp -25199
transform 1 0 10580 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _80_
timestamp -25199
transform 1 0 11040 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _81_
timestamp -25199
transform 1 0 13064 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _82_
timestamp -25199
transform 1 0 11040 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _83_
timestamp -25199
transform 1 0 12052 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _84_
timestamp -25199
transform 1 0 11040 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _85_
timestamp -25199
transform 1 0 11684 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _86_
timestamp -25199
transform 1 0 11040 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _87_
timestamp -25199
transform -1 0 11040 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _88_
timestamp -25199
transform 1 0 11500 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _89_
timestamp -25199
transform 1 0 11592 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _90_
timestamp -25199
transform 1 0 12052 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _91_
timestamp -25199
transform 1 0 12328 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _92_
timestamp -25199
transform 1 0 12604 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _93_
timestamp -25199
transform 1 0 11040 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _94_
timestamp -25199
transform 1 0 13064 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _95_
timestamp -25199
transform 1 0 13064 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -25199
transform 1 0 11500 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp -25199
transform -1 0 11408 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp -25199
transform -1 0 12880 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp -25199
transform 1 0 11500 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp -25199
transform 1 0 12144 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp -25199
transform -1 0 10672 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  clkload1
timestamp -25199
transform -1 0 11040 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  clkload2
timestamp -25199
transform 1 0 12236 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  fanout67
timestamp -25199
transform -1 0 10580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout68
timestamp -25199
transform 1 0 10212 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout69
timestamp -25199
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout70
timestamp -25199
transform -1 0 11132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout71
timestamp -25199
transform 1 0 11132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout72
timestamp -25199
transform -1 0 11776 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout73
timestamp -25199
transform 1 0 11500 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout74
timestamp -25199
transform -1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout75
timestamp -25199
transform -1 0 12144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout76
timestamp -25199
transform -1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout77
timestamp -25199
transform -1 0 12880 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout78
timestamp -25199
transform 1 0 12328 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout79
timestamp -25199
transform -1 0 12604 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout80
timestamp -25199
transform 1 0 11132 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6
timestamp 1636943256
transform 1 0 1656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18
timestamp -25199
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp -25199
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636943256
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636943256
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -25199
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636943256
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636943256
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -25199
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636943256
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636943256
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -25199
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp -25199
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120
timestamp 1636943256
transform 1 0 12144 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132
timestamp -25199
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636943256
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636943256
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -25199
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636943256
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636943256
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -25199
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636943256
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636943256
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -25199
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636943256
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636943256
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -25199
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636943256
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636943256
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -25199
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636943256
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6
timestamp 1636943256
transform 1 0 1656 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_18
timestamp 1636943256
transform 1 0 2760 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_30
timestamp 1636943256
transform 1 0 3864 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_42
timestamp 1636943256
transform 1 0 4968 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp -25199
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636943256
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636943256
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636943256
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_93
timestamp -25199
transform 1 0 9660 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_101
timestamp -25199
transform 1 0 10396 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_133
timestamp 1636943256
transform 1 0 13340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_145
timestamp 1636943256
transform 1 0 14444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_157
timestamp -25199
transform 1 0 15548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp -25199
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636943256
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636943256
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636943256
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636943256
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp -25199
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp -25199
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636943256
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636943256
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636943256
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636943256
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp -25199
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp -25199
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636943256
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_293
timestamp -25199
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6
timestamp 1636943256
transform 1 0 1656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp -25199
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp -25199
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636943256
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636943256
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636943256
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636943256
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp -25199
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -25199
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636943256
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_97
timestamp -25199
transform 1 0 10028 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp -25199
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636943256
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636943256
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636943256
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636943256
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp -25199
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp -25199
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636943256
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636943256
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636943256
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636943256
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp -25199
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp -25199
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636943256
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636943256
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636943256
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_289
timestamp -25199
transform 1 0 27692 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636943256
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636943256
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636943256
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636943256
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp -25199
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -25199
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636943256
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636943256
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636943256
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636943256
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_105
timestamp -25199
transform 1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_133
timestamp 1636943256
transform 1 0 13340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_145
timestamp 1636943256
transform 1 0 14444 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_157
timestamp -25199
transform 1 0 15548 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_165
timestamp -25199
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636943256
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636943256
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636943256
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636943256
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp -25199
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp -25199
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636943256
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636943256
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636943256
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636943256
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp -25199
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp -25199
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636943256
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_6
timestamp 1636943256
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_18
timestamp -25199
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp -25199
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636943256
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636943256
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636943256
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636943256
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp -25199
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -25199
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636943256
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_97
timestamp -25199
transform 1 0 10028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_132
timestamp -25199
transform 1 0 13248 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636943256
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636943256
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636943256
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636943256
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp -25199
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp -25199
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636943256
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636943256
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636943256
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636943256
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp -25199
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp -25199
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636943256
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636943256
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636943256
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_289
timestamp -25199
transform 1 0 27692 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_297
timestamp -25199
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6
timestamp 1636943256
transform 1 0 1656 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_18
timestamp 1636943256
transform 1 0 2760 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_30
timestamp 1636943256
transform 1 0 3864 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_42
timestamp 1636943256
transform 1 0 4968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp -25199
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636943256
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636943256
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636943256
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636943256
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp -25199
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -25199
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_122
timestamp 1636943256
transform 1 0 12328 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_134
timestamp 1636943256
transform 1 0 13432 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_146
timestamp 1636943256
transform 1 0 14536 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_158
timestamp -25199
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp -25199
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636943256
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636943256
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636943256
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636943256
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp -25199
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp -25199
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636943256
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636943256
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636943256
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636943256
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp -25199
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp -25199
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636943256
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636943256
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636943256
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -25199
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636943256
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636943256
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636943256
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636943256
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp -25199
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp -25199
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636943256
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_97
timestamp -25199
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_103
timestamp -25199
transform 1 0 10580 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_124
timestamp 1636943256
transform 1 0 12512 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp -25199
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636943256
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636943256
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636943256
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636943256
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp -25199
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp -25199
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636943256
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636943256
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1636943256
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1636943256
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp -25199
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp -25199
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636943256
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636943256
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1636943256
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_289
timestamp -25199
transform 1 0 27692 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_6
timestamp 1636943256
transform 1 0 1656 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_18
timestamp 1636943256
transform 1 0 2760 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_30
timestamp 1636943256
transform 1 0 3864 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_42
timestamp 1636943256
transform 1 0 4968 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp -25199
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636943256
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636943256
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636943256
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_93
timestamp -25199
transform 1 0 9660 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_133
timestamp 1636943256
transform 1 0 13340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_145
timestamp 1636943256
transform 1 0 14444 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_157
timestamp -25199
transform 1 0 15548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp -25199
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636943256
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636943256
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636943256
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1636943256
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp -25199
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp -25199
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636943256
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636943256
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636943256
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1636943256
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp -25199
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp -25199
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636943256
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp -25199
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_6
timestamp 1636943256
transform 1 0 1656 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_18
timestamp -25199
transform 1 0 2760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp -25199
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636943256
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636943256
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636943256
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636943256
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp -25199
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp -25199
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636943256
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_97
timestamp -25199
transform 1 0 10028 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_101
timestamp -25199
transform 1 0 10396 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_128
timestamp 1636943256
transform 1 0 12880 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636943256
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636943256
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636943256
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1636943256
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp -25199
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp -25199
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636943256
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636943256
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1636943256
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1636943256
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp -25199
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp -25199
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636943256
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1636943256
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1636943256
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_289
timestamp -25199
transform 1 0 27692 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636943256
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636943256
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636943256
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1636943256
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp -25199
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -25199
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636943256
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636943256
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636943256
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1636943256
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp -25199
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp -25199
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_122
timestamp 1636943256
transform 1 0 12328 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_134
timestamp 1636943256
transform 1 0 13432 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_146
timestamp 1636943256
transform 1 0 14536 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_158
timestamp -25199
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp -25199
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636943256
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1636943256
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1636943256
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1636943256
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp -25199
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp -25199
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636943256
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1636943256
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1636943256
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1636943256
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp -25199
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp -25199
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636943256
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_6
timestamp 1636943256
transform 1 0 1656 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_18
timestamp -25199
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp -25199
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636943256
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636943256
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636943256
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1636943256
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp -25199
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp -25199
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636943256
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_97
timestamp -25199
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_103
timestamp -25199
transform 1 0 10580 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_124
timestamp 1636943256
transform 1 0 12512 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp -25199
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636943256
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1636943256
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1636943256
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1636943256
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp -25199
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp -25199
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1636943256
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1636943256
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1636943256
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1636943256
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp -25199
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp -25199
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1636943256
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1636943256
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1636943256
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_289
timestamp -25199
transform 1 0 27692 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_297
timestamp -25199
transform 1 0 28428 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_6
timestamp 1636943256
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_18
timestamp 1636943256
transform 1 0 2760 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_30
timestamp 1636943256
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_42
timestamp 1636943256
transform 1 0 4968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp -25199
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636943256
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1636943256
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1636943256
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_93
timestamp -25199
transform 1 0 9660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp -25199
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_133
timestamp 1636943256
transform 1 0 13340 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_145
timestamp 1636943256
transform 1 0 14444 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_157
timestamp -25199
transform 1 0 15548 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp -25199
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1636943256
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1636943256
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1636943256
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1636943256
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp -25199
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp -25199
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1636943256
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1636943256
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1636943256
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1636943256
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp -25199
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp -25199
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1636943256
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636943256
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636943256
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp -25199
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636943256
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636943256
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1636943256
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1636943256
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp -25199
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp -25199
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1636943256
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1636943256
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_109
timestamp -25199
transform 1 0 11132 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_115
timestamp -25199
transform 1 0 11684 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_120
timestamp 1636943256
transform 1 0 12144 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_132
timestamp -25199
transform 1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1636943256
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1636943256
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1636943256
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1636943256
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp -25199
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp -25199
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1636943256
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1636943256
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1636943256
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1636943256
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp -25199
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp -25199
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1636943256
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1636943256
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1636943256
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_289
timestamp -25199
transform 1 0 27692 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_6
timestamp 1636943256
transform 1 0 1656 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_18
timestamp 1636943256
transform 1 0 2760 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_30
timestamp 1636943256
transform 1 0 3864 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_42
timestamp 1636943256
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp -25199
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636943256
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1636943256
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1636943256
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_93
timestamp -25199
transform 1 0 9660 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp -25199
transform 1 0 10396 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_134
timestamp 1636943256
transform 1 0 13432 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_146
timestamp 1636943256
transform 1 0 14536 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_158
timestamp -25199
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp -25199
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1636943256
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1636943256
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1636943256
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1636943256
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp -25199
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp -25199
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1636943256
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1636943256
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1636943256
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1636943256
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp -25199
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp -25199
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1636943256
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_293
timestamp -25199
transform 1 0 28060 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_6
timestamp 1636943256
transform 1 0 1656 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_18
timestamp -25199
transform 1 0 2760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp -25199
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636943256
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636943256
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1636943256
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1636943256
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp -25199
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp -25199
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1636943256
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_97
timestamp -25199
transform 1 0 10028 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_103
timestamp -25199
transform 1 0 10580 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_134
timestamp -25199
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1636943256
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1636943256
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1636943256
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1636943256
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp -25199
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp -25199
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1636943256
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1636943256
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1636943256
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1636943256
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp -25199
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp -25199
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1636943256
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1636943256
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1636943256
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_289
timestamp -25199
transform 1 0 27692 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636943256
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636943256
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636943256
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1636943256
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp -25199
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp -25199
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636943256
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1636943256
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1636943256
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_93
timestamp -25199
transform 1 0 9660 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_122
timestamp 1636943256
transform 1 0 12328 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_134
timestamp 1636943256
transform 1 0 13432 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_146
timestamp 1636943256
transform 1 0 14536 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_158
timestamp -25199
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp -25199
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1636943256
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1636943256
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1636943256
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1636943256
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp -25199
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp -25199
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1636943256
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1636943256
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1636943256
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1636943256
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp -25199
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp -25199
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1636943256
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_6
timestamp 1636943256
transform 1 0 1656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_18
timestamp -25199
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp -25199
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636943256
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1636943256
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1636943256
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1636943256
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp -25199
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp -25199
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1636943256
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_97
timestamp -25199
transform 1 0 10028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_103
timestamp -25199
transform 1 0 10580 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_125
timestamp 1636943256
transform 1 0 12604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp -25199
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1636943256
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1636943256
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1636943256
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1636943256
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp -25199
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp -25199
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1636943256
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1636943256
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1636943256
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1636943256
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp -25199
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp -25199
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1636943256
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1636943256
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1636943256
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_289
timestamp -25199
transform 1 0 27692 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp -25199
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_6
timestamp 1636943256
transform 1 0 1656 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_18
timestamp 1636943256
transform 1 0 2760 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_30
timestamp 1636943256
transform 1 0 3864 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_42
timestamp 1636943256
transform 1 0 4968 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp -25199
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636943256
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1636943256
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_81
timestamp -25199
transform 1 0 8556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_89
timestamp -25199
transform 1 0 9292 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_134
timestamp 1636943256
transform 1 0 13432 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_146
timestamp 1636943256
transform 1 0 14536 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_158
timestamp -25199
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp -25199
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1636943256
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1636943256
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1636943256
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1636943256
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp -25199
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp -25199
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1636943256
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1636943256
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1636943256
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1636943256
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp -25199
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp -25199
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1636943256
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636943256
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636943256
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp -25199
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636943256
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636943256
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1636943256
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1636943256
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp -25199
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp -25199
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1636943256
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_97
timestamp -25199
transform 1 0 10028 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_125
timestamp 1636943256
transform 1 0 12604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp -25199
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1636943256
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1636943256
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1636943256
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1636943256
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp -25199
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp -25199
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1636943256
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1636943256
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1636943256
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1636943256
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp -25199
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp -25199
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1636943256
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1636943256
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1636943256
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_289
timestamp -25199
transform 1 0 27692 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_6
timestamp 1636943256
transform 1 0 1656 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_18
timestamp 1636943256
transform 1 0 2760 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_30
timestamp 1636943256
transform 1 0 3864 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_42
timestamp 1636943256
transform 1 0 4968 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp -25199
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636943256
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1636943256
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1636943256
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_93
timestamp -25199
transform 1 0 9660 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp -25199
transform 1 0 10396 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_134
timestamp 1636943256
transform 1 0 13432 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_146
timestamp 1636943256
transform 1 0 14536 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_158
timestamp -25199
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp -25199
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1636943256
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1636943256
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1636943256
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1636943256
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp -25199
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp -25199
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1636943256
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1636943256
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1636943256
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1636943256
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp -25199
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp -25199
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1636943256
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp -25199
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_6
timestamp 1636943256
transform 1 0 1656 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_18
timestamp -25199
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp -25199
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636943256
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1636943256
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1636943256
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1636943256
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp -25199
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp -25199
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1636943256
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_97
timestamp -25199
transform 1 0 10028 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp -25199
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp -25199
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1636943256
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1636943256
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1636943256
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1636943256
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp -25199
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp -25199
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1636943256
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1636943256
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1636943256
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1636943256
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp -25199
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp -25199
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1636943256
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1636943256
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1636943256
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_289
timestamp -25199
transform 1 0 27692 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636943256
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636943256
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1636943256
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1636943256
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp -25199
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp -25199
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1636943256
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1636943256
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1636943256
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1636943256
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp -25199
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp -25199
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_122
timestamp 1636943256
transform 1 0 12328 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_134
timestamp 1636943256
transform 1 0 13432 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_146
timestamp 1636943256
transform 1 0 14536 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_158
timestamp -25199
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp -25199
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1636943256
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1636943256
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1636943256
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1636943256
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp -25199
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp -25199
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1636943256
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1636943256
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1636943256
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1636943256
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp -25199
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp -25199
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1636943256
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_6
timestamp 1636943256
transform 1 0 1656 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_18
timestamp -25199
transform 1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp -25199
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636943256
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1636943256
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1636943256
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1636943256
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp -25199
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp -25199
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1636943256
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_97
timestamp -25199
transform 1 0 10028 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_128
timestamp 1636943256
transform 1 0 12880 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1636943256
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1636943256
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1636943256
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1636943256
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp -25199
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp -25199
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1636943256
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1636943256
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1636943256
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1636943256
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp -25199
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp -25199
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1636943256
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1636943256
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1636943256
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_289
timestamp -25199
transform 1 0 27692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_297
timestamp -25199
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_6
timestamp 1636943256
transform 1 0 1656 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_18
timestamp 1636943256
transform 1 0 2760 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_30
timestamp 1636943256
transform 1 0 3864 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_42
timestamp 1636943256
transform 1 0 4968 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp -25199
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1636943256
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1636943256
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1636943256
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_93
timestamp -25199
transform 1 0 9660 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp -25199
transform 1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_133
timestamp 1636943256
transform 1 0 13340 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_145
timestamp 1636943256
transform 1 0 14444 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_157
timestamp -25199
transform 1 0 15548 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp -25199
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1636943256
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1636943256
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1636943256
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1636943256
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp -25199
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp -25199
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1636943256
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1636943256
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1636943256
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1636943256
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp -25199
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp -25199
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1636943256
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636943256
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636943256
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp -25199
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636943256
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1636943256
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1636943256
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1636943256
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp -25199
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp -25199
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1636943256
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_97
timestamp -25199
transform 1 0 10028 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_117
timestamp -25199
transform 1 0 11868 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_128
timestamp 1636943256
transform 1 0 12880 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1636943256
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1636943256
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1636943256
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1636943256
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp -25199
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp -25199
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1636943256
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1636943256
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1636943256
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1636943256
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp -25199
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp -25199
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1636943256
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1636943256
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1636943256
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_289
timestamp -25199
transform 1 0 27692 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_6
timestamp 1636943256
transform 1 0 1656 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_18
timestamp 1636943256
transform 1 0 2760 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_30
timestamp 1636943256
transform 1 0 3864 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_42
timestamp 1636943256
transform 1 0 4968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp -25199
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636943256
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1636943256
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1636943256
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_93
timestamp -25199
transform 1 0 9660 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp -25199
transform 1 0 10396 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_134
timestamp 1636943256
transform 1 0 13432 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_146
timestamp 1636943256
transform 1 0 14536 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_158
timestamp -25199
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp -25199
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1636943256
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1636943256
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1636943256
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1636943256
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp -25199
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp -25199
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1636943256
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1636943256
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1636943256
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1636943256
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp -25199
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp -25199
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1636943256
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_293
timestamp -25199
transform 1 0 28060 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_6
timestamp 1636943256
transform 1 0 1656 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_18
timestamp -25199
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp -25199
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636943256
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1636943256
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1636943256
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1636943256
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp -25199
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp -25199
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1636943256
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1636943256
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_109
timestamp -25199
transform 1 0 11132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_113
timestamp -25199
transform 1 0 11500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp -25199
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp -25199
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1636943256
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1636943256
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1636943256
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1636943256
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp -25199
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp -25199
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1636943256
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1636943256
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1636943256
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1636943256
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp -25199
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp -25199
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1636943256
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1636943256
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1636943256
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_289
timestamp -25199
transform 1 0 27692 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636943256
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1636943256
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1636943256
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1636943256
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp -25199
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp -25199
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1636943256
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1636943256
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1636943256
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1636943256
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp -25199
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp -25199
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_113
timestamp -25199
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_140
timestamp 1636943256
transform 1 0 13984 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_152
timestamp 1636943256
transform 1 0 15088 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp -25199
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1636943256
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1636943256
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1636943256
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1636943256
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp -25199
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp -25199
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1636943256
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1636943256
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1636943256
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1636943256
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp -25199
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp -25199
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1636943256
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_6
timestamp 1636943256
transform 1 0 1656 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_18
timestamp -25199
transform 1 0 2760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp -25199
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636943256
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636943256
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1636943256
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1636943256
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp -25199
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp -25199
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1636943256
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1636943256
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_109
timestamp -25199
transform 1 0 11132 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_117
timestamp -25199
transform 1 0 11868 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_150
timestamp 1636943256
transform 1 0 14904 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_162
timestamp 1636943256
transform 1 0 16008 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_174
timestamp 1636943256
transform 1 0 17112 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_186
timestamp -25199
transform 1 0 18216 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp -25199
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1636943256
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1636943256
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1636943256
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1636943256
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp -25199
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp -25199
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1636943256
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1636943256
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1636943256
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_289
timestamp -25199
transform 1 0 27692 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_297
timestamp -25199
transform 1 0 28428 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_6
timestamp 1636943256
transform 1 0 1656 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_18
timestamp 1636943256
transform 1 0 2760 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_30
timestamp 1636943256
transform 1 0 3864 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_42
timestamp 1636943256
transform 1 0 4968 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp -25199
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636943256
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1636943256
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1636943256
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1636943256
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp -25199
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp -25199
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp -25199
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp -25199
transform 1 0 12236 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_143
timestamp 1636943256
transform 1 0 14260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_155
timestamp 1636943256
transform 1 0 15364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp -25199
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1636943256
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1636943256
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1636943256
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1636943256
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp -25199
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp -25199
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1636943256
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1636943256
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1636943256
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1636943256
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp -25199
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp -25199
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1636943256
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636943256
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636943256
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp -25199
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1636943256
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1636943256
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1636943256
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1636943256
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp -25199
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp -25199
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1636943256
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1636943256
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1636943256
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_132
timestamp -25199
transform 1 0 13248 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_150
timestamp 1636943256
transform 1 0 14904 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_162
timestamp 1636943256
transform 1 0 16008 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_174
timestamp 1636943256
transform 1 0 17112 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_186
timestamp -25199
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp -25199
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1636943256
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1636943256
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1636943256
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1636943256
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp -25199
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp -25199
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1636943256
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1636943256
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1636943256
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_289
timestamp -25199
transform 1 0 27692 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_6
timestamp 1636943256
transform 1 0 1656 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_18
timestamp 1636943256
transform 1 0 2760 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_30
timestamp 1636943256
transform 1 0 3864 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_42
timestamp 1636943256
transform 1 0 4968 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp -25199
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1636943256
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1636943256
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1636943256
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1636943256
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp -25199
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp -25199
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_122
timestamp -25199
transform 1 0 12328 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_146
timestamp 1636943256
transform 1 0 14536 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_158
timestamp -25199
transform 1 0 15640 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp -25199
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1636943256
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1636943256
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1636943256
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1636943256
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp -25199
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp -25199
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1636943256
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1636943256
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1636943256
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1636943256
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp -25199
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp -25199
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1636943256
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp -25199
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_6
timestamp 1636943256
transform 1 0 1656 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_18
timestamp -25199
transform 1 0 2760 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp -25199
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636943256
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1636943256
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1636943256
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1636943256
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp -25199
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp -25199
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1636943256
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_97
timestamp -25199
transform 1 0 10028 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_105
timestamp -25199
transform 1 0 10764 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_129
timestamp -25199
transform 1 0 12972 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1636943256
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1636943256
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1636943256
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1636943256
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp -25199
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp -25199
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1636943256
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1636943256
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1636943256
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1636943256
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp -25199
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp -25199
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1636943256
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1636943256
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1636943256
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_289
timestamp -25199
transform 1 0 27692 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636943256
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1636943256
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1636943256
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1636943256
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp -25199
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp -25199
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1636943256
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1636943256
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1636943256
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1636943256
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp -25199
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp -25199
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1636943256
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_125
timestamp -25199
transform 1 0 12604 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_129
timestamp -25199
transform 1 0 12972 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_151
timestamp 1636943256
transform 1 0 14996 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp -25199
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp -25199
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1636943256
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1636943256
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1636943256
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1636943256
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp -25199
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp -25199
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1636943256
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1636943256
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1636943256
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1636943256
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp -25199
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp -25199
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1636943256
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_6
timestamp 1636943256
transform 1 0 1656 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_18
timestamp -25199
transform 1 0 2760 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp -25199
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1636943256
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1636943256
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1636943256
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1636943256
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp -25199
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp -25199
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1636943256
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1636943256
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1636943256
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1636943256
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp -25199
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp -25199
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_150
timestamp 1636943256
transform 1 0 14904 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_162
timestamp 1636943256
transform 1 0 16008 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_174
timestamp 1636943256
transform 1 0 17112 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_186
timestamp -25199
transform 1 0 18216 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp -25199
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1636943256
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1636943256
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1636943256
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1636943256
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp -25199
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp -25199
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1636943256
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1636943256
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1636943256
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_289
timestamp -25199
transform 1 0 27692 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_297
timestamp -25199
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_6
timestamp 1636943256
transform 1 0 1656 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_18
timestamp 1636943256
transform 1 0 2760 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_30
timestamp 1636943256
transform 1 0 3864 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_42
timestamp 1636943256
transform 1 0 4968 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp -25199
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1636943256
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1636943256
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1636943256
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1636943256
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp -25199
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp -25199
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1636943256
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_125
timestamp -25199
transform 1 0 12604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_129
timestamp -25199
transform 1 0 12972 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_151
timestamp 1636943256
transform 1 0 14996 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_163
timestamp -25199
transform 1 0 16100 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp -25199
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1636943256
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1636943256
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1636943256
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1636943256
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp -25199
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp -25199
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1636943256
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1636943256
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1636943256
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1636943256
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp -25199
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp -25199
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1636943256
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636943256
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636943256
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp -25199
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1636943256
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1636943256
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1636943256
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1636943256
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp -25199
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp -25199
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1636943256
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_97
timestamp -25199
transform 1 0 10028 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_105
timestamp -25199
transform 1 0 10764 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_129
timestamp -25199
transform 1 0 12972 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_137
timestamp -25199
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_150
timestamp 1636943256
transform 1 0 14904 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_162
timestamp 1636943256
transform 1 0 16008 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_174
timestamp 1636943256
transform 1 0 17112 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_186
timestamp -25199
transform 1 0 18216 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp -25199
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1636943256
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1636943256
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1636943256
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1636943256
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp -25199
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp -25199
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1636943256
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1636943256
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1636943256
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_289
timestamp -25199
transform 1 0 27692 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_6
timestamp 1636943256
transform 1 0 1656 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_18
timestamp 1636943256
transform 1 0 2760 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_30
timestamp 1636943256
transform 1 0 3864 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_42
timestamp 1636943256
transform 1 0 4968 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp -25199
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1636943256
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1636943256
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1636943256
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1636943256
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp -25199
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp -25199
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_126
timestamp -25199
transform 1 0 12696 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_151
timestamp 1636943256
transform 1 0 14996 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_163
timestamp -25199
transform 1 0 16100 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp -25199
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1636943256
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1636943256
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1636943256
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1636943256
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp -25199
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp -25199
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1636943256
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1636943256
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1636943256
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1636943256
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp -25199
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp -25199
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1636943256
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_293
timestamp -25199
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_6
timestamp 1636943256
transform 1 0 1656 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_18
timestamp -25199
transform 1 0 2760 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp -25199
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1636943256
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1636943256
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1636943256
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1636943256
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp -25199
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp -25199
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1636943256
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1636943256
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp -25199
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp -25199
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_150
timestamp 1636943256
transform 1 0 14904 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_162
timestamp 1636943256
transform 1 0 16008 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_174
timestamp 1636943256
transform 1 0 17112 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_186
timestamp -25199
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp -25199
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1636943256
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1636943256
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1636943256
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1636943256
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp -25199
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp -25199
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1636943256
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1636943256
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1636943256
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_289
timestamp -25199
transform 1 0 27692 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1636943256
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1636943256
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1636943256
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1636943256
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp -25199
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp -25199
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1636943256
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1636943256
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1636943256
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1636943256
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp -25199
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp -25199
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_122
timestamp 1636943256
transform 1 0 12328 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_134
timestamp 1636943256
transform 1 0 13432 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_146
timestamp 1636943256
transform 1 0 14536 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_158
timestamp -25199
transform 1 0 15640 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp -25199
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1636943256
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1636943256
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1636943256
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1636943256
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp -25199
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp -25199
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1636943256
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1636943256
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1636943256
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1636943256
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp -25199
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp -25199
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1636943256
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_6
timestamp 1636943256
transform 1 0 1656 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_18
timestamp -25199
transform 1 0 2760 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp -25199
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636943256
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1636943256
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1636943256
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1636943256
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp -25199
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp -25199
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1636943256
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_97
timestamp -25199
transform 1 0 10028 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_105
timestamp -25199
transform 1 0 10764 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp -25199
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1636943256
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1636943256
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1636943256
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1636943256
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp -25199
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp -25199
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1636943256
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1636943256
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1636943256
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1636943256
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp -25199
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp -25199
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1636943256
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1636943256
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1636943256
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_289
timestamp -25199
transform 1 0 27692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_297
timestamp -25199
transform 1 0 28428 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_6
timestamp 1636943256
transform 1 0 1656 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_18
timestamp 1636943256
transform 1 0 2760 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_30
timestamp 1636943256
transform 1 0 3864 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_42
timestamp 1636943256
transform 1 0 4968 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp -25199
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1636943256
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1636943256
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1636943256
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1636943256
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp -25199
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp -25199
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_113
timestamp -25199
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_140
timestamp 1636943256
transform 1 0 13984 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_152
timestamp 1636943256
transform 1 0 15088 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp -25199
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1636943256
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1636943256
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1636943256
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1636943256
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp -25199
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp -25199
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1636943256
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1636943256
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1636943256
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1636943256
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp -25199
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp -25199
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1636943256
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636943256
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1636943256
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp -25199
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636943256
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1636943256
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1636943256
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1636943256
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp -25199
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp -25199
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1636943256
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_97
timestamp -25199
transform 1 0 10028 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_105
timestamp -25199
transform 1 0 10764 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_129
timestamp -25199
transform 1 0 12972 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp -25199
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1636943256
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1636943256
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1636943256
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1636943256
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp -25199
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp -25199
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1636943256
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1636943256
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1636943256
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1636943256
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp -25199
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp -25199
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1636943256
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1636943256
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1636943256
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_289
timestamp -25199
transform 1 0 27692 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_6
timestamp 1636943256
transform 1 0 1656 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_18
timestamp 1636943256
transform 1 0 2760 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_30
timestamp 1636943256
transform 1 0 3864 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_42
timestamp 1636943256
transform 1 0 4968 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp -25199
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1636943256
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1636943256
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1636943256
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_93
timestamp -25199
transform 1 0 9660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_101
timestamp -25199
transform 1 0 10396 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp -25199
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_136
timestamp 1636943256
transform 1 0 13616 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_148
timestamp 1636943256
transform 1 0 14720 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_160
timestamp -25199
transform 1 0 15824 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1636943256
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1636943256
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1636943256
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1636943256
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp -25199
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp -25199
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1636943256
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1636943256
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1636943256
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1636943256
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp -25199
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp -25199
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1636943256
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_293
timestamp -25199
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_6
timestamp 1636943256
transform 1 0 1656 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_18
timestamp -25199
transform 1 0 2760 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp -25199
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1636943256
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1636943256
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1636943256
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1636943256
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp -25199
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp -25199
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp -25199
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp -25199
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1636943256
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1636943256
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1636943256
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1636943256
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp -25199
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp -25199
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1636943256
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1636943256
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1636943256
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1636943256
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp -25199
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp -25199
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1636943256
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1636943256
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1636943256
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_289
timestamp -25199
transform 1 0 27692 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1636943256
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1636943256
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1636943256
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1636943256
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp -25199
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp -25199
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1636943256
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1636943256
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1636943256
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_93
timestamp -25199
transform 1 0 9660 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_101
timestamp -25199
transform 1 0 10396 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1636943256
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1636943256
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1636943256
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp -25199
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp -25199
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1636943256
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1636943256
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1636943256
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1636943256
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp -25199
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp -25199
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1636943256
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1636943256
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1636943256
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1636943256
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp -25199
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp -25199
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1636943256
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_12
timestamp 1636943256
transform 1 0 2208 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp -25199
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1636943256
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1636943256
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_53
timestamp -25199
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_57
timestamp 1636943256
transform 1 0 6348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_69
timestamp 1636943256
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp -25199
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1636943256
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1636943256
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_109
timestamp -25199
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_116
timestamp 1636943256
transform 1 0 11776 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_128
timestamp 1636943256
transform 1 0 12880 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1636943256
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1636943256
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_165
timestamp -25199
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_169
timestamp 1636943256
transform 1 0 16652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_181
timestamp 1636943256
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_193
timestamp -25199
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1636943256
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1636943256
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_221
timestamp -25199
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_225
timestamp 1636943256
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_237
timestamp 1636943256
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp -25199
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1636943256
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1636943256
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_277
timestamp -25199
transform 1 0 26588 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_281
timestamp 1636943256
transform 1 0 26956 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp -25199
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp -25199
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp -25199
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp -25199
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp -25199
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp -25199
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp -25199
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp -25199
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp -25199
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp -25199
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp -25199
transform -1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp -25199
transform -1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp -25199
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp -25199
transform -1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp -25199
transform -1 0 1656 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp -25199
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp -25199
transform -1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp -25199
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp -25199
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp -25199
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp -25199
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp -25199
transform -1 0 1656 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp -25199
transform 1 0 1380 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp -25199
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp -25199
transform -1 0 1656 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp -25199
transform 1 0 1380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp -25199
transform -1 0 1656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp -25199
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp -25199
transform -1 0 1656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp -25199
transform 1 0 1380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp -25199
transform -1 0 1932 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp -25199
transform -1 0 2208 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp -25199
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp -25199
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  output35
timestamp -25199
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output36
timestamp -25199
transform 1 0 28060 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output37
timestamp -25199
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output38
timestamp -25199
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output39
timestamp -25199
transform 1 0 28060 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output40
timestamp -25199
transform 1 0 28060 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output41
timestamp -25199
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output42
timestamp -25199
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output43
timestamp -25199
transform 1 0 28060 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output44
timestamp -25199
transform 1 0 28060 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output45
timestamp -25199
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output46
timestamp -25199
transform 1 0 28060 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output47
timestamp -25199
transform 1 0 28060 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output48
timestamp -25199
transform 1 0 28060 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output49
timestamp -25199
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output50
timestamp -25199
transform 1 0 28060 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output51
timestamp -25199
transform 1 0 28060 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output52
timestamp -25199
transform 1 0 28060 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output53
timestamp -25199
transform 1 0 28060 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output54
timestamp -25199
transform 1 0 28060 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output55
timestamp -25199
transform 1 0 28060 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output56
timestamp -25199
transform 1 0 28060 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output57
timestamp -25199
transform 1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output58
timestamp -25199
transform 1 0 28060 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output59
timestamp -25199
transform 1 0 28060 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output60
timestamp -25199
transform 1 0 28060 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output61
timestamp -25199
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output62
timestamp -25199
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output63
timestamp -25199
transform 1 0 28060 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output64
timestamp -25199
transform 1 0 28060 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output65
timestamp -25199
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output66
timestamp -25199
transform 1 0 28060 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_47
timestamp -25199
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -25199
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_48
timestamp -25199
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -25199
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_49
timestamp -25199
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -25199
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_50
timestamp -25199
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -25199
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_51
timestamp -25199
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -25199
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_52
timestamp -25199
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -25199
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_53
timestamp -25199
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -25199
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_54
timestamp -25199
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -25199
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_55
timestamp -25199
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -25199
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_56
timestamp -25199
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -25199
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_57
timestamp -25199
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -25199
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_58
timestamp -25199
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -25199
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_59
timestamp -25199
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -25199
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_60
timestamp -25199
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -25199
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_61
timestamp -25199
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -25199
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_62
timestamp -25199
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -25199
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_63
timestamp -25199
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -25199
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_64
timestamp -25199
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -25199
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_65
timestamp -25199
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -25199
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_66
timestamp -25199
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -25199
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_67
timestamp -25199
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -25199
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_68
timestamp -25199
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -25199
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_69
timestamp -25199
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -25199
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_70
timestamp -25199
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -25199
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_71
timestamp -25199
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -25199
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_72
timestamp -25199
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp -25199
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_73
timestamp -25199
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp -25199
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_74
timestamp -25199
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp -25199
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_75
timestamp -25199
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp -25199
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_76
timestamp -25199
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp -25199
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_77
timestamp -25199
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp -25199
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_78
timestamp -25199
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp -25199
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_79
timestamp -25199
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp -25199
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_80
timestamp -25199
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp -25199
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_81
timestamp -25199
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp -25199
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_82
timestamp -25199
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp -25199
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_83
timestamp -25199
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp -25199
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_84
timestamp -25199
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp -25199
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_85
timestamp -25199
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp -25199
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_86
timestamp -25199
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp -25199
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_87
timestamp -25199
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp -25199
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_88
timestamp -25199
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp -25199
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_89
timestamp -25199
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp -25199
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_90
timestamp -25199
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp -25199
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_91
timestamp -25199
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp -25199
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_92
timestamp -25199
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp -25199
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_93
timestamp -25199
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp -25199
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_94
timestamp -25199
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_95
timestamp -25199
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_96
timestamp -25199
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_97
timestamp -25199
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_98
timestamp -25199
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_99
timestamp -25199
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_100
timestamp -25199
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_101
timestamp -25199
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_102
timestamp -25199
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_103
timestamp -25199
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_104
timestamp -25199
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_105
timestamp -25199
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_106
timestamp -25199
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_107
timestamp -25199
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_108
timestamp -25199
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_109
timestamp -25199
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_110
timestamp -25199
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_111
timestamp -25199
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_112
timestamp -25199
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_113
timestamp -25199
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_114
timestamp -25199
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_115
timestamp -25199
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_116
timestamp -25199
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_117
timestamp -25199
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_118
timestamp -25199
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_119
timestamp -25199
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_120
timestamp -25199
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_121
timestamp -25199
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_122
timestamp -25199
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_123
timestamp -25199
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_124
timestamp -25199
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_125
timestamp -25199
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_126
timestamp -25199
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_127
timestamp -25199
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_128
timestamp -25199
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_129
timestamp -25199
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_130
timestamp -25199
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_131
timestamp -25199
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_132
timestamp -25199
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_133
timestamp -25199
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_134
timestamp -25199
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_135
timestamp -25199
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_136
timestamp -25199
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_137
timestamp -25199
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_138
timestamp -25199
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_139
timestamp -25199
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_140
timestamp -25199
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_141
timestamp -25199
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_142
timestamp -25199
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_143
timestamp -25199
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_144
timestamp -25199
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_145
timestamp -25199
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_146
timestamp -25199
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_147
timestamp -25199
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_148
timestamp -25199
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_149
timestamp -25199
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_150
timestamp -25199
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_151
timestamp -25199
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_152
timestamp -25199
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_153
timestamp -25199
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_154
timestamp -25199
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_155
timestamp -25199
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_156
timestamp -25199
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_157
timestamp -25199
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_158
timestamp -25199
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_159
timestamp -25199
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_160
timestamp -25199
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_161
timestamp -25199
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_162
timestamp -25199
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_163
timestamp -25199
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_164
timestamp -25199
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_165
timestamp -25199
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_166
timestamp -25199
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_167
timestamp -25199
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_168
timestamp -25199
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_169
timestamp -25199
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_170
timestamp -25199
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_171
timestamp -25199
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_172
timestamp -25199
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_173
timestamp -25199
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_174
timestamp -25199
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_175
timestamp -25199
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_176
timestamp -25199
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_177
timestamp -25199
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_178
timestamp -25199
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_179
timestamp -25199
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_180
timestamp -25199
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_181
timestamp -25199
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_182
timestamp -25199
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_183
timestamp -25199
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_184
timestamp -25199
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_185
timestamp -25199
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_186
timestamp -25199
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_187
timestamp -25199
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_188
timestamp -25199
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_189
timestamp -25199
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_190
timestamp -25199
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_191
timestamp -25199
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_192
timestamp -25199
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_193
timestamp -25199
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_194
timestamp -25199
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_195
timestamp -25199
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_196
timestamp -25199
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_197
timestamp -25199
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_198
timestamp -25199
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_199
timestamp -25199
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_200
timestamp -25199
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_201
timestamp -25199
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_202
timestamp -25199
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_203
timestamp -25199
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_204
timestamp -25199
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_205
timestamp -25199
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_206
timestamp -25199
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_207
timestamp -25199
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_208
timestamp -25199
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_209
timestamp -25199
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_210
timestamp -25199
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_211
timestamp -25199
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_212
timestamp -25199
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_213
timestamp -25199
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_214
timestamp -25199
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_215
timestamp -25199
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_216
timestamp -25199
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_217
timestamp -25199
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_218
timestamp -25199
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_219
timestamp -25199
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_220
timestamp -25199
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_221
timestamp -25199
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_222
timestamp -25199
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_223
timestamp -25199
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_224
timestamp -25199
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_225
timestamp -25199
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_226
timestamp -25199
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_227
timestamp -25199
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_228
timestamp -25199
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_229
timestamp -25199
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_230
timestamp -25199
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_231
timestamp -25199
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_232
timestamp -25199
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_233
timestamp -25199
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_234
timestamp -25199
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_235
timestamp -25199
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_236
timestamp -25199
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_237
timestamp -25199
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_238
timestamp -25199
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_239
timestamp -25199
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_240
timestamp -25199
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_241
timestamp -25199
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_242
timestamp -25199
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_243
timestamp -25199
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_244
timestamp -25199
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_245
timestamp -25199
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_246
timestamp -25199
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_247
timestamp -25199
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_248
timestamp -25199
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_249
timestamp -25199
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_250
timestamp -25199
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_251
timestamp -25199
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_252
timestamp -25199
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp -25199
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_254
timestamp -25199
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_255
timestamp -25199
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_256
timestamp -25199
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_257
timestamp -25199
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp -25199
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_259
timestamp -25199
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_260
timestamp -25199
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_261
timestamp -25199
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_262
timestamp -25199
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp -25199
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_264
timestamp -25199
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp -25199
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_266
timestamp -25199
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_267
timestamp -25199
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp -25199
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_269
timestamp -25199
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_270
timestamp -25199
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_271
timestamp -25199
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_272
timestamp -25199
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp -25199
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_274
timestamp -25199
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_275
timestamp -25199
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_276
timestamp -25199
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_277
timestamp -25199
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp -25199
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_279
timestamp -25199
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_280
timestamp -25199
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_281
timestamp -25199
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_282
timestamp -25199
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp -25199
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_284
timestamp -25199
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_285
timestamp -25199
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_286
timestamp -25199
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_287
timestamp -25199
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp -25199
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_289
timestamp -25199
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_290
timestamp -25199
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_291
timestamp -25199
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_292
timestamp -25199
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp -25199
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_294
timestamp -25199
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_295
timestamp -25199
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_296
timestamp -25199
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_297
timestamp -25199
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_298
timestamp -25199
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_299
timestamp -25199
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_300
timestamp -25199
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_301
timestamp -25199
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_302
timestamp -25199
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_303
timestamp -25199
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_304
timestamp -25199
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_305
timestamp -25199
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_306
timestamp -25199
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_307
timestamp -25199
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_308
timestamp -25199
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_309
timestamp -25199
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_310
timestamp -25199
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_311
timestamp -25199
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_312
timestamp -25199
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_313
timestamp -25199
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_314
timestamp -25199
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_315
timestamp -25199
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_316
timestamp -25199
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_317
timestamp -25199
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_318
timestamp -25199
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_319
timestamp -25199
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_320
timestamp -25199
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_321
timestamp -25199
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_322
timestamp -25199
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_323
timestamp -25199
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_324
timestamp -25199
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_325
timestamp -25199
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_326
timestamp -25199
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_327
timestamp -25199
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_328
timestamp -25199
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_329
timestamp -25199
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_330
timestamp -25199
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_331
timestamp -25199
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_332
timestamp -25199
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_333
timestamp -25199
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_334
timestamp -25199
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_335
timestamp -25199
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_336
timestamp -25199
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_337
timestamp -25199
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_338
timestamp -25199
transform 1 0 26864 0 1 27200
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 824 800 944 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 29200 2184 30000 2304 0 FreeSans 480 0 0 0 pm_current_s0_o[0]
port 1 nsew signal output
flabel metal3 s 29200 3000 30000 3120 0 FreeSans 480 0 0 0 pm_current_s0_o[1]
port 2 nsew signal output
flabel metal3 s 29200 3816 30000 3936 0 FreeSans 480 0 0 0 pm_current_s0_o[2]
port 3 nsew signal output
flabel metal3 s 29200 4632 30000 4752 0 FreeSans 480 0 0 0 pm_current_s0_o[3]
port 4 nsew signal output
flabel metal3 s 29200 5448 30000 5568 0 FreeSans 480 0 0 0 pm_current_s0_o[4]
port 5 nsew signal output
flabel metal3 s 29200 6264 30000 6384 0 FreeSans 480 0 0 0 pm_current_s0_o[5]
port 6 nsew signal output
flabel metal3 s 29200 7080 30000 7200 0 FreeSans 480 0 0 0 pm_current_s0_o[6]
port 7 nsew signal output
flabel metal3 s 29200 7896 30000 8016 0 FreeSans 480 0 0 0 pm_current_s0_o[7]
port 8 nsew signal output
flabel metal3 s 29200 8712 30000 8832 0 FreeSans 480 0 0 0 pm_current_s1_o[0]
port 9 nsew signal output
flabel metal3 s 29200 9528 30000 9648 0 FreeSans 480 0 0 0 pm_current_s1_o[1]
port 10 nsew signal output
flabel metal3 s 29200 10344 30000 10464 0 FreeSans 480 0 0 0 pm_current_s1_o[2]
port 11 nsew signal output
flabel metal3 s 29200 11160 30000 11280 0 FreeSans 480 0 0 0 pm_current_s1_o[3]
port 12 nsew signal output
flabel metal3 s 29200 11976 30000 12096 0 FreeSans 480 0 0 0 pm_current_s1_o[4]
port 13 nsew signal output
flabel metal3 s 29200 12792 30000 12912 0 FreeSans 480 0 0 0 pm_current_s1_o[5]
port 14 nsew signal output
flabel metal3 s 29200 13608 30000 13728 0 FreeSans 480 0 0 0 pm_current_s1_o[6]
port 15 nsew signal output
flabel metal3 s 29200 14424 30000 14544 0 FreeSans 480 0 0 0 pm_current_s1_o[7]
port 16 nsew signal output
flabel metal3 s 29200 15240 30000 15360 0 FreeSans 480 0 0 0 pm_current_s2_o[0]
port 17 nsew signal output
flabel metal3 s 29200 16056 30000 16176 0 FreeSans 480 0 0 0 pm_current_s2_o[1]
port 18 nsew signal output
flabel metal3 s 29200 16872 30000 16992 0 FreeSans 480 0 0 0 pm_current_s2_o[2]
port 19 nsew signal output
flabel metal3 s 29200 17688 30000 17808 0 FreeSans 480 0 0 0 pm_current_s2_o[3]
port 20 nsew signal output
flabel metal3 s 29200 18504 30000 18624 0 FreeSans 480 0 0 0 pm_current_s2_o[4]
port 21 nsew signal output
flabel metal3 s 29200 19320 30000 19440 0 FreeSans 480 0 0 0 pm_current_s2_o[5]
port 22 nsew signal output
flabel metal3 s 29200 20136 30000 20256 0 FreeSans 480 0 0 0 pm_current_s2_o[6]
port 23 nsew signal output
flabel metal3 s 29200 20952 30000 21072 0 FreeSans 480 0 0 0 pm_current_s2_o[7]
port 24 nsew signal output
flabel metal3 s 29200 21768 30000 21888 0 FreeSans 480 0 0 0 pm_current_s3_o[0]
port 25 nsew signal output
flabel metal3 s 29200 22584 30000 22704 0 FreeSans 480 0 0 0 pm_current_s3_o[1]
port 26 nsew signal output
flabel metal3 s 29200 23400 30000 23520 0 FreeSans 480 0 0 0 pm_current_s3_o[2]
port 27 nsew signal output
flabel metal3 s 29200 24216 30000 24336 0 FreeSans 480 0 0 0 pm_current_s3_o[3]
port 28 nsew signal output
flabel metal3 s 29200 25032 30000 25152 0 FreeSans 480 0 0 0 pm_current_s3_o[4]
port 29 nsew signal output
flabel metal3 s 29200 25848 30000 25968 0 FreeSans 480 0 0 0 pm_current_s3_o[5]
port 30 nsew signal output
flabel metal3 s 29200 26664 30000 26784 0 FreeSans 480 0 0 0 pm_current_s3_o[6]
port 31 nsew signal output
flabel metal3 s 29200 27480 30000 27600 0 FreeSans 480 0 0 0 pm_current_s3_o[7]
port 32 nsew signal output
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 pm_new_s0_i[0]
port 33 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 pm_new_s0_i[1]
port 34 nsew signal input
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 pm_new_s0_i[2]
port 35 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 pm_new_s0_i[3]
port 36 nsew signal input
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 pm_new_s0_i[4]
port 37 nsew signal input
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 pm_new_s0_i[5]
port 38 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 pm_new_s0_i[6]
port 39 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 pm_new_s0_i[7]
port 40 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 pm_new_s1_i[0]
port 41 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 pm_new_s1_i[1]
port 42 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 pm_new_s1_i[2]
port 43 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 pm_new_s1_i[3]
port 44 nsew signal input
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 pm_new_s1_i[4]
port 45 nsew signal input
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 pm_new_s1_i[5]
port 46 nsew signal input
flabel metal3 s 0 14696 800 14816 0 FreeSans 480 0 0 0 pm_new_s1_i[6]
port 47 nsew signal input
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 pm_new_s1_i[7]
port 48 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 pm_new_s2_i[0]
port 49 nsew signal input
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 pm_new_s2_i[1]
port 50 nsew signal input
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 pm_new_s2_i[2]
port 51 nsew signal input
flabel metal3 s 0 18776 800 18896 0 FreeSans 480 0 0 0 pm_new_s2_i[3]
port 52 nsew signal input
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 pm_new_s2_i[4]
port 53 nsew signal input
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 pm_new_s2_i[5]
port 54 nsew signal input
flabel metal3 s 0 21224 800 21344 0 FreeSans 480 0 0 0 pm_new_s2_i[6]
port 55 nsew signal input
flabel metal3 s 0 22040 800 22160 0 FreeSans 480 0 0 0 pm_new_s2_i[7]
port 56 nsew signal input
flabel metal3 s 0 22856 800 22976 0 FreeSans 480 0 0 0 pm_new_s3_i[0]
port 57 nsew signal input
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 pm_new_s3_i[1]
port 58 nsew signal input
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 pm_new_s3_i[2]
port 59 nsew signal input
flabel metal3 s 0 25304 800 25424 0 FreeSans 480 0 0 0 pm_new_s3_i[3]
port 60 nsew signal input
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 pm_new_s3_i[4]
port 61 nsew signal input
flabel metal3 s 0 26936 800 27056 0 FreeSans 480 0 0 0 pm_new_s3_i[5]
port 62 nsew signal input
flabel metal3 s 0 27752 800 27872 0 FreeSans 480 0 0 0 pm_new_s3_i[6]
port 63 nsew signal input
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 pm_new_s3_i[7]
port 64 nsew signal input
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 rst_n
port 65 nsew signal input
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 valid_i
port 66 nsew signal input
flabel metal4 s 2904 2128 3304 27792 0 FreeSans 1920 90 0 0 vccd1
port 67 nsew power bidirectional
flabel metal4 s 10904 2128 11304 27792 0 FreeSans 1920 90 0 0 vccd1
port 67 nsew power bidirectional
flabel metal4 s 18904 2128 19304 27792 0 FreeSans 1920 90 0 0 vccd1
port 67 nsew power bidirectional
flabel metal4 s 26904 2128 27304 27792 0 FreeSans 1920 90 0 0 vccd1
port 67 nsew power bidirectional
flabel metal4 s 3644 2128 4044 27792 0 FreeSans 1920 90 0 0 vssd1
port 68 nsew ground bidirectional
flabel metal4 s 11644 2128 12044 27792 0 FreeSans 1920 90 0 0 vssd1
port 68 nsew ground bidirectional
flabel metal4 s 19644 2128 20044 27792 0 FreeSans 1920 90 0 0 vssd1
port 68 nsew ground bidirectional
flabel metal4 s 27644 2128 28044 27792 0 FreeSans 1920 90 0 0 vssd1
port 68 nsew ground bidirectional
rlabel metal1 14996 27744 14996 27744 0 vccd1
rlabel metal1 14996 27200 14996 27200 0 vssd1
rlabel metal1 11592 2958 11592 2958 0 _00_
rlabel metal1 11914 3638 11914 3638 0 _01_
rlabel metal2 12466 4250 12466 4250 0 _02_
rlabel metal1 11224 4658 11224 4658 0 _03_
rlabel metal1 10902 5746 10902 5746 0 _04_
rlabel metal1 11592 6222 11592 6222 0 _05_
rlabel metal1 11270 7514 11270 7514 0 _06_
rlabel metal1 11730 8398 11730 8398 0 _07_
rlabel metal1 11638 9486 11638 9486 0 _08_
rlabel metal1 12650 10132 12650 10132 0 _09_
rlabel metal1 11316 10778 11316 10778 0 _10_
rlabel metal1 11454 10506 11454 10506 0 _11_
rlabel metal1 11224 12274 11224 12274 0 _12_
rlabel metal1 12282 12750 12282 12750 0 _13_
rlabel metal1 11270 13362 11270 13362 0 _14_
rlabel metal1 10902 14450 10902 14450 0 _15_
rlabel metal2 11454 22202 11454 22202 0 _16_
rlabel metal2 13478 22780 13478 22780 0 _17_
rlabel metal2 11546 24004 11546 24004 0 _18_
rlabel metal2 13018 24548 13018 24548 0 _19_
rlabel metal2 11454 25500 11454 25500 0 _20_
rlabel metal2 13018 26010 13018 26010 0 _21_
rlabel metal2 11454 26588 11454 26588 0 _22_
rlabel metal2 10626 26588 10626 26588 0 _23_
rlabel metal1 11638 16014 11638 16014 0 _24_
rlabel metal2 12098 16116 12098 16116 0 _25_
rlabel metal2 12466 17340 12466 17340 0 _26_
rlabel metal2 12742 18428 12742 18428 0 _27_
rlabel metal2 13018 19516 13018 19516 0 _28_
rlabel metal1 11500 19482 11500 19482 0 _29_
rlabel metal1 13708 20366 13708 20366 0 _30_
rlabel metal2 13478 21692 13478 21692 0 _31_
rlabel metal1 6900 14994 6900 14994 0 clk
rlabel metal1 11868 17646 11868 17646 0 clknet_0_clk
rlabel metal1 11546 12716 11546 12716 0 clknet_2_0__leaf_clk
rlabel metal2 10718 8092 10718 8092 0 clknet_2_1__leaf_clk
rlabel metal2 13110 22032 13110 22032 0 clknet_2_2__leaf_clk
rlabel metal1 11822 17102 11822 17102 0 clknet_2_3__leaf_clk
rlabel metal1 10580 3162 10580 3162 0 net1
rlabel metal1 2185 11254 2185 11254 0 net10
rlabel metal1 12052 10778 12052 10778 0 net11
rlabel metal1 6118 12614 6118 12614 0 net12
rlabel metal2 10902 13056 10902 13056 0 net13
rlabel metal1 12604 13362 12604 13362 0 net14
rlabel metal1 11776 14042 11776 14042 0 net15
rlabel metal1 10948 15130 10948 15130 0 net16
rlabel metal2 10902 16320 10902 16320 0 net17
rlabel metal1 11960 15538 11960 15538 0 net18
rlabel metal2 14582 18054 14582 18054 0 net19
rlabel metal1 12834 3570 12834 3570 0 net2
rlabel metal2 14582 19006 14582 19006 0 net20
rlabel metal1 13662 19958 13662 19958 0 net21
rlabel metal1 11684 19414 11684 19414 0 net22
rlabel metal2 14582 21148 14582 21148 0 net23
rlabel metal1 14582 22134 14582 22134 0 net24
rlabel metal1 11592 22746 11592 22746 0 net25
rlabel metal2 14582 23426 14582 23426 0 net26
rlabel metal1 11730 23766 11730 23766 0 net27
rlabel metal1 12052 24242 12052 24242 0 net28
rlabel metal1 10672 26010 10672 26010 0 net29
rlabel metal1 12926 4726 12926 4726 0 net3
rlabel metal1 13386 26214 13386 26214 0 net30
rlabel metal1 11730 27098 11730 27098 0 net31
rlabel metal1 11040 27098 11040 27098 0 net32
rlabel metal1 13478 3400 13478 3400 0 net33
rlabel metal1 11362 4182 11362 4182 0 net34
rlabel metal2 20654 2618 20654 2618 0 net35
rlabel metal1 20470 3502 20470 3502 0 net36
rlabel metal1 13294 4080 13294 4080 0 net37
rlabel metal2 12558 4386 12558 4386 0 net38
rlabel metal1 12466 5712 12466 5712 0 net39
rlabel metal1 2185 6086 2185 6086 0 net4
rlabel metal2 28106 6426 28106 6426 0 net40
rlabel metal2 12466 7616 12466 7616 0 net41
rlabel metal1 13294 8432 13294 8432 0 net42
rlabel metal2 28106 9146 28106 9146 0 net43
rlabel metal1 12765 10030 12765 10030 0 net44
rlabel via1 12489 11050 12489 11050 0 net45
rlabel metal1 12926 11628 12926 11628 0 net46
rlabel metal1 11500 12818 11500 12818 0 net47
rlabel via1 13363 12954 13363 12954 0 net48
rlabel via1 12397 13498 12397 13498 0 net49
rlabel metal2 10074 6528 10074 6528 0 net5
rlabel metal1 14490 14382 14490 14382 0 net50
rlabel metal1 11132 16082 11132 16082 0 net51
rlabel metal2 21390 15980 21390 15980 0 net52
rlabel metal2 14490 17340 14490 17340 0 net53
rlabel metal2 14490 18428 14490 18428 0 net54
rlabel metal2 23506 19040 23506 19040 0 net55
rlabel metal1 12098 19482 12098 19482 0 net56
rlabel metal1 14582 20842 14582 20842 0 net57
rlabel metal2 17894 21726 17894 21726 0 net58
rlabel metal1 13547 21930 13547 21930 0 net59
rlabel metal1 10534 6426 10534 6426 0 net6
rlabel via1 14927 22746 14927 22746 0 net60
rlabel metal1 12282 23834 12282 23834 0 net61
rlabel metal2 13386 24480 13386 24480 0 net62
rlabel metal1 11316 25874 11316 25874 0 net63
rlabel via1 13547 26010 13547 26010 0 net64
rlabel metal2 21390 26656 21390 26656 0 net65
rlabel metal2 21298 27132 21298 27132 0 net66
rlabel metal2 13018 4896 13018 4896 0 net67
rlabel metal2 10810 13124 10810 13124 0 net68
rlabel metal1 11132 8398 11132 8398 0 net69
rlabel metal1 2185 8330 2185 8330 0 net7
rlabel metal1 14260 18802 14260 18802 0 net70
rlabel metal2 12098 24650 12098 24650 0 net71
rlabel metal2 12190 26656 12190 26656 0 net72
rlabel metal1 11776 19278 11776 19278 0 net73
rlabel metal1 12098 2618 12098 2618 0 net74
rlabel metal2 12466 12529 12466 12529 0 net75
rlabel metal1 12190 2414 12190 2414 0 net76
rlabel metal2 13754 18870 13754 18870 0 net77
rlabel via1 13846 22661 13846 22661 0 net78
rlabel metal1 12236 26010 12236 26010 0 net79
rlabel metal1 10856 8602 10856 8602 0 net8
rlabel metal2 12466 21182 12466 21182 0 net80
rlabel metal2 1610 9792 1610 9792 0 net9
rlabel metal2 28382 2295 28382 2295 0 pm_current_s0_o[0]
rlabel metal2 28382 3247 28382 3247 0 pm_current_s0_o[1]
rlabel metal2 28382 3961 28382 3961 0 pm_current_s0_o[2]
rlabel metal2 28382 4913 28382 4913 0 pm_current_s0_o[3]
rlabel metal2 28382 5559 28382 5559 0 pm_current_s0_o[4]
rlabel metal2 28382 6511 28382 6511 0 pm_current_s0_o[5]
rlabel metal2 28382 7225 28382 7225 0 pm_current_s0_o[6]
rlabel metal2 28382 8177 28382 8177 0 pm_current_s0_o[7]
rlabel metal2 28382 8823 28382 8823 0 pm_current_s1_o[0]
rlabel metal2 28382 9775 28382 9775 0 pm_current_s1_o[1]
rlabel metal2 28382 10489 28382 10489 0 pm_current_s1_o[2]
rlabel metal2 28382 11441 28382 11441 0 pm_current_s1_o[3]
rlabel metal2 28382 12087 28382 12087 0 pm_current_s1_o[4]
rlabel metal2 28382 13039 28382 13039 0 pm_current_s1_o[5]
rlabel metal2 28382 13753 28382 13753 0 pm_current_s1_o[6]
rlabel metal2 28382 14705 28382 14705 0 pm_current_s1_o[7]
rlabel metal2 28382 15351 28382 15351 0 pm_current_s2_o[0]
rlabel metal2 28382 16303 28382 16303 0 pm_current_s2_o[1]
rlabel metal2 28382 17017 28382 17017 0 pm_current_s2_o[2]
rlabel metal2 28382 17969 28382 17969 0 pm_current_s2_o[3]
rlabel metal2 28382 18615 28382 18615 0 pm_current_s2_o[4]
rlabel metal2 28382 19567 28382 19567 0 pm_current_s2_o[5]
rlabel metal2 28382 20281 28382 20281 0 pm_current_s2_o[6]
rlabel metal2 28382 21233 28382 21233 0 pm_current_s2_o[7]
rlabel metal2 28382 21879 28382 21879 0 pm_current_s3_o[0]
rlabel metal2 28382 22831 28382 22831 0 pm_current_s3_o[1]
rlabel metal2 28382 23545 28382 23545 0 pm_current_s3_o[2]
rlabel metal2 28382 24497 28382 24497 0 pm_current_s3_o[3]
rlabel metal2 28382 25143 28382 25143 0 pm_current_s3_o[4]
rlabel metal3 28850 25908 28850 25908 0 pm_current_s3_o[5]
rlabel metal2 28382 26809 28382 26809 0 pm_current_s3_o[6]
rlabel via2 28382 27523 28382 27523 0 pm_current_s3_o[7]
rlabel metal3 751 3332 751 3332 0 pm_new_s0_i[0]
rlabel metal3 751 4148 751 4148 0 pm_new_s0_i[1]
rlabel metal3 751 4964 751 4964 0 pm_new_s0_i[2]
rlabel metal3 751 5780 751 5780 0 pm_new_s0_i[3]
rlabel metal3 751 6596 751 6596 0 pm_new_s0_i[4]
rlabel metal3 751 7412 751 7412 0 pm_new_s0_i[5]
rlabel metal3 751 8228 751 8228 0 pm_new_s0_i[6]
rlabel metal3 751 9044 751 9044 0 pm_new_s0_i[7]
rlabel metal3 1050 9860 1050 9860 0 pm_new_s1_i[0]
rlabel metal3 751 10676 751 10676 0 pm_new_s1_i[1]
rlabel metal3 751 11492 751 11492 0 pm_new_s1_i[2]
rlabel metal3 751 12308 751 12308 0 pm_new_s1_i[3]
rlabel metal3 751 13124 751 13124 0 pm_new_s1_i[4]
rlabel metal3 751 13940 751 13940 0 pm_new_s1_i[5]
rlabel metal3 751 14756 751 14756 0 pm_new_s1_i[6]
rlabel metal3 751 15572 751 15572 0 pm_new_s1_i[7]
rlabel metal3 751 16388 751 16388 0 pm_new_s2_i[0]
rlabel metal3 751 17204 751 17204 0 pm_new_s2_i[1]
rlabel metal3 1050 18020 1050 18020 0 pm_new_s2_i[2]
rlabel metal1 1150 19346 1150 19346 0 pm_new_s2_i[3]
rlabel metal3 751 19652 751 19652 0 pm_new_s2_i[4]
rlabel metal3 751 20468 751 20468 0 pm_new_s2_i[5]
rlabel metal3 751 21284 751 21284 0 pm_new_s2_i[6]
rlabel metal3 751 22100 751 22100 0 pm_new_s2_i[7]
rlabel metal3 751 22916 751 22916 0 pm_new_s3_i[0]
rlabel metal3 751 23732 751 23732 0 pm_new_s3_i[1]
rlabel metal3 751 24548 751 24548 0 pm_new_s3_i[2]
rlabel metal3 751 25364 751 25364 0 pm_new_s3_i[3]
rlabel metal3 751 26180 751 26180 0 pm_new_s3_i[4]
rlabel metal3 751 26996 751 26996 0 pm_new_s3_i[5]
rlabel metal3 820 27812 820 27812 0 pm_new_s3_i[6]
rlabel metal3 866 28628 866 28628 0 pm_new_s3_i[7]
rlabel metal3 751 1700 751 1700 0 rst_n
rlabel metal3 751 2516 751 2516 0 valid_i
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
