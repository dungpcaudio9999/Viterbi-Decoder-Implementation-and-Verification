VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sync_fifo
  CLASS BLOCK ;
  FOREIGN sync_fifo ;
  ORIGIN 0.000 0.000 ;
  SIZE 182.365 BY 193.085 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END clk
  PIN empty_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 24.520 182.365 25.120 ;
    END
  END empty_o
  PIN full_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 15.000 182.365 15.600 ;
    END
  END full_o
  PIN rd_data_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 34.040 182.365 34.640 ;
    END
  END rd_data_o[0]
  PIN rd_data_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 129.240 182.365 129.840 ;
    END
  END rd_data_o[10]
  PIN rd_data_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 138.760 182.365 139.360 ;
    END
  END rd_data_o[11]
  PIN rd_data_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 148.280 182.365 148.880 ;
    END
  END rd_data_o[12]
  PIN rd_data_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 157.800 182.365 158.400 ;
    END
  END rd_data_o[13]
  PIN rd_data_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 167.320 182.365 167.920 ;
    END
  END rd_data_o[14]
  PIN rd_data_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 176.840 182.365 177.440 ;
    END
  END rd_data_o[15]
  PIN rd_data_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 43.560 182.365 44.160 ;
    END
  END rd_data_o[1]
  PIN rd_data_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 53.080 182.365 53.680 ;
    END
  END rd_data_o[2]
  PIN rd_data_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 62.600 182.365 63.200 ;
    END
  END rd_data_o[3]
  PIN rd_data_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 72.120 182.365 72.720 ;
    END
  END rd_data_o[4]
  PIN rd_data_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 81.640 182.365 82.240 ;
    END
  END rd_data_o[5]
  PIN rd_data_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 91.160 182.365 91.760 ;
    END
  END rd_data_o[6]
  PIN rd_data_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 100.680 182.365 101.280 ;
    END
  END rd_data_o[7]
  PIN rd_data_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 110.200 182.365 110.800 ;
    END
  END rd_data_o[8]
  PIN rd_data_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 178.365 119.720 182.365 120.320 ;
    END
  END rd_data_o[9]
  PIN rd_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END rd_en_i
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END rst_n
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 179.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 179.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 179.760 ;
    END
  END vssd1
  PIN wr_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END wr_data_i[0]
  PIN wr_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END wr_data_i[10]
  PIN wr_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END wr_data_i[11]
  PIN wr_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END wr_data_i[12]
  PIN wr_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END wr_data_i[13]
  PIN wr_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END wr_data_i[14]
  PIN wr_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END wr_data_i[15]
  PIN wr_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END wr_data_i[1]
  PIN wr_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END wr_data_i[2]
  PIN wr_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END wr_data_i[3]
  PIN wr_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END wr_data_i[4]
  PIN wr_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END wr_data_i[5]
  PIN wr_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END wr_data_i[6]
  PIN wr_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END wr_data_i[7]
  PIN wr_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END wr_data_i[8]
  PIN wr_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END wr_data_i[9]
  PIN wr_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END wr_en_i
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 176.830 179.605 ;
      LAYER li1 ;
        RECT 5.520 10.795 176.640 179.605 ;
      LAYER met1 ;
        RECT 5.520 10.640 177.030 179.760 ;
      LAYER met2 ;
        RECT 6.070 5.595 177.010 186.845 ;
      LAYER met3 ;
        RECT 4.400 185.960 178.365 186.825 ;
        RECT 4.000 177.840 178.365 185.960 ;
        RECT 4.400 176.440 177.965 177.840 ;
        RECT 4.000 168.320 178.365 176.440 ;
        RECT 4.400 166.920 177.965 168.320 ;
        RECT 4.000 158.800 178.365 166.920 ;
        RECT 4.400 157.400 177.965 158.800 ;
        RECT 4.000 149.280 178.365 157.400 ;
        RECT 4.400 147.880 177.965 149.280 ;
        RECT 4.000 139.760 178.365 147.880 ;
        RECT 4.400 138.360 177.965 139.760 ;
        RECT 4.000 130.240 178.365 138.360 ;
        RECT 4.400 128.840 177.965 130.240 ;
        RECT 4.000 120.720 178.365 128.840 ;
        RECT 4.400 119.320 177.965 120.720 ;
        RECT 4.000 111.200 178.365 119.320 ;
        RECT 4.400 109.800 177.965 111.200 ;
        RECT 4.000 101.680 178.365 109.800 ;
        RECT 4.400 100.280 177.965 101.680 ;
        RECT 4.000 92.160 178.365 100.280 ;
        RECT 4.400 90.760 177.965 92.160 ;
        RECT 4.000 82.640 178.365 90.760 ;
        RECT 4.400 81.240 177.965 82.640 ;
        RECT 4.000 73.120 178.365 81.240 ;
        RECT 4.400 71.720 177.965 73.120 ;
        RECT 4.000 63.600 178.365 71.720 ;
        RECT 4.400 62.200 177.965 63.600 ;
        RECT 4.000 54.080 178.365 62.200 ;
        RECT 4.400 52.680 177.965 54.080 ;
        RECT 4.000 44.560 178.365 52.680 ;
        RECT 4.400 43.160 177.965 44.560 ;
        RECT 4.000 35.040 178.365 43.160 ;
        RECT 4.400 33.640 177.965 35.040 ;
        RECT 4.000 25.520 178.365 33.640 ;
        RECT 4.400 24.120 177.965 25.520 ;
        RECT 4.000 16.000 178.365 24.120 ;
        RECT 4.400 14.600 177.965 16.000 ;
        RECT 4.000 6.480 178.365 14.600 ;
        RECT 4.400 5.615 178.365 6.480 ;
      LAYER met4 ;
        RECT 75.735 34.175 153.345 177.305 ;
  END
END sync_fifo
END LIBRARY

