VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tbu
  CLASS BLOCK ;
  FOREIGN tbu ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 150.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END clk
  PIN dec_bits_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END dec_bits_i[0]
  PIN dec_bits_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END dec_bits_i[1]
  PIN dec_bits_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END dec_bits_i[2]
  PIN dec_bits_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END dec_bits_i[3]
  PIN decoded_bit_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 36.760 150.000 37.360 ;
    END
  END decoded_bit_o
  PIN pm_new_s0_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END pm_new_s0_i[0]
  PIN pm_new_s0_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END pm_new_s0_i[1]
  PIN pm_new_s0_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END pm_new_s0_i[2]
  PIN pm_new_s0_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END pm_new_s0_i[3]
  PIN pm_new_s0_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END pm_new_s0_i[4]
  PIN pm_new_s0_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END pm_new_s0_i[5]
  PIN pm_new_s0_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END pm_new_s0_i[6]
  PIN pm_new_s0_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END pm_new_s0_i[7]
  PIN pm_new_s1_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END pm_new_s1_i[0]
  PIN pm_new_s1_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END pm_new_s1_i[1]
  PIN pm_new_s1_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END pm_new_s1_i[2]
  PIN pm_new_s1_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END pm_new_s1_i[3]
  PIN pm_new_s1_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END pm_new_s1_i[4]
  PIN pm_new_s1_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END pm_new_s1_i[5]
  PIN pm_new_s1_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END pm_new_s1_i[6]
  PIN pm_new_s1_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END pm_new_s1_i[7]
  PIN pm_new_s2_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END pm_new_s2_i[0]
  PIN pm_new_s2_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END pm_new_s2_i[1]
  PIN pm_new_s2_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END pm_new_s2_i[2]
  PIN pm_new_s2_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END pm_new_s2_i[3]
  PIN pm_new_s2_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END pm_new_s2_i[4]
  PIN pm_new_s2_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END pm_new_s2_i[5]
  PIN pm_new_s2_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END pm_new_s2_i[6]
  PIN pm_new_s2_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END pm_new_s2_i[7]
  PIN pm_new_s3_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END pm_new_s3_i[0]
  PIN pm_new_s3_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END pm_new_s3_i[1]
  PIN pm_new_s3_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END pm_new_s3_i[2]
  PIN pm_new_s3_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END pm_new_s3_i[3]
  PIN pm_new_s3_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END pm_new_s3_i[4]
  PIN pm_new_s3_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END pm_new_s3_i[5]
  PIN pm_new_s3_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END pm_new_s3_i[6]
  PIN pm_new_s3_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END pm_new_s3_i[7]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END rst_n
  PIN valid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END valid_i
  PIN valid_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 146.000 111.560 150.000 112.160 ;
    END
  END valid_o
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.520 10.640 16.520 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.520 10.640 56.520 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.520 10.640 96.520 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.520 10.640 136.520 138.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 18.220 10.640 20.220 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.220 10.640 60.220 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.220 10.640 100.220 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.220 10.640 140.220 138.960 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 144.630 138.910 ;
      LAYER li1 ;
        RECT 5.520 10.795 144.440 138.805 ;
      LAYER met1 ;
        RECT 5.130 10.640 144.440 138.960 ;
      LAYER met2 ;
        RECT 5.150 10.695 142.050 138.905 ;
      LAYER met3 ;
        RECT 4.000 126.160 146.000 138.885 ;
        RECT 4.400 124.760 146.000 126.160 ;
        RECT 4.000 123.440 146.000 124.760 ;
        RECT 4.400 122.040 146.000 123.440 ;
        RECT 4.000 120.720 146.000 122.040 ;
        RECT 4.400 119.320 146.000 120.720 ;
        RECT 4.000 118.000 146.000 119.320 ;
        RECT 4.400 116.600 146.000 118.000 ;
        RECT 4.000 115.280 146.000 116.600 ;
        RECT 4.400 113.880 146.000 115.280 ;
        RECT 4.000 112.560 146.000 113.880 ;
        RECT 4.400 111.160 145.600 112.560 ;
        RECT 4.000 109.840 146.000 111.160 ;
        RECT 4.400 108.440 146.000 109.840 ;
        RECT 4.000 107.120 146.000 108.440 ;
        RECT 4.400 105.720 146.000 107.120 ;
        RECT 4.000 104.400 146.000 105.720 ;
        RECT 4.400 103.000 146.000 104.400 ;
        RECT 4.000 101.680 146.000 103.000 ;
        RECT 4.400 100.280 146.000 101.680 ;
        RECT 4.000 98.960 146.000 100.280 ;
        RECT 4.400 97.560 146.000 98.960 ;
        RECT 4.000 96.240 146.000 97.560 ;
        RECT 4.400 94.840 146.000 96.240 ;
        RECT 4.000 93.520 146.000 94.840 ;
        RECT 4.400 92.120 146.000 93.520 ;
        RECT 4.000 90.800 146.000 92.120 ;
        RECT 4.400 89.400 146.000 90.800 ;
        RECT 4.000 88.080 146.000 89.400 ;
        RECT 4.400 86.680 146.000 88.080 ;
        RECT 4.000 85.360 146.000 86.680 ;
        RECT 4.400 83.960 146.000 85.360 ;
        RECT 4.000 82.640 146.000 83.960 ;
        RECT 4.400 81.240 146.000 82.640 ;
        RECT 4.000 79.920 146.000 81.240 ;
        RECT 4.400 78.520 146.000 79.920 ;
        RECT 4.000 77.200 146.000 78.520 ;
        RECT 4.400 75.800 146.000 77.200 ;
        RECT 4.000 74.480 146.000 75.800 ;
        RECT 4.400 73.080 146.000 74.480 ;
        RECT 4.000 71.760 146.000 73.080 ;
        RECT 4.400 70.360 146.000 71.760 ;
        RECT 4.000 69.040 146.000 70.360 ;
        RECT 4.400 67.640 146.000 69.040 ;
        RECT 4.000 66.320 146.000 67.640 ;
        RECT 4.400 64.920 146.000 66.320 ;
        RECT 4.000 63.600 146.000 64.920 ;
        RECT 4.400 62.200 146.000 63.600 ;
        RECT 4.000 60.880 146.000 62.200 ;
        RECT 4.400 59.480 146.000 60.880 ;
        RECT 4.000 58.160 146.000 59.480 ;
        RECT 4.400 56.760 146.000 58.160 ;
        RECT 4.000 55.440 146.000 56.760 ;
        RECT 4.400 54.040 146.000 55.440 ;
        RECT 4.000 52.720 146.000 54.040 ;
        RECT 4.400 51.320 146.000 52.720 ;
        RECT 4.000 50.000 146.000 51.320 ;
        RECT 4.400 48.600 146.000 50.000 ;
        RECT 4.000 47.280 146.000 48.600 ;
        RECT 4.400 45.880 146.000 47.280 ;
        RECT 4.000 44.560 146.000 45.880 ;
        RECT 4.400 43.160 146.000 44.560 ;
        RECT 4.000 41.840 146.000 43.160 ;
        RECT 4.400 40.440 146.000 41.840 ;
        RECT 4.000 39.120 146.000 40.440 ;
        RECT 4.400 37.760 146.000 39.120 ;
        RECT 4.400 37.720 145.600 37.760 ;
        RECT 4.000 36.400 145.600 37.720 ;
        RECT 4.400 36.360 145.600 36.400 ;
        RECT 4.400 35.000 146.000 36.360 ;
        RECT 4.000 33.680 146.000 35.000 ;
        RECT 4.400 32.280 146.000 33.680 ;
        RECT 4.000 30.960 146.000 32.280 ;
        RECT 4.400 29.560 146.000 30.960 ;
        RECT 4.000 28.240 146.000 29.560 ;
        RECT 4.400 26.840 146.000 28.240 ;
        RECT 4.000 25.520 146.000 26.840 ;
        RECT 4.400 24.120 146.000 25.520 ;
        RECT 4.000 22.800 146.000 24.120 ;
        RECT 4.400 21.400 146.000 22.800 ;
        RECT 4.000 10.715 146.000 21.400 ;
      LAYER met4 ;
        RECT 8.575 56.615 14.120 109.985 ;
        RECT 16.920 56.615 17.185 109.985 ;
  END
END tbu
END LIBRARY

