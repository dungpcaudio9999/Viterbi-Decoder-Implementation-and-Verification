module piso (clk,
    fifo_empty_i,
    fifo_rd_en_o,
    rst_n,
    valid_serial_o,
    data_serial_o,
    fifo_data_i);
 input clk;
 input fifo_empty_i;
 output fifo_rd_en_o;
 input rst_n;
 output valid_serial_o;
 output [1:0] data_serial_o;
 input [15:0] fifo_data_i;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire \count[0] ;
 wire \count[1] ;
 wire \count[2] ;
 wire \count[3] ;
 wire \shift_reg[10] ;
 wire \shift_reg[11] ;
 wire \shift_reg[12] ;
 wire \shift_reg[13] ;
 wire \shift_reg[14] ;
 wire \shift_reg[15] ;
 wire \shift_reg[2] ;
 wire \shift_reg[3] ;
 wire \shift_reg[4] ;
 wire \shift_reg[5] ;
 wire \shift_reg[6] ;
 wire \shift_reg[7] ;
 wire \shift_reg[8] ;
 wire \shift_reg[9] ;
 wire \state[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 sky130_fd_sc_hd__inv_2 _046_ (.A(\state[1] ),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _047_ (.A(\count[0] ),
    .Y(_018_));
 sky130_fd_sc_hd__nor2_1 _048_ (.A(net21),
    .B(\state[1] ),
    .Y(_019_));
 sky130_fd_sc_hd__or2_1 _049_ (.A(net21),
    .B(\state[1] ),
    .X(_020_));
 sky130_fd_sc_hd__nor2_1 _050_ (.A(net17),
    .B(net34),
    .Y(_037_));
 sky130_fd_sc_hd__and2b_1 _051_ (.A_N(\state[1] ),
    .B(net21),
    .X(_021_));
 sky130_fd_sc_hd__nor2_1 _052_ (.A(\count[0] ),
    .B(\count[1] ),
    .Y(_022_));
 sky130_fd_sc_hd__and2b_1 _053_ (.A_N(\count[2] ),
    .B(_022_),
    .X(_023_));
 sky130_fd_sc_hd__or4_1 _054_ (.A(\count[2] ),
    .B(\count[3] ),
    .C(\count[0] ),
    .D(\count[1] ),
    .X(_024_));
 sky130_fd_sc_hd__and2b_1 _055_ (.A_N(net21),
    .B(\state[1] ),
    .X(_025_));
 sky130_fd_sc_hd__a21o_1 _056_ (.A1(net30),
    .A2(net26),
    .B1(net33),
    .X(_038_));
 sky130_fd_sc_hd__a31o_1 _057_ (.A1(_018_),
    .A2(net28),
    .A3(net25),
    .B1(net32),
    .X(_039_));
 sky130_fd_sc_hd__and2_1 _058_ (.A(\count[0] ),
    .B(\count[1] ),
    .X(_026_));
 sky130_fd_sc_hd__o31a_1 _059_ (.A1(net32),
    .A2(_022_),
    .A3(_026_),
    .B1(_038_),
    .X(_040_));
 sky130_fd_sc_hd__and3b_1 _060_ (.A_N(_022_),
    .B(net25),
    .C(\count[2] ),
    .X(_027_));
 sky130_fd_sc_hd__a311o_1 _061_ (.A1(\count[3] ),
    .A2(_023_),
    .A3(net25),
    .B1(_027_),
    .C1(net32),
    .X(_041_));
 sky130_fd_sc_hd__and3b_1 _062_ (.A_N(_023_),
    .B(net25),
    .C(\count[3] ),
    .X(_042_));
 sky130_fd_sc_hd__a32o_1 _063_ (.A1(\shift_reg[14] ),
    .A2(net29),
    .A3(net25),
    .B1(net6),
    .B2(net32),
    .X(_043_));
 sky130_fd_sc_hd__a32o_1 _064_ (.A1(\shift_reg[15] ),
    .A2(net30),
    .A3(net24),
    .B1(net7),
    .B2(net33),
    .X(_044_));
 sky130_fd_sc_hd__a22o_1 _065_ (.A1(\shift_reg[2] ),
    .A2(_019_),
    .B1(net32),
    .B2(net1),
    .X(_000_));
 sky130_fd_sc_hd__a22o_1 _066_ (.A1(\shift_reg[3] ),
    .A2(_019_),
    .B1(net32),
    .B2(net8),
    .X(_001_));
 sky130_fd_sc_hd__a32o_1 _067_ (.A1(\shift_reg[2] ),
    .A2(net27),
    .A3(net23),
    .B1(net9),
    .B2(net36),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _068_ (.A0(\shift_reg[4] ),
    .A1(_028_),
    .S(net35),
    .X(_002_));
 sky130_fd_sc_hd__a32o_1 _069_ (.A1(\shift_reg[3] ),
    .A2(net27),
    .A3(net23),
    .B1(net10),
    .B2(net36),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _070_ (.A0(\shift_reg[5] ),
    .A1(_029_),
    .S(net35),
    .X(_003_));
 sky130_fd_sc_hd__a32o_1 _071_ (.A1(\shift_reg[4] ),
    .A2(net27),
    .A3(net23),
    .B1(net11),
    .B2(net36),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _072_ (.A0(\shift_reg[6] ),
    .A1(_030_),
    .S(net35),
    .X(_004_));
 sky130_fd_sc_hd__a32o_1 _073_ (.A1(\shift_reg[5] ),
    .A2(net27),
    .A3(net23),
    .B1(net12),
    .B2(net36),
    .X(_031_));
 sky130_fd_sc_hd__mux2_1 _074_ (.A0(\shift_reg[7] ),
    .A1(_031_),
    .S(net35),
    .X(_005_));
 sky130_fd_sc_hd__a32o_1 _075_ (.A1(\shift_reg[6] ),
    .A2(net28),
    .A3(net24),
    .B1(net13),
    .B2(net36),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _076_ (.A0(\shift_reg[8] ),
    .A1(_032_),
    .S(net35),
    .X(_006_));
 sky130_fd_sc_hd__a32o_1 _077_ (.A1(\shift_reg[7] ),
    .A2(net27),
    .A3(net23),
    .B1(net14),
    .B2(net36),
    .X(_033_));
 sky130_fd_sc_hd__mux2_1 _078_ (.A0(\shift_reg[9] ),
    .A1(_033_),
    .S(net34),
    .X(_007_));
 sky130_fd_sc_hd__a32o_1 _079_ (.A1(\shift_reg[8] ),
    .A2(net27),
    .A3(net23),
    .B1(net15),
    .B2(net37),
    .X(_034_));
 sky130_fd_sc_hd__mux2_1 _080_ (.A0(\shift_reg[10] ),
    .A1(_034_),
    .S(net34),
    .X(_008_));
 sky130_fd_sc_hd__a32o_1 _081_ (.A1(\shift_reg[9] ),
    .A2(net29),
    .A3(net24),
    .B1(net16),
    .B2(net37),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _082_ (.A0(\shift_reg[11] ),
    .A1(_035_),
    .S(net34),
    .X(_009_));
 sky130_fd_sc_hd__a32o_1 _083_ (.A1(\shift_reg[10] ),
    .A2(net29),
    .A3(net24),
    .B1(net2),
    .B2(net37),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _084_ (.A0(\shift_reg[12] ),
    .A1(_036_),
    .S(_020_),
    .X(_010_));
 sky130_fd_sc_hd__a32o_1 _085_ (.A1(\shift_reg[11] ),
    .A2(net29),
    .A3(net24),
    .B1(net3),
    .B2(net37),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _086_ (.A0(\shift_reg[13] ),
    .A1(_014_),
    .S(net34),
    .X(_011_));
 sky130_fd_sc_hd__a32o_1 _087_ (.A1(\shift_reg[12] ),
    .A2(net29),
    .A3(net26),
    .B1(net4),
    .B2(net37),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _088_ (.A0(\shift_reg[14] ),
    .A1(_015_),
    .S(_020_),
    .X(_012_));
 sky130_fd_sc_hd__a32o_1 _089_ (.A1(\shift_reg[13] ),
    .A2(net29),
    .A3(net26),
    .B1(net5),
    .B2(net37),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _090_ (.A0(\shift_reg[15] ),
    .A1(_016_),
    .S(net34),
    .X(_013_));
 sky130_fd_sc_hd__a21o_1 _091_ (.A1(net30),
    .A2(net25),
    .B1(net33),
    .X(_045_));
 sky130_fd_sc_hd__dfrtp_1 _092_ (.CLK(clknet_1_0__leaf_clk),
    .D(_000_),
    .RESET_B(net38),
    .Q(\shift_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _093_ (.CLK(clknet_1_0__leaf_clk),
    .D(_001_),
    .RESET_B(net38),
    .Q(\shift_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _094_ (.CLK(clknet_1_0__leaf_clk),
    .D(_002_),
    .RESET_B(net38),
    .Q(\shift_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _095_ (.CLK(clknet_1_0__leaf_clk),
    .D(_003_),
    .RESET_B(net38),
    .Q(\shift_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _096_ (.CLK(clknet_1_0__leaf_clk),
    .D(_004_),
    .RESET_B(net38),
    .Q(\shift_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _097_ (.CLK(clknet_1_0__leaf_clk),
    .D(_005_),
    .RESET_B(net38),
    .Q(\shift_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _098_ (.CLK(clknet_1_0__leaf_clk),
    .D(_006_),
    .RESET_B(net39),
    .Q(\shift_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _099_ (.CLK(clknet_1_1__leaf_clk),
    .D(_007_),
    .RESET_B(net39),
    .Q(\shift_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _100_ (.CLK(clknet_1_1__leaf_clk),
    .D(_008_),
    .RESET_B(net39),
    .Q(\shift_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _101_ (.CLK(clknet_1_1__leaf_clk),
    .D(_009_),
    .RESET_B(net39),
    .Q(\shift_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _102_ (.CLK(clknet_1_1__leaf_clk),
    .D(_010_),
    .RESET_B(net40),
    .Q(\shift_reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 _103_ (.CLK(clknet_1_1__leaf_clk),
    .D(_011_),
    .RESET_B(net39),
    .Q(\shift_reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 _104_ (.CLK(clknet_1_1__leaf_clk),
    .D(_012_),
    .RESET_B(net41),
    .Q(\shift_reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 _105_ (.CLK(clknet_1_1__leaf_clk),
    .D(_013_),
    .RESET_B(net42),
    .Q(\shift_reg[15] ));
 sky130_fd_sc_hd__dfrtp_1 _106_ (.CLK(clknet_1_1__leaf_clk),
    .D(_037_),
    .RESET_B(net42),
    .Q(net21));
 sky130_fd_sc_hd__dfrtp_1 _107_ (.CLK(clknet_1_0__leaf_clk),
    .D(_043_),
    .RESET_B(net40),
    .Q(net19));
 sky130_fd_sc_hd__dfrtp_1 _108_ (.CLK(clknet_1_1__leaf_clk),
    .D(_044_),
    .RESET_B(net41),
    .Q(net20));
 sky130_fd_sc_hd__dfrtp_1 _109_ (.CLK(clknet_1_1__leaf_clk),
    .D(_045_),
    .RESET_B(net41),
    .Q(net22));
 sky130_fd_sc_hd__dfrtp_1 _110_ (.CLK(clknet_1_0__leaf_clk),
    .D(_039_),
    .RESET_B(net40),
    .Q(\count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _111_ (.CLK(clknet_1_1__leaf_clk),
    .D(_040_),
    .RESET_B(net40),
    .Q(\count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _112_ (.CLK(clknet_1_0__leaf_clk),
    .D(_041_),
    .RESET_B(net40),
    .Q(\count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _113_ (.CLK(clknet_1_0__leaf_clk),
    .D(_042_),
    .RESET_B(net40),
    .Q(\count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _114_ (.CLK(clknet_1_1__leaf_clk),
    .D(_038_),
    .RESET_B(net41),
    .Q(\state[1] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_65 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(fifo_data_i[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(fifo_data_i[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(fifo_data_i[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(fifo_data_i[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(fifo_data_i[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(fifo_data_i[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(fifo_data_i[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(fifo_data_i[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(fifo_data_i[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(fifo_data_i[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(fifo_data_i[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(fifo_data_i[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(fifo_data_i[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(fifo_data_i[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(fifo_data_i[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(fifo_data_i[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(fifo_empty_i),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(rst_n),
    .X(net18));
 sky130_fd_sc_hd__buf_4 output19 (.A(net19),
    .X(data_serial_o[0]));
 sky130_fd_sc_hd__buf_4 output20 (.A(net20),
    .X(data_serial_o[1]));
 sky130_fd_sc_hd__buf_4 output21 (.A(net21),
    .X(fifo_rd_en_o));
 sky130_fd_sc_hd__buf_4 output22 (.A(net22),
    .X(valid_serial_o));
 sky130_fd_sc_hd__clkbuf_2 fanout23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 fanout24 (.A(net26),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout25 (.A(net26),
    .X(net25));
 sky130_fd_sc_hd__buf_1 fanout26 (.A(_025_),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__buf_1 fanout28 (.A(net31),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 fanout29 (.A(net31),
    .X(net29));
 sky130_fd_sc_hd__buf_1 fanout30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__buf_1 fanout31 (.A(_024_),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 fanout32 (.A(_021_),
    .X(net32));
 sky130_fd_sc_hd__buf_1 fanout33 (.A(_021_),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 fanout34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 fanout35 (.A(_020_),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout36 (.A(_017_),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 fanout37 (.A(_017_),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 fanout39 (.A(net42),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 fanout40 (.A(net42),
    .X(net40));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 fanout42 (.A(net18),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload0 (.A(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(fifo_data_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(fifo_data_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(fifo_data_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(fifo_data_i[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(fifo_data_i[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(fifo_data_i[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(fifo_data_i[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(fifo_data_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(fifo_data_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(fifo_data_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(fifo_data_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(fifo_data_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(fifo_data_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(fifo_data_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(fifo_data_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(fifo_data_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(fifo_empty_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(rst_n));
 sky130_fd_sc_hd__decap_4 FILLER_0_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_101 ();
endmodule
