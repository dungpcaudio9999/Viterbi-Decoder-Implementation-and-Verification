magic
tech sky130A
magscale 1 2
timestamp 1769198312
<< viali >>
rect 2513 17289 2547 17323
rect 3065 17289 3099 17323
rect 3617 17289 3651 17323
rect 6009 17289 6043 17323
rect 7481 17289 7515 17323
rect 8033 17289 8067 17323
rect 8585 17289 8619 17323
rect 9689 17289 9723 17323
rect 10241 17289 10275 17323
rect 11069 17289 11103 17323
rect 16405 17289 16439 17323
rect 2145 17221 2179 17255
rect 3893 17221 3927 17255
rect 4353 17221 4387 17255
rect 4629 17221 4663 17255
rect 5825 17221 5859 17255
rect 6653 17221 6687 17255
rect 8217 17221 8251 17255
rect 8769 17221 8803 17255
rect 10425 17221 10459 17255
rect 15485 17221 15519 17255
rect 17233 17221 17267 17255
rect 1501 17153 1535 17187
rect 1777 17153 1811 17187
rect 2605 17153 2639 17187
rect 3157 17153 3191 17187
rect 4813 17153 4847 17187
rect 5365 17153 5399 17187
rect 6101 17153 6135 17187
rect 6837 17153 6871 17187
rect 7021 17153 7055 17187
rect 7113 17153 7147 17187
rect 7573 17153 7607 17187
rect 8953 17153 8987 17187
rect 9229 17153 9263 17187
rect 9781 17153 9815 17187
rect 10885 17153 10919 17187
rect 11161 17153 11195 17187
rect 11529 17153 11563 17187
rect 12541 17153 12575 17187
rect 13645 17153 13679 17187
rect 13746 17157 13780 17191
rect 14197 17153 14231 17187
rect 15301 17153 15335 17187
rect 15669 17153 15703 17187
rect 15761 17153 15795 17187
rect 15945 17153 15979 17187
rect 16306 17153 16340 17187
rect 16681 17153 16715 17187
rect 16865 17153 16899 17187
rect 17601 17153 17635 17187
rect 18521 17153 18555 17187
rect 5181 17085 5215 17119
rect 11805 17085 11839 17119
rect 12817 17085 12851 17119
rect 14473 17085 14507 17119
rect 18245 17085 18279 17119
rect 1961 17017 1995 17051
rect 2789 17017 2823 17051
rect 4537 17017 4571 17051
rect 6469 17017 6503 17051
rect 8401 17017 8435 17051
rect 10609 17017 10643 17051
rect 15117 17017 15151 17051
rect 17049 17017 17083 17051
rect 1685 16949 1719 16983
rect 2237 16949 2271 16983
rect 3341 16949 3375 16983
rect 3985 16949 4019 16983
rect 4997 16949 5031 16983
rect 5549 16949 5583 16983
rect 6929 16949 6963 16983
rect 7297 16949 7331 16983
rect 7757 16949 7791 16983
rect 9137 16949 9171 16983
rect 9413 16949 9447 16983
rect 9965 16949 9999 16983
rect 11345 16949 11379 16983
rect 13461 16949 13495 16983
rect 13921 16949 13955 16983
rect 15945 16949 15979 16983
rect 16129 16949 16163 16983
rect 17417 16949 17451 16983
rect 1961 16745 1995 16779
rect 4169 16745 4203 16779
rect 4721 16745 4755 16779
rect 6561 16745 6595 16779
rect 12265 16745 12299 16779
rect 14657 16745 14691 16779
rect 15485 16745 15519 16779
rect 17509 16745 17543 16779
rect 2053 16677 2087 16711
rect 9873 16677 9907 16711
rect 12081 16677 12115 16711
rect 13277 16677 13311 16711
rect 14933 16677 14967 16711
rect 15577 16677 15611 16711
rect 17141 16677 17175 16711
rect 2237 16609 2271 16643
rect 6377 16609 6411 16643
rect 6837 16609 6871 16643
rect 7757 16609 7791 16643
rect 8493 16609 8527 16643
rect 8769 16609 8803 16643
rect 9505 16609 9539 16643
rect 11437 16609 11471 16643
rect 12541 16609 12575 16643
rect 13645 16609 13679 16643
rect 1409 16541 1443 16575
rect 1685 16541 1719 16575
rect 5549 16541 5583 16575
rect 6009 16541 6043 16575
rect 7021 16541 7055 16575
rect 7481 16541 7515 16575
rect 8401 16541 8435 16575
rect 9413 16541 9447 16575
rect 11713 16541 11747 16575
rect 11989 16541 12023 16575
rect 13001 16541 13035 16575
rect 13737 16541 13771 16575
rect 14289 16541 14323 16575
rect 15301 16541 15335 16575
rect 15853 16541 15887 16575
rect 16957 16541 16991 16575
rect 17141 16541 17175 16575
rect 17417 16541 17451 16575
rect 17693 16541 17727 16575
rect 17785 16541 17819 16575
rect 17877 16541 17911 16575
rect 18061 16541 18095 16575
rect 18337 16541 18371 16575
rect 10057 16473 10091 16507
rect 12449 16473 12483 16507
rect 12725 16473 12759 16507
rect 12909 16473 12943 16507
rect 13280 16473 13314 16507
rect 14381 16473 14415 16507
rect 14749 16473 14783 16507
rect 15117 16473 15151 16507
rect 15209 16473 15243 16507
rect 16865 16473 16899 16507
rect 1593 16405 1627 16439
rect 9781 16405 9815 16439
rect 11897 16405 11931 16439
rect 12239 16405 12273 16439
rect 13093 16405 13127 16439
rect 13369 16405 13403 16439
rect 14105 16405 14139 16439
rect 17233 16405 17267 16439
rect 1869 16201 1903 16235
rect 5733 16201 5767 16235
rect 9229 16201 9263 16235
rect 11713 16201 11747 16235
rect 13001 16201 13035 16235
rect 13277 16201 13311 16235
rect 14013 16201 14047 16235
rect 15117 16201 15151 16235
rect 15685 16201 15719 16235
rect 15853 16201 15887 16235
rect 16865 16201 16899 16235
rect 17417 16201 17451 16235
rect 17969 16201 18003 16235
rect 18521 16201 18555 16235
rect 8585 16133 8619 16167
rect 12081 16133 12115 16167
rect 12357 16133 12391 16167
rect 15485 16133 15519 16167
rect 17049 16133 17083 16167
rect 1409 16065 1443 16099
rect 1685 16065 1719 16099
rect 4261 16065 4295 16099
rect 5181 16065 5215 16099
rect 5365 16065 5399 16099
rect 5641 16065 5675 16099
rect 5825 16065 5859 16099
rect 6929 16065 6963 16099
rect 9137 16065 9171 16099
rect 10241 16065 10275 16099
rect 10885 16065 10919 16099
rect 10977 16065 11011 16099
rect 11897 16065 11931 16099
rect 11989 16065 12023 16099
rect 12245 16065 12279 16099
rect 12541 16065 12575 16099
rect 12633 16065 12667 16099
rect 12909 16065 12943 16099
rect 13829 16065 13863 16099
rect 15301 16065 15335 16099
rect 17509 16065 17543 16099
rect 18245 16065 18279 16099
rect 4169 15997 4203 16031
rect 4997 15997 5031 16031
rect 7021 15997 7055 16031
rect 9321 15997 9355 16031
rect 10057 15997 10091 16031
rect 11069 15997 11103 16031
rect 1593 15929 1627 15963
rect 7297 15929 7331 15963
rect 10517 15929 10551 15963
rect 5273 15861 5307 15895
rect 8493 15861 8527 15895
rect 8769 15861 8803 15895
rect 10425 15861 10459 15895
rect 12817 15861 12851 15895
rect 13737 15861 13771 15895
rect 15669 15861 15703 15895
rect 18061 15861 18095 15895
rect 7021 15657 7055 15691
rect 11253 15657 11287 15691
rect 13645 15657 13679 15691
rect 8217 15589 8251 15623
rect 12081 15589 12115 15623
rect 13369 15589 13403 15623
rect 13829 15589 13863 15623
rect 4997 15521 5031 15555
rect 6745 15521 6779 15555
rect 9597 15521 9631 15555
rect 10057 15521 10091 15555
rect 14105 15521 14139 15555
rect 14381 15521 14415 15555
rect 15945 15521 15979 15555
rect 16681 15521 16715 15555
rect 5273 15453 5307 15487
rect 5641 15453 5675 15487
rect 6653 15453 6687 15487
rect 9413 15453 9447 15487
rect 9689 15453 9723 15487
rect 9781 15453 9815 15487
rect 9873 15453 9907 15487
rect 10609 15453 10643 15487
rect 10757 15453 10791 15487
rect 11074 15453 11108 15487
rect 12357 15453 12391 15487
rect 13093 15453 13127 15487
rect 14473 15453 14507 15487
rect 15393 15453 15427 15487
rect 15577 15453 15611 15487
rect 15761 15453 15795 15487
rect 16129 15453 16163 15487
rect 16773 15453 16807 15487
rect 5917 15385 5951 15419
rect 8401 15385 8435 15419
rect 8769 15385 8803 15419
rect 10885 15385 10919 15419
rect 10977 15385 11011 15419
rect 13369 15385 13403 15419
rect 13461 15385 13495 15419
rect 13661 15385 13695 15419
rect 8493 15317 8527 15351
rect 8585 15317 8619 15351
rect 11897 15317 11931 15351
rect 13185 15317 13219 15351
rect 17141 15317 17175 15351
rect 1593 15113 1627 15147
rect 8769 15113 8803 15147
rect 13553 15113 13587 15147
rect 1409 14977 1443 15011
rect 1685 14977 1719 15011
rect 4445 14977 4479 15011
rect 4629 14977 4663 15011
rect 4997 14977 5031 15011
rect 8125 14977 8159 15011
rect 8769 14977 8803 15011
rect 9045 14977 9079 15011
rect 12633 14977 12667 15011
rect 13461 14977 13495 15011
rect 13645 14977 13679 15011
rect 15485 14977 15519 15011
rect 15669 14977 15703 15011
rect 15761 14977 15795 15011
rect 4537 14909 4571 14943
rect 5089 14909 5123 14943
rect 7941 14909 7975 14943
rect 8309 14909 8343 14943
rect 8861 14909 8895 14943
rect 15577 14909 15611 14943
rect 5365 14841 5399 14875
rect 12449 14773 12483 14807
rect 15301 14773 15335 14807
rect 12725 14569 12759 14603
rect 10609 14501 10643 14535
rect 12173 14501 12207 14535
rect 4261 14433 4295 14467
rect 4537 14433 4571 14467
rect 6469 14433 6503 14467
rect 9505 14433 9539 14467
rect 10885 14433 10919 14467
rect 12817 14433 12851 14467
rect 14565 14433 14599 14467
rect 4169 14365 4203 14399
rect 6561 14365 6595 14399
rect 8585 14365 8619 14399
rect 8769 14365 8803 14399
rect 9321 14365 9355 14399
rect 10057 14365 10091 14399
rect 10149 14365 10183 14399
rect 10241 14365 10275 14399
rect 10425 14365 10459 14399
rect 10977 14365 11011 14399
rect 11437 14365 11471 14399
rect 13093 14365 13127 14399
rect 16405 14365 16439 14399
rect 16589 14365 16623 14399
rect 8677 14297 8711 14331
rect 9413 14297 9447 14331
rect 12449 14297 12483 14331
rect 14197 14297 14231 14331
rect 14381 14297 14415 14331
rect 6929 14229 6963 14263
rect 8953 14229 8987 14263
rect 9781 14229 9815 14263
rect 11253 14229 11287 14263
rect 12357 14229 12391 14263
rect 12541 14229 12575 14263
rect 16497 14229 16531 14263
rect 4997 14025 5031 14059
rect 7205 14025 7239 14059
rect 9597 14025 9631 14059
rect 10793 14025 10827 14059
rect 13737 14025 13771 14059
rect 16957 14025 16991 14059
rect 17417 14025 17451 14059
rect 4537 13957 4571 13991
rect 5365 13957 5399 13991
rect 6929 13957 6963 13991
rect 7481 13957 7515 13991
rect 8493 13957 8527 13991
rect 8585 13957 8619 13991
rect 13093 13957 13127 13991
rect 1409 13889 1443 13923
rect 1685 13889 1719 13923
rect 5457 13889 5491 13923
rect 6653 13889 6687 13923
rect 6837 13889 6871 13923
rect 7021 13889 7055 13923
rect 7297 13889 7331 13923
rect 7665 13889 7699 13923
rect 8401 13889 8435 13923
rect 8769 13889 8803 13923
rect 8861 13889 8895 13923
rect 9781 13889 9815 13923
rect 11069 13889 11103 13923
rect 11253 13889 11287 13923
rect 11529 13889 11563 13923
rect 11621 13889 11655 13923
rect 11897 13889 11931 13923
rect 12081 13889 12115 13923
rect 12357 13889 12391 13923
rect 12633 13889 12667 13923
rect 13001 13889 13035 13923
rect 13553 13889 13587 13923
rect 13645 13889 13679 13923
rect 14473 13889 14507 13923
rect 15853 13889 15887 13923
rect 16037 13889 16071 13923
rect 16129 13889 16163 13923
rect 16221 13889 16255 13923
rect 17049 13889 17083 13923
rect 5273 13821 5307 13855
rect 9965 13821 9999 13855
rect 10977 13821 11011 13855
rect 11161 13821 11195 13855
rect 12449 13821 12483 13855
rect 13277 13821 13311 13855
rect 13369 13821 13403 13855
rect 14381 13821 14415 13855
rect 15209 13821 15243 13855
rect 16497 13821 16531 13855
rect 16865 13821 16899 13855
rect 4905 13753 4939 13787
rect 8217 13753 8251 13787
rect 1593 13685 1627 13719
rect 5825 13685 5859 13719
rect 13921 13685 13955 13719
rect 4353 13481 4387 13515
rect 5917 13481 5951 13515
rect 6469 13481 6503 13515
rect 13645 13481 13679 13515
rect 14289 13481 14323 13515
rect 14473 13481 14507 13515
rect 14657 13481 14691 13515
rect 16589 13481 16623 13515
rect 8677 13413 8711 13447
rect 4077 13345 4111 13379
rect 12725 13345 12759 13379
rect 13001 13345 13035 13379
rect 17141 13345 17175 13379
rect 17785 13345 17819 13379
rect 18245 13345 18279 13379
rect 3985 13277 4019 13311
rect 5457 13277 5491 13311
rect 5733 13277 5767 13311
rect 8401 13277 8435 13311
rect 13645 13277 13679 13311
rect 13921 13277 13955 13311
rect 14749 13277 14783 13311
rect 15393 13277 15427 13311
rect 15485 13277 15519 13311
rect 15669 13277 15703 13311
rect 15761 13277 15795 13311
rect 16221 13277 16255 13311
rect 16405 13277 16439 13311
rect 17233 13277 17267 13311
rect 17877 13277 17911 13311
rect 6101 13209 6135 13243
rect 6285 13209 6319 13243
rect 8677 13209 8711 13243
rect 14105 13209 14139 13243
rect 14305 13209 14339 13243
rect 5549 13141 5583 13175
rect 8493 13141 8527 13175
rect 13829 13141 13863 13175
rect 15209 13141 15243 13175
rect 17601 13141 17635 13175
rect 7941 12937 7975 12971
rect 8585 12937 8619 12971
rect 15025 12869 15059 12903
rect 15669 12869 15703 12903
rect 16037 12869 16071 12903
rect 1409 12801 1443 12835
rect 1685 12801 1719 12835
rect 6009 12801 6043 12835
rect 8125 12801 8159 12835
rect 8217 12801 8251 12835
rect 8360 12801 8394 12835
rect 8493 12791 8527 12825
rect 8841 12801 8875 12835
rect 8950 12801 8984 12835
rect 9050 12804 9084 12838
rect 9229 12801 9263 12835
rect 10425 12801 10459 12835
rect 10609 12801 10643 12835
rect 10793 12801 10827 12835
rect 10885 12801 10919 12835
rect 10977 12801 11011 12835
rect 11069 12801 11103 12835
rect 11253 12801 11287 12835
rect 14933 12801 14967 12835
rect 15189 12801 15223 12835
rect 15485 12801 15519 12835
rect 15761 12801 15795 12835
rect 18061 12801 18095 12835
rect 15853 12733 15887 12767
rect 18337 12733 18371 12767
rect 1593 12665 1627 12699
rect 10977 12665 11011 12699
rect 6101 12597 6135 12631
rect 15393 12597 15427 12631
rect 15761 12597 15795 12631
rect 8585 12393 8619 12427
rect 12449 12393 12483 12427
rect 13369 12393 13403 12427
rect 5365 12325 5399 12359
rect 8401 12325 8435 12359
rect 13093 12325 13127 12359
rect 4445 12257 4479 12291
rect 6009 12257 6043 12291
rect 6101 12257 6135 12291
rect 6929 12257 6963 12291
rect 9321 12257 9355 12291
rect 11345 12257 11379 12291
rect 12817 12257 12851 12291
rect 4353 12189 4387 12223
rect 5181 12189 5215 12223
rect 6837 12189 6871 12223
rect 9137 12189 9171 12223
rect 9413 12189 9447 12223
rect 9597 12189 9631 12223
rect 11253 12189 11287 12223
rect 11897 12189 11931 12223
rect 12173 12189 12207 12223
rect 12725 12189 12759 12223
rect 17141 12189 17175 12223
rect 17417 12189 17451 12223
rect 17877 12189 17911 12223
rect 4813 12121 4847 12155
rect 6193 12121 6227 12155
rect 8769 12121 8803 12155
rect 11805 12121 11839 12155
rect 12265 12121 12299 12155
rect 12449 12121 12483 12155
rect 13185 12121 13219 12155
rect 17233 12121 17267 12155
rect 17693 12121 17727 12155
rect 4721 12053 4755 12087
rect 4997 12053 5031 12087
rect 5089 12053 5123 12087
rect 6561 12053 6595 12087
rect 7205 12053 7239 12087
rect 8569 12053 8603 12087
rect 8953 12053 8987 12087
rect 9505 12053 9539 12087
rect 11621 12053 11655 12087
rect 13385 12053 13419 12087
rect 13553 12053 13587 12087
rect 17601 12053 17635 12087
rect 18061 12053 18095 12087
rect 4261 11849 4295 11883
rect 4445 11849 4479 11883
rect 8493 11849 8527 11883
rect 10701 11849 10735 11883
rect 16129 11849 16163 11883
rect 17049 11849 17083 11883
rect 8585 11781 8619 11815
rect 15025 11781 15059 11815
rect 16313 11781 16347 11815
rect 16957 11781 16991 11815
rect 1409 11713 1443 11747
rect 1685 11713 1719 11747
rect 3433 11713 3467 11747
rect 4077 11713 4111 11747
rect 4353 11713 4387 11747
rect 4537 11713 4571 11747
rect 6561 11713 6595 11747
rect 9873 11713 9907 11747
rect 10333 11713 10367 11747
rect 10425 11713 10459 11747
rect 14013 11713 14047 11747
rect 14197 11713 14231 11747
rect 14289 11713 14323 11747
rect 14473 11713 14507 11747
rect 14749 11713 14783 11747
rect 15301 11713 15335 11747
rect 15393 11713 15427 11747
rect 15485 11713 15519 11747
rect 15669 11713 15703 11747
rect 15761 11713 15795 11747
rect 15945 11713 15979 11747
rect 16221 11713 16255 11747
rect 16399 11713 16433 11747
rect 17693 11713 17727 11747
rect 17877 11713 17911 11747
rect 18061 11713 18095 11747
rect 18245 11713 18279 11747
rect 3341 11645 3375 11679
rect 3801 11645 3835 11679
rect 3893 11645 3927 11679
rect 6653 11645 6687 11679
rect 8769 11645 8803 11679
rect 9689 11645 9723 11679
rect 10057 11645 10091 11679
rect 10241 11645 10275 11679
rect 10517 11645 10551 11679
rect 16865 11645 16899 11679
rect 17969 11645 18003 11679
rect 1593 11577 1627 11611
rect 14197 11577 14231 11611
rect 14565 11577 14599 11611
rect 14657 11577 14691 11611
rect 14933 11577 14967 11611
rect 17509 11577 17543 11611
rect 6929 11509 6963 11543
rect 8125 11509 8159 11543
rect 17417 11509 17451 11543
rect 6837 11305 6871 11339
rect 13461 11305 13495 11339
rect 14841 11305 14875 11339
rect 7297 11169 7331 11203
rect 7481 11169 7515 11203
rect 9229 11169 9263 11203
rect 9505 11169 9539 11203
rect 18061 11169 18095 11203
rect 18153 11169 18187 11203
rect 7205 11101 7239 11135
rect 9137 11101 9171 11135
rect 13737 11101 13771 11135
rect 15025 11101 15059 11135
rect 15117 11101 15151 11135
rect 15301 11101 15335 11135
rect 15393 11101 15427 11135
rect 17969 11101 18003 11135
rect 13461 11033 13495 11067
rect 13645 11033 13679 11067
rect 17601 10965 17635 10999
rect 1593 10761 1627 10795
rect 13369 10761 13403 10795
rect 17233 10761 17267 10795
rect 10977 10693 11011 10727
rect 12541 10693 12575 10727
rect 18153 10693 18187 10727
rect 1409 10625 1443 10659
rect 1685 10625 1719 10659
rect 5273 10625 5307 10659
rect 8677 10625 8711 10659
rect 10425 10625 10459 10659
rect 10885 10625 10919 10659
rect 11069 10625 11103 10659
rect 11713 10625 11747 10659
rect 12817 10625 12851 10659
rect 13093 10625 13127 10659
rect 13185 10625 13219 10659
rect 14197 10625 14231 10659
rect 16681 10625 16715 10659
rect 16957 10625 16991 10659
rect 17049 10625 17083 10659
rect 5365 10557 5399 10591
rect 10517 10557 10551 10591
rect 11805 10557 11839 10591
rect 12173 10557 12207 10591
rect 8493 10489 8527 10523
rect 10793 10489 10827 10523
rect 12081 10489 12115 10523
rect 16773 10489 16807 10523
rect 5641 10421 5675 10455
rect 12541 10421 12575 10455
rect 12725 10421 12759 10455
rect 12909 10421 12943 10455
rect 14289 10421 14323 10455
rect 18061 10421 18095 10455
rect 4629 10217 4663 10251
rect 4813 10217 4847 10251
rect 7757 10217 7791 10251
rect 9137 10217 9171 10251
rect 13001 10217 13035 10251
rect 5181 10149 5215 10183
rect 7021 10149 7055 10183
rect 8217 10149 8251 10183
rect 8953 10149 8987 10183
rect 12909 10149 12943 10183
rect 14841 10149 14875 10183
rect 15669 10149 15703 10183
rect 17417 10149 17451 10183
rect 7389 10081 7423 10115
rect 8677 10081 8711 10115
rect 14289 10081 14323 10115
rect 14381 10081 14415 10115
rect 15025 10081 15059 10115
rect 15209 10081 15243 10115
rect 16773 10081 16807 10115
rect 17693 10081 17727 10115
rect 1409 10013 1443 10047
rect 1685 10013 1719 10047
rect 4905 10013 4939 10047
rect 5273 10013 5307 10047
rect 5457 10013 5491 10047
rect 6469 10013 6503 10047
rect 6653 10013 6687 10047
rect 6837 10013 6871 10047
rect 7941 10013 7975 10047
rect 8585 10013 8619 10047
rect 15301 10013 15335 10047
rect 15761 10013 15795 10047
rect 15945 10013 15979 10047
rect 16221 10013 16255 10047
rect 16313 10013 16347 10047
rect 16497 10013 16531 10047
rect 16681 10013 16715 10047
rect 16865 10013 16899 10047
rect 17049 10013 17083 10047
rect 17325 10013 17359 10047
rect 17877 10013 17911 10047
rect 4445 9945 4479 9979
rect 5181 9945 5215 9979
rect 5365 9945 5399 9979
rect 6561 9945 6595 9979
rect 8125 9945 8159 9979
rect 9321 9945 9355 9979
rect 12541 9945 12575 9979
rect 14473 9945 14507 9979
rect 1593 9877 1627 9911
rect 4645 9877 4679 9911
rect 4997 9877 5031 9911
rect 6009 9877 6043 9911
rect 6285 9877 6319 9911
rect 6929 9877 6963 9911
rect 9111 9877 9145 9911
rect 16037 9877 16071 9911
rect 17969 9877 18003 9911
rect 18337 9877 18371 9911
rect 2237 9673 2271 9707
rect 4629 9673 4663 9707
rect 16681 9673 16715 9707
rect 3341 9605 3375 9639
rect 4537 9605 4571 9639
rect 6101 9605 6135 9639
rect 8125 9605 8159 9639
rect 17049 9605 17083 9639
rect 17417 9605 17451 9639
rect 1593 9537 1627 9571
rect 1685 9537 1719 9571
rect 1869 9537 1903 9571
rect 1961 9537 1995 9571
rect 2105 9537 2139 9571
rect 2329 9537 2363 9571
rect 2789 9537 2823 9571
rect 3249 9537 3283 9571
rect 3433 9537 3467 9571
rect 6193 9537 6227 9571
rect 6561 9537 6595 9571
rect 6653 9537 6687 9571
rect 6929 9537 6963 9571
rect 8033 9537 8067 9571
rect 8309 9537 8343 9571
rect 12265 9537 12299 9571
rect 16865 9537 16899 9571
rect 16957 9537 16991 9571
rect 17233 9537 17267 9571
rect 17325 9537 17359 9571
rect 17601 9537 17635 9571
rect 17785 9537 17819 9571
rect 2697 9469 2731 9503
rect 4445 9469 4479 9503
rect 5641 9469 5675 9503
rect 5917 9469 5951 9503
rect 6377 9469 6411 9503
rect 6837 9469 6871 9503
rect 2513 9401 2547 9435
rect 8309 9401 8343 9435
rect 3065 9333 3099 9367
rect 4997 9333 5031 9367
rect 12357 9333 12391 9367
rect 17601 9333 17635 9367
rect 1961 9129 1995 9163
rect 4353 9129 4387 9163
rect 9413 9129 9447 9163
rect 10241 9129 10275 9163
rect 12449 9129 12483 9163
rect 9597 9061 9631 9095
rect 12173 9061 12207 9095
rect 12633 9061 12667 9095
rect 1685 8993 1719 9027
rect 4445 8993 4479 9027
rect 6193 8993 6227 9027
rect 6653 8993 6687 9027
rect 8033 8993 8067 9027
rect 9781 8993 9815 9027
rect 13461 8993 13495 9027
rect 1593 8925 1627 8959
rect 3433 8925 3467 8959
rect 3985 8925 4019 8959
rect 5825 8925 5859 8959
rect 5917 8925 5951 8959
rect 6101 8925 6135 8959
rect 6285 8925 6319 8959
rect 6469 8925 6503 8959
rect 8125 8925 8159 8959
rect 9873 8925 9907 8959
rect 10793 8925 10827 8959
rect 11069 8925 11103 8959
rect 11897 8925 11931 8959
rect 12909 8925 12943 8959
rect 13093 8925 13127 8959
rect 13553 8925 13587 8959
rect 9459 8891 9493 8925
rect 3617 8857 3651 8891
rect 3801 8857 3835 8891
rect 4629 8857 4663 8891
rect 5457 8857 5491 8891
rect 5641 8857 5675 8891
rect 9229 8857 9263 8891
rect 10517 8857 10551 8891
rect 11989 8857 12023 8891
rect 12173 8857 12207 8891
rect 12265 8857 12299 8891
rect 13277 8857 13311 8891
rect 4077 8789 4111 8823
rect 4169 8789 4203 8823
rect 5181 8789 5215 8823
rect 7757 8789 7791 8823
rect 10701 8789 10735 8823
rect 10885 8789 10919 8823
rect 12465 8789 12499 8823
rect 13921 8789 13955 8823
rect 6837 8585 6871 8619
rect 4997 8517 5031 8551
rect 5825 8517 5859 8551
rect 6469 8517 6503 8551
rect 9781 8517 9815 8551
rect 10149 8517 10183 8551
rect 1869 8449 1903 8483
rect 4905 8449 4939 8483
rect 5549 8449 5583 8483
rect 5917 8449 5951 8483
rect 6377 8449 6411 8483
rect 6653 8449 6687 8483
rect 7573 8449 7607 8483
rect 9505 8449 9539 8483
rect 9597 8449 9631 8483
rect 10057 8449 10091 8483
rect 10241 8449 10275 8483
rect 11989 8449 12023 8483
rect 12633 8449 12667 8483
rect 1593 8381 1627 8415
rect 2513 8381 2547 8415
rect 5181 8381 5215 8415
rect 12081 8381 12115 8415
rect 12541 8381 12575 8415
rect 4537 8313 4571 8347
rect 5365 8313 5399 8347
rect 9781 8313 9815 8347
rect 13001 8313 13035 8347
rect 6101 8245 6135 8279
rect 7757 8245 7791 8279
rect 12265 8245 12299 8279
rect 6929 8041 6963 8075
rect 8033 8041 8067 8075
rect 4721 7973 4755 8007
rect 8585 7973 8619 8007
rect 1409 7905 1443 7939
rect 3525 7905 3559 7939
rect 4445 7905 4479 7939
rect 7481 7905 7515 7939
rect 1685 7837 1719 7871
rect 2513 7837 2547 7871
rect 4353 7837 4387 7871
rect 6285 7837 6319 7871
rect 6469 7837 6503 7871
rect 6561 7837 6595 7871
rect 6653 7837 6687 7871
rect 7021 7837 7055 7871
rect 7297 7837 7331 7871
rect 7849 7837 7883 7871
rect 8309 7837 8343 7871
rect 18061 7837 18095 7871
rect 7665 7769 7699 7803
rect 8401 7769 8435 7803
rect 18337 7769 18371 7803
rect 8217 7701 8251 7735
rect 1593 7497 1627 7531
rect 9137 7497 9171 7531
rect 9505 7497 9539 7531
rect 12081 7497 12115 7531
rect 13277 7497 13311 7531
rect 2145 7429 2179 7463
rect 3433 7429 3467 7463
rect 8953 7429 8987 7463
rect 14013 7429 14047 7463
rect 1409 7361 1443 7395
rect 1869 7361 1903 7395
rect 2053 7361 2087 7395
rect 2237 7361 2271 7395
rect 2789 7361 2823 7395
rect 3157 7361 3191 7395
rect 4629 7361 4663 7395
rect 4905 7361 4939 7395
rect 5365 7361 5399 7395
rect 6561 7361 6595 7395
rect 6653 7361 6687 7395
rect 6837 7361 6871 7395
rect 6929 7361 6963 7395
rect 7021 7361 7055 7395
rect 7205 7361 7239 7395
rect 7849 7361 7883 7395
rect 9229 7361 9263 7395
rect 9321 7361 9355 7395
rect 10333 7361 10367 7395
rect 10517 7361 10551 7395
rect 10885 7361 10919 7395
rect 11713 7361 11747 7395
rect 12817 7361 12851 7395
rect 13001 7361 13035 7395
rect 13461 7361 13495 7395
rect 13829 7361 13863 7395
rect 14105 7361 14139 7395
rect 14197 7361 14231 7395
rect 1685 7293 1719 7327
rect 2513 7293 2547 7327
rect 4721 7293 4755 7327
rect 4813 7293 4847 7327
rect 5089 7293 5123 7327
rect 5549 7293 5583 7327
rect 10241 7293 10275 7327
rect 11805 7293 11839 7327
rect 7021 7225 7055 7259
rect 7665 7225 7699 7259
rect 10885 7225 10919 7259
rect 5181 7157 5215 7191
rect 6377 7157 6411 7191
rect 13185 7157 13219 7191
rect 14381 7157 14415 7191
rect 8217 6953 8251 6987
rect 9137 6953 9171 6987
rect 14565 6953 14599 6987
rect 14841 6885 14875 6919
rect 4813 6817 4847 6851
rect 10057 6817 10091 6851
rect 10241 6817 10275 6851
rect 12909 6817 12943 6851
rect 13093 6817 13127 6851
rect 14105 6817 14139 6851
rect 2145 6749 2179 6783
rect 4537 6749 4571 6783
rect 7757 6749 7791 6783
rect 8125 6749 8159 6783
rect 8401 6749 8435 6783
rect 8769 6749 8803 6783
rect 8953 6749 8987 6783
rect 9229 6749 9263 6783
rect 9597 6749 9631 6783
rect 9781 6749 9815 6783
rect 9873 6749 9907 6783
rect 9965 6749 9999 6783
rect 11069 6749 11103 6783
rect 11253 6749 11287 6783
rect 11345 6749 11379 6783
rect 11437 6749 11471 6783
rect 12265 6749 12299 6783
rect 12541 6749 12575 6783
rect 13185 6749 13219 6783
rect 14289 6749 14323 6783
rect 14381 6749 14415 6783
rect 14657 6749 14691 6783
rect 15209 6749 15243 6783
rect 1961 6681 1995 6715
rect 4629 6681 4663 6715
rect 8677 6681 8711 6715
rect 11713 6681 11747 6715
rect 2329 6613 2363 6647
rect 4169 6613 4203 6647
rect 7941 6613 7975 6647
rect 9413 6613 9447 6647
rect 12357 6613 12391 6647
rect 12725 6613 12759 6647
rect 13553 6613 13587 6647
rect 14749 6613 14783 6647
rect 1593 6409 1627 6443
rect 6377 6409 6411 6443
rect 8861 6409 8895 6443
rect 13737 6409 13771 6443
rect 1409 6273 1443 6307
rect 1961 6273 1995 6307
rect 2789 6273 2823 6307
rect 6561 6273 6595 6307
rect 6837 6273 6871 6307
rect 7021 6273 7055 6307
rect 7941 6273 7975 6307
rect 8217 6273 8251 6307
rect 8777 6273 8811 6307
rect 9045 6273 9079 6307
rect 11069 6273 11103 6307
rect 11161 6273 11195 6307
rect 11529 6273 11563 6307
rect 11621 6273 11655 6307
rect 11805 6273 11839 6307
rect 11897 6273 11931 6307
rect 12173 6273 12207 6307
rect 12357 6273 12391 6307
rect 13001 6273 13035 6307
rect 13185 6273 13219 6307
rect 13369 6273 13403 6307
rect 13553 6273 13587 6307
rect 2053 6205 2087 6239
rect 2881 6205 2915 6239
rect 13277 6205 13311 6239
rect 3157 6137 3191 6171
rect 6653 6137 6687 6171
rect 6745 6137 6779 6171
rect 11345 6137 11379 6171
rect 2329 6069 2363 6103
rect 7665 6069 7699 6103
rect 8125 6069 8159 6103
rect 9137 6069 9171 6103
rect 12081 6069 12115 6103
rect 12173 6069 12207 6103
rect 1409 5865 1443 5899
rect 6377 5865 6411 5899
rect 7021 5865 7055 5899
rect 7297 5865 7331 5899
rect 9413 5865 9447 5899
rect 13093 5865 13127 5899
rect 9689 5797 9723 5831
rect 5457 5729 5491 5763
rect 1869 5661 1903 5695
rect 2145 5661 2179 5695
rect 2513 5661 2547 5695
rect 2697 5661 2731 5695
rect 2789 5661 2823 5695
rect 2973 5661 3007 5695
rect 4537 5661 4571 5695
rect 4629 5661 4663 5695
rect 4813 5661 4847 5695
rect 4997 5661 5031 5695
rect 5273 5661 5307 5695
rect 5733 5661 5767 5695
rect 5917 5661 5951 5695
rect 6009 5661 6043 5695
rect 6101 5661 6135 5695
rect 6469 5661 6503 5695
rect 6561 5661 6595 5695
rect 6745 5661 6779 5695
rect 6837 5661 6871 5695
rect 7665 5661 7699 5695
rect 9965 5661 9999 5695
rect 12449 5661 12483 5695
rect 12633 5661 12667 5695
rect 12725 5661 12759 5695
rect 12817 5661 12851 5695
rect 12909 5661 12943 5695
rect 2237 5593 2271 5627
rect 7281 5593 7315 5627
rect 7481 5593 7515 5627
rect 7849 5593 7883 5627
rect 9229 5593 9263 5627
rect 9689 5593 9723 5627
rect 9873 5593 9907 5627
rect 2329 5525 2363 5559
rect 2973 5525 3007 5559
rect 5089 5525 5123 5559
rect 7113 5525 7147 5559
rect 9429 5525 9463 5559
rect 9597 5525 9631 5559
rect 4997 5321 5031 5355
rect 6101 5321 6135 5355
rect 10977 5321 11011 5355
rect 13461 5321 13495 5355
rect 3617 5253 3651 5287
rect 3709 5253 3743 5287
rect 6469 5253 6503 5287
rect 6929 5253 6963 5287
rect 10609 5253 10643 5287
rect 12541 5253 12575 5287
rect 12909 5253 12943 5287
rect 1409 5185 1443 5219
rect 1685 5185 1719 5219
rect 3433 5185 3467 5219
rect 3801 5185 3835 5219
rect 4261 5185 4295 5219
rect 4445 5185 4479 5219
rect 4537 5185 4571 5219
rect 4813 5185 4847 5219
rect 5917 5185 5951 5219
rect 6377 5185 6411 5219
rect 6561 5185 6595 5219
rect 6837 5185 6871 5219
rect 7113 5185 7147 5219
rect 7941 5185 7975 5219
rect 9229 5185 9263 5219
rect 10517 5185 10551 5219
rect 10793 5185 10827 5219
rect 11072 5185 11106 5219
rect 11253 5185 11287 5219
rect 11345 5185 11379 5219
rect 12633 5185 12667 5219
rect 13001 5185 13035 5219
rect 13093 5185 13127 5219
rect 13369 5185 13403 5219
rect 14013 5185 14047 5219
rect 4629 5117 4663 5151
rect 5733 5117 5767 5151
rect 7849 5117 7883 5151
rect 9137 5117 9171 5151
rect 13461 5117 13495 5151
rect 3985 5049 4019 5083
rect 7113 5049 7147 5083
rect 9597 5049 9631 5083
rect 11345 5049 11379 5083
rect 1593 4981 1627 5015
rect 7665 4981 7699 5015
rect 12725 4981 12759 5015
rect 13185 4981 13219 5015
rect 14105 4981 14139 5015
rect 6561 4777 6595 4811
rect 8677 4777 8711 4811
rect 3065 4641 3099 4675
rect 6745 4641 6779 4675
rect 8493 4641 8527 4675
rect 10885 4641 10919 4675
rect 12541 4641 12575 4675
rect 14565 4641 14599 4675
rect 14749 4641 14783 4675
rect 14933 4641 14967 4675
rect 2053 4573 2087 4607
rect 6837 4573 6871 4607
rect 8217 4573 8251 4607
rect 8309 4573 8343 4607
rect 8401 4573 8435 4607
rect 10793 4573 10827 4607
rect 11253 4573 11287 4607
rect 12725 4573 12759 4607
rect 13001 4573 13035 4607
rect 13185 4573 13219 4607
rect 14473 4573 14507 4607
rect 15117 4573 15151 4607
rect 11345 4505 11379 4539
rect 7941 4437 7975 4471
rect 11161 4437 11195 4471
rect 12909 4437 12943 4471
rect 13093 4437 13127 4471
rect 14105 4437 14139 4471
rect 2513 4233 2547 4267
rect 5365 4233 5399 4267
rect 3893 4165 3927 4199
rect 1961 4097 1995 4131
rect 2329 4097 2363 4131
rect 4629 4097 4663 4131
rect 5457 4097 5491 4131
rect 6745 4097 6779 4131
rect 12449 4097 12483 4131
rect 12633 4097 12667 4131
rect 1685 4029 1719 4063
rect 2145 4029 2179 4063
rect 4905 4029 4939 4063
rect 5641 4029 5675 4063
rect 6837 4029 6871 4063
rect 12633 3961 12667 3995
rect 4997 3893 5031 3927
rect 6469 3893 6503 3927
rect 17969 3893 18003 3927
rect 1593 3689 1627 3723
rect 4353 3689 4387 3723
rect 9045 3689 9079 3723
rect 12173 3689 12207 3723
rect 8769 3621 8803 3655
rect 10517 3621 10551 3655
rect 1961 3553 1995 3587
rect 2421 3553 2455 3587
rect 4169 3553 4203 3587
rect 4721 3553 4755 3587
rect 8493 3553 8527 3587
rect 9689 3553 9723 3587
rect 10333 3553 10367 3587
rect 11989 3553 12023 3587
rect 17785 3553 17819 3587
rect 1409 3485 1443 3519
rect 1685 3485 1719 3519
rect 2053 3485 2087 3519
rect 2513 3485 2547 3519
rect 2697 3485 2731 3519
rect 2881 3485 2915 3519
rect 3893 3485 3927 3519
rect 3985 3485 4019 3519
rect 4077 3485 4111 3519
rect 4813 3485 4847 3519
rect 7941 3485 7975 3519
rect 8125 3485 8159 3519
rect 8401 3485 8435 3519
rect 8953 3485 8987 3519
rect 9229 3485 9263 3519
rect 9597 3485 9631 3519
rect 9781 3485 9815 3519
rect 9965 3485 9999 3519
rect 10241 3485 10275 3519
rect 12357 3485 12391 3519
rect 12449 3485 12483 3519
rect 17509 3485 17543 3519
rect 18061 3485 18095 3519
rect 3249 3417 3283 3451
rect 3433 3417 3467 3451
rect 8033 3417 8067 3451
rect 9873 3417 9907 3451
rect 18337 3417 18371 3451
rect 3617 3349 3651 3383
rect 4445 3349 4479 3383
rect 9505 3349 9539 3383
rect 2145 3145 2179 3179
rect 2605 3145 2639 3179
rect 5365 3145 5399 3179
rect 7757 3145 7791 3179
rect 9965 3145 9999 3179
rect 10793 3145 10827 3179
rect 10885 3145 10919 3179
rect 11897 3145 11931 3179
rect 11989 3145 12023 3179
rect 12725 3145 12759 3179
rect 13553 3145 13587 3179
rect 2513 3077 2547 3111
rect 5273 3077 5307 3111
rect 8217 3077 8251 3111
rect 12817 3077 12851 3111
rect 13645 3077 13679 3111
rect 2053 3009 2087 3043
rect 3433 3009 3467 3043
rect 4169 3009 4203 3043
rect 4445 3009 4479 3043
rect 6469 3009 6503 3043
rect 7389 3009 7423 3043
rect 8033 3009 8067 3043
rect 8401 3009 8435 3043
rect 8677 3009 8711 3043
rect 8861 3009 8895 3043
rect 10057 3009 10091 3043
rect 17509 3009 17543 3043
rect 18521 3009 18555 3043
rect 1869 2941 1903 2975
rect 2697 2941 2731 2975
rect 3157 2941 3191 2975
rect 3893 2941 3927 2975
rect 4629 2941 4663 2975
rect 5457 2941 5491 2975
rect 6653 2941 6687 2975
rect 7481 2941 7515 2975
rect 8493 2941 8527 2975
rect 9873 2941 9907 2975
rect 10609 2941 10643 2975
rect 12081 2941 12115 2975
rect 13001 2941 13035 2975
rect 13737 2941 13771 2975
rect 17693 2941 17727 2975
rect 18245 2941 18279 2975
rect 4905 2873 4939 2907
rect 13185 2873 13219 2907
rect 4261 2805 4295 2839
rect 10425 2805 10459 2839
rect 11253 2805 11287 2839
rect 11529 2805 11563 2839
rect 12357 2805 12391 2839
rect 1593 2601 1627 2635
rect 1869 2601 1903 2635
rect 2881 2601 2915 2635
rect 3893 2601 3927 2635
rect 2329 2465 2363 2499
rect 2513 2465 2547 2499
rect 15393 2465 15427 2499
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 2697 2397 2731 2431
rect 3617 2397 3651 2431
rect 3801 2397 3835 2431
rect 3985 2397 4019 2431
rect 4537 2397 4571 2431
rect 5089 2397 5123 2431
rect 5641 2397 5675 2431
rect 5733 2397 5767 2431
rect 6653 2397 6687 2431
rect 7665 2397 7699 2431
rect 8217 2397 8251 2431
rect 8769 2397 8803 2431
rect 9689 2397 9723 2431
rect 10241 2397 10275 2431
rect 10333 2397 10367 2431
rect 11345 2397 11379 2431
rect 11529 2397 11563 2431
rect 12541 2397 12575 2431
rect 12633 2397 12667 2431
rect 13645 2397 13679 2431
rect 14105 2397 14139 2431
rect 14657 2397 14691 2431
rect 15209 2397 15243 2431
rect 16221 2397 16255 2431
rect 16681 2397 16715 2431
rect 16957 2397 16991 2431
rect 17233 2397 17267 2431
rect 17785 2397 17819 2431
rect 2973 2329 3007 2363
rect 3341 2329 3375 2363
rect 4261 2329 4295 2363
rect 4813 2329 4847 2363
rect 5365 2329 5399 2363
rect 6009 2329 6043 2363
rect 6929 2329 6963 2363
rect 7389 2329 7423 2363
rect 7941 2329 7975 2363
rect 8493 2329 8527 2363
rect 9413 2329 9447 2363
rect 9965 2329 9999 2363
rect 10609 2329 10643 2363
rect 11069 2329 11103 2363
rect 11805 2329 11839 2363
rect 12265 2329 12299 2363
rect 12909 2329 12943 2363
rect 13369 2329 13403 2363
rect 14381 2329 14415 2363
rect 14933 2329 14967 2363
rect 15945 2329 15979 2363
rect 17509 2329 17543 2363
rect 18061 2329 18095 2363
rect 2237 2261 2271 2295
<< metal1 >>
rect 7006 17688 7012 17740
rect 7064 17728 7070 17740
rect 15010 17728 15016 17740
rect 7064 17700 15016 17728
rect 7064 17688 7070 17700
rect 15010 17688 15016 17700
rect 15068 17688 15074 17740
rect 12250 17552 12256 17604
rect 12308 17592 12314 17604
rect 16758 17592 16764 17604
rect 12308 17564 16764 17592
rect 12308 17552 12314 17564
rect 16758 17552 16764 17564
rect 16816 17552 16822 17604
rect 7742 17484 7748 17536
rect 7800 17524 7806 17536
rect 15378 17524 15384 17536
rect 7800 17496 15384 17524
rect 7800 17484 7806 17496
rect 15378 17484 15384 17496
rect 15436 17484 15442 17536
rect 15746 17484 15752 17536
rect 15804 17524 15810 17536
rect 16482 17524 16488 17536
rect 15804 17496 16488 17524
rect 15804 17484 15810 17496
rect 16482 17484 16488 17496
rect 16540 17484 16546 17536
rect 1104 17434 18860 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 18860 17434
rect 1104 17360 18860 17382
rect 2498 17280 2504 17332
rect 2556 17280 2562 17332
rect 3050 17280 3056 17332
rect 3108 17280 3114 17332
rect 3602 17280 3608 17332
rect 3660 17320 3666 17332
rect 5997 17323 6055 17329
rect 5997 17320 6009 17323
rect 3660 17292 3924 17320
rect 3660 17280 3666 17292
rect 1946 17212 1952 17264
rect 2004 17252 2010 17264
rect 2133 17255 2191 17261
rect 2133 17252 2145 17255
rect 2004 17224 2145 17252
rect 2004 17212 2010 17224
rect 2133 17221 2145 17224
rect 2179 17221 2191 17255
rect 2133 17215 2191 17221
rect 1486 17144 1492 17196
rect 1544 17144 1550 17196
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17153 1823 17187
rect 2516 17184 2544 17280
rect 2593 17187 2651 17193
rect 2593 17184 2605 17187
rect 2516 17156 2605 17184
rect 1765 17147 1823 17153
rect 2593 17153 2605 17156
rect 2639 17153 2651 17187
rect 3068 17184 3096 17280
rect 3896 17261 3924 17292
rect 4080 17292 6009 17320
rect 3881 17255 3939 17261
rect 3881 17221 3893 17255
rect 3927 17221 3939 17255
rect 3881 17215 3939 17221
rect 3145 17187 3203 17193
rect 3145 17184 3157 17187
rect 3068 17156 3157 17184
rect 2593 17147 2651 17153
rect 3145 17153 3157 17156
rect 3191 17153 3203 17187
rect 3145 17147 3203 17153
rect 1302 17076 1308 17128
rect 1360 17116 1366 17128
rect 1780 17116 1808 17147
rect 3418 17144 3424 17196
rect 3476 17184 3482 17196
rect 4080 17184 4108 17292
rect 5997 17289 6009 17292
rect 6043 17289 6055 17323
rect 5997 17283 6055 17289
rect 6730 17280 6736 17332
rect 6788 17320 6794 17332
rect 7006 17320 7012 17332
rect 6788 17292 7012 17320
rect 6788 17280 6794 17292
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 7466 17280 7472 17332
rect 7524 17280 7530 17332
rect 8018 17280 8024 17332
rect 8076 17320 8082 17332
rect 8076 17292 8248 17320
rect 8076 17280 8082 17292
rect 4154 17212 4160 17264
rect 4212 17252 4218 17264
rect 4341 17255 4399 17261
rect 4341 17252 4353 17255
rect 4212 17224 4353 17252
rect 4212 17212 4218 17224
rect 4341 17221 4353 17224
rect 4387 17221 4399 17255
rect 4341 17215 4399 17221
rect 4617 17255 4675 17261
rect 4617 17221 4629 17255
rect 4663 17252 4675 17255
rect 5813 17255 5871 17261
rect 4663 17224 5304 17252
rect 4663 17221 4675 17224
rect 4617 17215 4675 17221
rect 5276 17196 5304 17224
rect 5813 17221 5825 17255
rect 5859 17252 5871 17255
rect 6362 17252 6368 17264
rect 5859 17224 6368 17252
rect 5859 17221 5871 17224
rect 5813 17215 5871 17221
rect 6362 17212 6368 17224
rect 6420 17252 6426 17264
rect 6641 17255 6699 17261
rect 6641 17252 6653 17255
rect 6420 17224 6653 17252
rect 6420 17212 6426 17224
rect 6641 17221 6653 17224
rect 6687 17221 6699 17255
rect 6641 17215 6699 17221
rect 6914 17212 6920 17264
rect 6972 17252 6978 17264
rect 6972 17224 7144 17252
rect 6972 17212 6978 17224
rect 3476 17156 4108 17184
rect 3476 17144 3482 17156
rect 4706 17144 4712 17196
rect 4764 17184 4770 17196
rect 4801 17187 4859 17193
rect 4801 17184 4813 17187
rect 4764 17156 4813 17184
rect 4764 17144 4770 17156
rect 4801 17153 4813 17156
rect 4847 17153 4859 17187
rect 4801 17147 4859 17153
rect 5258 17144 5264 17196
rect 5316 17184 5322 17196
rect 5353 17187 5411 17193
rect 5353 17184 5365 17187
rect 5316 17156 5365 17184
rect 5316 17144 5322 17156
rect 5353 17153 5365 17156
rect 5399 17153 5411 17187
rect 5353 17147 5411 17153
rect 5902 17144 5908 17196
rect 5960 17184 5966 17196
rect 6089 17187 6147 17193
rect 6089 17184 6101 17187
rect 5960 17156 6101 17184
rect 5960 17144 5966 17156
rect 6089 17153 6101 17156
rect 6135 17153 6147 17187
rect 6546 17184 6552 17196
rect 6089 17147 6147 17153
rect 6196 17156 6552 17184
rect 5169 17119 5227 17125
rect 1360 17088 1808 17116
rect 1964 17088 5120 17116
rect 1360 17076 1366 17088
rect 1964 17057 1992 17088
rect 1949 17051 2007 17057
rect 1949 17017 1961 17051
rect 1995 17017 2007 17051
rect 1949 17011 2007 17017
rect 2777 17051 2835 17057
rect 2777 17017 2789 17051
rect 2823 17048 2835 17051
rect 4525 17051 4583 17057
rect 2823 17020 4476 17048
rect 2823 17017 2835 17020
rect 2777 17011 2835 17017
rect 1670 16940 1676 16992
rect 1728 16940 1734 16992
rect 2038 16940 2044 16992
rect 2096 16980 2102 16992
rect 2225 16983 2283 16989
rect 2225 16980 2237 16983
rect 2096 16952 2237 16980
rect 2096 16940 2102 16952
rect 2225 16949 2237 16952
rect 2271 16949 2283 16983
rect 2225 16943 2283 16949
rect 3329 16983 3387 16989
rect 3329 16949 3341 16983
rect 3375 16980 3387 16983
rect 3510 16980 3516 16992
rect 3375 16952 3516 16980
rect 3375 16949 3387 16952
rect 3329 16943 3387 16949
rect 3510 16940 3516 16952
rect 3568 16940 3574 16992
rect 3878 16940 3884 16992
rect 3936 16980 3942 16992
rect 3973 16983 4031 16989
rect 3973 16980 3985 16983
rect 3936 16952 3985 16980
rect 3936 16940 3942 16952
rect 3973 16949 3985 16952
rect 4019 16949 4031 16983
rect 4448 16980 4476 17020
rect 4525 17017 4537 17051
rect 4571 17048 4583 17051
rect 4614 17048 4620 17060
rect 4571 17020 4620 17048
rect 4571 17017 4583 17020
rect 4525 17011 4583 17017
rect 4614 17008 4620 17020
rect 4672 17008 4678 17060
rect 5092 17048 5120 17088
rect 5169 17085 5181 17119
rect 5215 17116 5227 17119
rect 5920 17116 5948 17144
rect 5215 17088 5948 17116
rect 5215 17085 5227 17088
rect 5169 17079 5227 17085
rect 6196 17048 6224 17156
rect 6546 17144 6552 17156
rect 6604 17184 6610 17196
rect 6825 17187 6883 17193
rect 6825 17184 6837 17187
rect 6604 17156 6837 17184
rect 6604 17144 6610 17156
rect 6825 17153 6837 17156
rect 6871 17153 6883 17187
rect 6825 17147 6883 17153
rect 7006 17144 7012 17196
rect 7064 17144 7070 17196
rect 7116 17193 7144 17224
rect 7101 17187 7159 17193
rect 7101 17153 7113 17187
rect 7147 17153 7159 17187
rect 7484 17184 7512 17280
rect 8220 17261 8248 17292
rect 8570 17280 8576 17332
rect 8628 17280 8634 17332
rect 9674 17280 9680 17332
rect 9732 17280 9738 17332
rect 10226 17280 10232 17332
rect 10284 17320 10290 17332
rect 10284 17292 10456 17320
rect 10284 17280 10290 17292
rect 8205 17255 8263 17261
rect 8205 17221 8217 17255
rect 8251 17221 8263 17255
rect 8205 17215 8263 17221
rect 7561 17187 7619 17193
rect 7561 17184 7573 17187
rect 7484 17156 7573 17184
rect 7101 17147 7159 17153
rect 7561 17153 7573 17156
rect 7607 17153 7619 17187
rect 8588 17184 8616 17280
rect 8757 17255 8815 17261
rect 8757 17221 8769 17255
rect 8803 17252 8815 17255
rect 8803 17224 9168 17252
rect 8803 17221 8815 17224
rect 8757 17215 8815 17221
rect 9140 17196 9168 17224
rect 8941 17187 8999 17193
rect 8941 17184 8953 17187
rect 8588 17156 8953 17184
rect 7561 17147 7619 17153
rect 8941 17153 8953 17156
rect 8987 17153 8999 17187
rect 8941 17147 8999 17153
rect 9122 17144 9128 17196
rect 9180 17184 9186 17196
rect 9217 17187 9275 17193
rect 9217 17184 9229 17187
rect 9180 17156 9229 17184
rect 9180 17144 9186 17156
rect 9217 17153 9229 17156
rect 9263 17153 9275 17187
rect 9692 17184 9720 17280
rect 10428 17261 10456 17292
rect 10778 17280 10784 17332
rect 10836 17320 10842 17332
rect 11057 17323 11115 17329
rect 11057 17320 11069 17323
rect 10836 17292 11069 17320
rect 10836 17280 10842 17292
rect 11057 17289 11069 17292
rect 11103 17289 11115 17323
rect 11057 17283 11115 17289
rect 10413 17255 10471 17261
rect 10413 17221 10425 17255
rect 10459 17221 10471 17255
rect 11072 17252 11100 17283
rect 12986 17280 12992 17332
rect 13044 17320 13050 17332
rect 13998 17320 14004 17332
rect 13044 17292 14004 17320
rect 13044 17280 13050 17292
rect 13998 17280 14004 17292
rect 14056 17280 14062 17332
rect 15194 17280 15200 17332
rect 15252 17320 15258 17332
rect 16022 17320 16028 17332
rect 15252 17292 16028 17320
rect 15252 17280 15258 17292
rect 16022 17280 16028 17292
rect 16080 17320 16086 17332
rect 16393 17323 16451 17329
rect 16393 17320 16405 17323
rect 16080 17292 16405 17320
rect 16080 17280 16086 17292
rect 16393 17289 16405 17292
rect 16439 17289 16451 17323
rect 16393 17283 16451 17289
rect 16850 17280 16856 17332
rect 16908 17320 16914 17332
rect 16908 17292 17264 17320
rect 16908 17280 16914 17292
rect 15473 17255 15531 17261
rect 15473 17252 15485 17255
rect 11072 17224 11560 17252
rect 10413 17215 10471 17221
rect 9769 17187 9827 17193
rect 9769 17184 9781 17187
rect 9692 17156 9781 17184
rect 9217 17147 9275 17153
rect 9769 17153 9781 17156
rect 9815 17153 9827 17187
rect 9769 17147 9827 17153
rect 10873 17187 10931 17193
rect 10873 17153 10885 17187
rect 10919 17184 10931 17187
rect 11149 17187 11207 17193
rect 11149 17184 11161 17187
rect 10919 17156 11161 17184
rect 10919 17153 10931 17156
rect 10873 17147 10931 17153
rect 11149 17153 11161 17156
rect 11195 17184 11207 17187
rect 11330 17184 11336 17196
rect 11195 17156 11336 17184
rect 11195 17153 11207 17156
rect 11149 17147 11207 17153
rect 11330 17144 11336 17156
rect 11388 17144 11394 17196
rect 11532 17193 11560 17224
rect 14200 17224 15485 17252
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17153 11575 17187
rect 11517 17147 11575 17153
rect 12434 17144 12440 17196
rect 12492 17184 12498 17196
rect 12529 17187 12587 17193
rect 12529 17184 12541 17187
rect 12492 17156 12541 17184
rect 12492 17144 12498 17156
rect 12529 17153 12541 17156
rect 12575 17153 12587 17187
rect 13262 17184 13268 17196
rect 12529 17147 12587 17153
rect 12912 17156 13268 17184
rect 6638 17076 6644 17128
rect 6696 17116 6702 17128
rect 11698 17116 11704 17128
rect 6696 17088 11704 17116
rect 6696 17076 6702 17088
rect 11698 17076 11704 17088
rect 11756 17076 11762 17128
rect 11790 17076 11796 17128
rect 11848 17076 11854 17128
rect 12802 17076 12808 17128
rect 12860 17076 12866 17128
rect 5092 17020 6224 17048
rect 6270 17008 6276 17060
rect 6328 17048 6334 17060
rect 6457 17051 6515 17057
rect 6457 17048 6469 17051
rect 6328 17020 6469 17048
rect 6328 17008 6334 17020
rect 6457 17017 6469 17020
rect 6503 17017 6515 17051
rect 6457 17011 6515 17017
rect 8389 17051 8447 17057
rect 8389 17017 8401 17051
rect 8435 17048 8447 17051
rect 10042 17048 10048 17060
rect 8435 17020 10048 17048
rect 8435 17017 8447 17020
rect 8389 17011 8447 17017
rect 10042 17008 10048 17020
rect 10100 17008 10106 17060
rect 10597 17051 10655 17057
rect 10597 17017 10609 17051
rect 10643 17048 10655 17051
rect 10686 17048 10692 17060
rect 10643 17020 10692 17048
rect 10643 17017 10655 17020
rect 10597 17011 10655 17017
rect 10686 17008 10692 17020
rect 10744 17008 10750 17060
rect 11882 17008 11888 17060
rect 11940 17048 11946 17060
rect 12912 17048 12940 17156
rect 13262 17144 13268 17156
rect 13320 17184 13326 17196
rect 13633 17187 13691 17193
rect 13633 17184 13645 17187
rect 13320 17156 13645 17184
rect 13320 17144 13326 17156
rect 13633 17153 13645 17156
rect 13679 17153 13691 17187
rect 13633 17147 13691 17153
rect 13734 17191 13792 17197
rect 13734 17157 13746 17191
rect 13780 17184 13792 17191
rect 13906 17184 13912 17196
rect 13780 17157 13912 17184
rect 13734 17156 13912 17157
rect 13734 17151 13792 17156
rect 13906 17144 13912 17156
rect 13964 17144 13970 17196
rect 14090 17144 14096 17196
rect 14148 17184 14154 17196
rect 14200 17193 14228 17224
rect 15473 17221 15485 17224
rect 15519 17221 15531 17255
rect 15473 17215 15531 17221
rect 15764 17224 16436 17252
rect 15764 17196 15792 17224
rect 14185 17187 14243 17193
rect 14185 17184 14197 17187
rect 14148 17156 14197 17184
rect 14148 17144 14154 17156
rect 14185 17153 14197 17156
rect 14231 17153 14243 17187
rect 14185 17147 14243 17153
rect 14642 17144 14648 17196
rect 14700 17184 14706 17196
rect 15102 17184 15108 17196
rect 14700 17156 15108 17184
rect 14700 17144 14706 17156
rect 15102 17144 15108 17156
rect 15160 17184 15166 17196
rect 15289 17187 15347 17193
rect 15289 17184 15301 17187
rect 15160 17156 15301 17184
rect 15160 17144 15166 17156
rect 15289 17153 15301 17156
rect 15335 17153 15347 17187
rect 15289 17147 15347 17153
rect 15654 17144 15660 17196
rect 15712 17144 15718 17196
rect 15746 17144 15752 17196
rect 15804 17144 15810 17196
rect 15930 17144 15936 17196
rect 15988 17144 15994 17196
rect 16022 17144 16028 17196
rect 16080 17184 16086 17196
rect 16294 17188 16352 17193
rect 16224 17187 16352 17188
rect 16224 17184 16306 17187
rect 16080 17160 16306 17184
rect 16080 17156 16252 17160
rect 16080 17144 16086 17156
rect 16294 17153 16306 17160
rect 16340 17153 16352 17187
rect 16408 17184 16436 17224
rect 16482 17212 16488 17264
rect 16540 17252 16546 17264
rect 17236 17261 17264 17292
rect 17221 17255 17279 17261
rect 16540 17224 16988 17252
rect 16540 17212 16546 17224
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 16408 17156 16681 17184
rect 16294 17147 16352 17153
rect 16669 17153 16681 17156
rect 16715 17153 16727 17187
rect 16669 17147 16727 17153
rect 16758 17144 16764 17196
rect 16816 17184 16822 17196
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 16816 17156 16865 17184
rect 16816 17144 16822 17156
rect 16853 17153 16865 17156
rect 16899 17153 16911 17187
rect 16960 17184 16988 17224
rect 17221 17221 17233 17255
rect 17267 17221 17279 17255
rect 17221 17215 17279 17221
rect 17589 17187 17647 17193
rect 17589 17184 17601 17187
rect 16960 17156 17601 17184
rect 16853 17147 16911 17153
rect 17589 17153 17601 17156
rect 17635 17153 17647 17187
rect 17589 17147 17647 17153
rect 18506 17144 18512 17196
rect 18564 17144 18570 17196
rect 14458 17076 14464 17128
rect 14516 17076 14522 17128
rect 16206 17076 16212 17128
rect 16264 17116 16270 17128
rect 18233 17119 18291 17125
rect 18233 17116 18245 17119
rect 16264 17088 18245 17116
rect 16264 17076 16270 17088
rect 18233 17085 18245 17088
rect 18279 17085 18291 17119
rect 18233 17079 18291 17085
rect 11940 17020 12940 17048
rect 11940 17008 11946 17020
rect 15010 17008 15016 17060
rect 15068 17048 15074 17060
rect 15105 17051 15163 17057
rect 15105 17048 15117 17051
rect 15068 17020 15117 17048
rect 15068 17008 15074 17020
rect 15105 17017 15117 17020
rect 15151 17017 15163 17051
rect 15105 17011 15163 17017
rect 15286 17008 15292 17060
rect 15344 17048 15350 17060
rect 17037 17051 17095 17057
rect 17037 17048 17049 17051
rect 15344 17020 17049 17048
rect 15344 17008 15350 17020
rect 17037 17017 17049 17020
rect 17083 17017 17095 17051
rect 17037 17011 17095 17017
rect 4798 16980 4804 16992
rect 4448 16952 4804 16980
rect 3973 16943 4031 16949
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 4985 16983 5043 16989
rect 4985 16949 4997 16983
rect 5031 16980 5043 16983
rect 5350 16980 5356 16992
rect 5031 16952 5356 16980
rect 5031 16949 5043 16952
rect 4985 16943 5043 16949
rect 5350 16940 5356 16952
rect 5408 16940 5414 16992
rect 5537 16983 5595 16989
rect 5537 16949 5549 16983
rect 5583 16980 5595 16983
rect 5902 16980 5908 16992
rect 5583 16952 5908 16980
rect 5583 16949 5595 16952
rect 5537 16943 5595 16949
rect 5902 16940 5908 16952
rect 5960 16940 5966 16992
rect 6914 16940 6920 16992
rect 6972 16940 6978 16992
rect 7285 16983 7343 16989
rect 7285 16949 7297 16983
rect 7331 16980 7343 16983
rect 7558 16980 7564 16992
rect 7331 16952 7564 16980
rect 7331 16949 7343 16952
rect 7285 16943 7343 16949
rect 7558 16940 7564 16952
rect 7616 16940 7622 16992
rect 7745 16983 7803 16989
rect 7745 16949 7757 16983
rect 7791 16980 7803 16983
rect 7926 16980 7932 16992
rect 7791 16952 7932 16980
rect 7791 16949 7803 16952
rect 7745 16943 7803 16949
rect 7926 16940 7932 16952
rect 7984 16940 7990 16992
rect 9030 16940 9036 16992
rect 9088 16980 9094 16992
rect 9125 16983 9183 16989
rect 9125 16980 9137 16983
rect 9088 16952 9137 16980
rect 9088 16940 9094 16952
rect 9125 16949 9137 16952
rect 9171 16949 9183 16983
rect 9125 16943 9183 16949
rect 9401 16983 9459 16989
rect 9401 16949 9413 16983
rect 9447 16980 9459 16983
rect 9582 16980 9588 16992
rect 9447 16952 9588 16980
rect 9447 16949 9459 16952
rect 9401 16943 9459 16949
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 9953 16983 10011 16989
rect 9953 16949 9965 16983
rect 9999 16980 10011 16983
rect 10226 16980 10232 16992
rect 9999 16952 10232 16980
rect 9999 16949 10011 16952
rect 9953 16943 10011 16949
rect 10226 16940 10232 16952
rect 10284 16940 10290 16992
rect 11330 16940 11336 16992
rect 11388 16940 11394 16992
rect 12894 16940 12900 16992
rect 12952 16980 12958 16992
rect 13449 16983 13507 16989
rect 13449 16980 13461 16983
rect 12952 16952 13461 16980
rect 12952 16940 12958 16952
rect 13449 16949 13461 16952
rect 13495 16949 13507 16983
rect 13449 16943 13507 16949
rect 13906 16940 13912 16992
rect 13964 16940 13970 16992
rect 14642 16940 14648 16992
rect 14700 16980 14706 16992
rect 15562 16980 15568 16992
rect 14700 16952 15568 16980
rect 14700 16940 14706 16952
rect 15562 16940 15568 16952
rect 15620 16940 15626 16992
rect 15933 16983 15991 16989
rect 15933 16949 15945 16983
rect 15979 16980 15991 16983
rect 16022 16980 16028 16992
rect 15979 16952 16028 16980
rect 15979 16949 15991 16952
rect 15933 16943 15991 16949
rect 16022 16940 16028 16952
rect 16080 16940 16086 16992
rect 16114 16940 16120 16992
rect 16172 16940 16178 16992
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 17405 16983 17463 16989
rect 17405 16980 17417 16983
rect 16724 16952 17417 16980
rect 16724 16940 16730 16952
rect 17405 16949 17417 16952
rect 17451 16949 17463 16983
rect 17405 16943 17463 16949
rect 1104 16890 18860 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 18860 16890
rect 1104 16816 18860 16838
rect 1946 16736 1952 16788
rect 2004 16736 2010 16788
rect 4154 16736 4160 16788
rect 4212 16736 4218 16788
rect 4706 16736 4712 16788
rect 4764 16736 4770 16788
rect 6549 16779 6607 16785
rect 6549 16745 6561 16779
rect 6595 16776 6607 16779
rect 7006 16776 7012 16788
rect 6595 16748 7012 16776
rect 6595 16745 6607 16748
rect 6549 16739 6607 16745
rect 7006 16736 7012 16748
rect 7064 16736 7070 16788
rect 12250 16736 12256 16788
rect 12308 16736 12314 16788
rect 12710 16776 12716 16788
rect 12406 16748 12716 16776
rect 1670 16668 1676 16720
rect 1728 16708 1734 16720
rect 2041 16711 2099 16717
rect 2041 16708 2053 16711
rect 1728 16680 2053 16708
rect 1728 16668 1734 16680
rect 2041 16677 2053 16680
rect 2087 16677 2099 16711
rect 2041 16671 2099 16677
rect 8496 16680 8892 16708
rect 1302 16600 1308 16652
rect 1360 16640 1366 16652
rect 2225 16643 2283 16649
rect 2225 16640 2237 16643
rect 1360 16612 2237 16640
rect 1360 16600 1366 16612
rect 2225 16609 2237 16612
rect 2271 16609 2283 16643
rect 2225 16603 2283 16609
rect 6365 16643 6423 16649
rect 6365 16609 6377 16643
rect 6411 16640 6423 16643
rect 6825 16643 6883 16649
rect 6411 16612 6776 16640
rect 6411 16609 6423 16612
rect 6365 16603 6423 16609
rect 1394 16532 1400 16584
rect 1452 16572 1458 16584
rect 1673 16575 1731 16581
rect 1673 16572 1685 16575
rect 1452 16544 1685 16572
rect 1452 16532 1458 16544
rect 1673 16541 1685 16544
rect 1719 16541 1731 16575
rect 1673 16535 1731 16541
rect 5537 16575 5595 16581
rect 5537 16541 5549 16575
rect 5583 16541 5595 16575
rect 5537 16535 5595 16541
rect 5552 16504 5580 16535
rect 5810 16532 5816 16584
rect 5868 16572 5874 16584
rect 5997 16575 6055 16581
rect 5997 16572 6009 16575
rect 5868 16544 6009 16572
rect 5868 16532 5874 16544
rect 5997 16541 6009 16544
rect 6043 16572 6055 16575
rect 6638 16572 6644 16584
rect 6043 16544 6644 16572
rect 6043 16541 6055 16544
rect 5997 16535 6055 16541
rect 6638 16532 6644 16544
rect 6696 16532 6702 16584
rect 6748 16572 6776 16612
rect 6825 16609 6837 16643
rect 6871 16640 6883 16643
rect 6914 16640 6920 16652
rect 6871 16612 6920 16640
rect 6871 16609 6883 16612
rect 6825 16603 6883 16609
rect 6914 16600 6920 16612
rect 6972 16600 6978 16652
rect 7742 16600 7748 16652
rect 7800 16600 7806 16652
rect 8496 16649 8524 16680
rect 8481 16643 8539 16649
rect 8481 16609 8493 16643
rect 8527 16609 8539 16643
rect 8481 16603 8539 16609
rect 8754 16600 8760 16652
rect 8812 16600 8818 16652
rect 8864 16640 8892 16680
rect 9214 16668 9220 16720
rect 9272 16708 9278 16720
rect 9861 16711 9919 16717
rect 9861 16708 9873 16711
rect 9272 16680 9873 16708
rect 9272 16668 9278 16680
rect 9861 16677 9873 16680
rect 9907 16677 9919 16711
rect 9861 16671 9919 16677
rect 12069 16711 12127 16717
rect 12069 16677 12081 16711
rect 12115 16708 12127 16711
rect 12406 16708 12434 16748
rect 12710 16736 12716 16748
rect 12768 16776 12774 16788
rect 12768 16748 13676 16776
rect 12768 16736 12774 16748
rect 12115 16680 12434 16708
rect 13265 16711 13323 16717
rect 12115 16677 12127 16680
rect 12069 16671 12127 16677
rect 13265 16677 13277 16711
rect 13311 16677 13323 16711
rect 13265 16671 13323 16677
rect 9493 16643 9551 16649
rect 9493 16640 9505 16643
rect 8864 16612 9505 16640
rect 9493 16609 9505 16612
rect 9539 16640 9551 16643
rect 9950 16640 9956 16652
rect 9539 16612 9956 16640
rect 9539 16609 9551 16612
rect 9493 16603 9551 16609
rect 9950 16600 9956 16612
rect 10008 16640 10014 16652
rect 10008 16612 10272 16640
rect 10008 16600 10014 16612
rect 7006 16572 7012 16584
rect 6748 16544 7012 16572
rect 7006 16532 7012 16544
rect 7064 16532 7070 16584
rect 7466 16532 7472 16584
rect 7524 16532 7530 16584
rect 8389 16575 8447 16581
rect 8389 16541 8401 16575
rect 8435 16572 8447 16575
rect 9401 16575 9459 16581
rect 9401 16572 9413 16575
rect 8435 16544 9413 16572
rect 8435 16541 8447 16544
rect 8389 16535 8447 16541
rect 9401 16541 9413 16544
rect 9447 16572 9459 16575
rect 10244 16572 10272 16612
rect 11054 16600 11060 16652
rect 11112 16640 11118 16652
rect 11425 16643 11483 16649
rect 11425 16640 11437 16643
rect 11112 16612 11437 16640
rect 11112 16600 11118 16612
rect 11425 16609 11437 16612
rect 11471 16609 11483 16643
rect 12526 16640 12532 16652
rect 11425 16603 11483 16609
rect 11624 16612 11836 16640
rect 11624 16572 11652 16612
rect 9447 16544 10180 16572
rect 10244 16544 11652 16572
rect 9447 16541 9459 16544
rect 9401 16535 9459 16541
rect 5626 16504 5632 16516
rect 1596 16476 5632 16504
rect 1596 16445 1624 16476
rect 5626 16464 5632 16476
rect 5684 16464 5690 16516
rect 10045 16507 10103 16513
rect 10045 16473 10057 16507
rect 10091 16473 10103 16507
rect 10152 16504 10180 16544
rect 11698 16532 11704 16584
rect 11756 16532 11762 16584
rect 11808 16572 11836 16612
rect 11992 16612 12532 16640
rect 11882 16572 11888 16584
rect 11808 16544 11888 16572
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 11992 16581 12020 16612
rect 12526 16600 12532 16612
rect 12584 16600 12590 16652
rect 11977 16575 12035 16581
rect 11977 16541 11989 16575
rect 12023 16541 12035 16575
rect 11977 16535 12035 16541
rect 12158 16532 12164 16584
rect 12216 16572 12222 16584
rect 12989 16575 13047 16581
rect 12989 16572 13001 16575
rect 12216 16544 13001 16572
rect 12216 16532 12222 16544
rect 12989 16541 13001 16544
rect 13035 16541 13047 16575
rect 13280 16572 13308 16671
rect 13648 16649 13676 16748
rect 14642 16736 14648 16788
rect 14700 16736 14706 16788
rect 15286 16776 15292 16788
rect 14936 16748 15292 16776
rect 14936 16717 14964 16748
rect 15286 16736 15292 16748
rect 15344 16736 15350 16788
rect 15473 16779 15531 16785
rect 15473 16745 15485 16779
rect 15519 16776 15531 16779
rect 15654 16776 15660 16788
rect 15519 16748 15660 16776
rect 15519 16745 15531 16748
rect 15473 16739 15531 16745
rect 15654 16736 15660 16748
rect 15712 16736 15718 16788
rect 16758 16736 16764 16788
rect 16816 16776 16822 16788
rect 17497 16779 17555 16785
rect 17497 16776 17509 16779
rect 16816 16748 17509 16776
rect 16816 16736 16822 16748
rect 17497 16745 17509 16748
rect 17543 16745 17555 16779
rect 17497 16739 17555 16745
rect 14921 16711 14979 16717
rect 14921 16677 14933 16711
rect 14967 16677 14979 16711
rect 14921 16671 14979 16677
rect 15102 16668 15108 16720
rect 15160 16708 15166 16720
rect 15565 16711 15623 16717
rect 15565 16708 15577 16711
rect 15160 16680 15577 16708
rect 15160 16668 15166 16680
rect 15565 16677 15577 16680
rect 15611 16677 15623 16711
rect 16206 16708 16212 16720
rect 15565 16671 15623 16677
rect 15856 16680 16212 16708
rect 13633 16643 13691 16649
rect 13633 16609 13645 16643
rect 13679 16609 13691 16643
rect 15856 16640 15884 16680
rect 16206 16668 16212 16680
rect 16264 16668 16270 16720
rect 17129 16711 17187 16717
rect 17129 16677 17141 16711
rect 17175 16708 17187 16711
rect 18046 16708 18052 16720
rect 17175 16680 18052 16708
rect 17175 16677 17187 16680
rect 17129 16671 17187 16677
rect 18046 16668 18052 16680
rect 18104 16668 18110 16720
rect 13633 16603 13691 16609
rect 14200 16612 14504 16640
rect 12989 16535 13047 16541
rect 13096 16544 13308 16572
rect 13725 16575 13783 16581
rect 12342 16504 12348 16516
rect 10152 16476 12348 16504
rect 10045 16467 10103 16473
rect 1581 16439 1639 16445
rect 1581 16405 1593 16439
rect 1627 16405 1639 16439
rect 1581 16399 1639 16405
rect 9766 16396 9772 16448
rect 9824 16396 9830 16448
rect 10060 16436 10088 16467
rect 12342 16464 12348 16476
rect 12400 16464 12406 16516
rect 12437 16507 12495 16513
rect 12437 16473 12449 16507
rect 12483 16473 12495 16507
rect 12437 16467 12495 16473
rect 10870 16436 10876 16448
rect 10060 16408 10876 16436
rect 10870 16396 10876 16408
rect 10928 16396 10934 16448
rect 11238 16396 11244 16448
rect 11296 16436 11302 16448
rect 11885 16439 11943 16445
rect 11885 16436 11897 16439
rect 11296 16408 11897 16436
rect 11296 16396 11302 16408
rect 11885 16405 11897 16408
rect 11931 16405 11943 16439
rect 11885 16399 11943 16405
rect 11974 16396 11980 16448
rect 12032 16436 12038 16448
rect 12227 16439 12285 16445
rect 12227 16436 12239 16439
rect 12032 16408 12239 16436
rect 12032 16396 12038 16408
rect 12227 16405 12239 16408
rect 12273 16405 12285 16439
rect 12452 16436 12480 16467
rect 12710 16464 12716 16516
rect 12768 16464 12774 16516
rect 12897 16507 12955 16513
rect 12897 16473 12909 16507
rect 12943 16504 12955 16507
rect 13096 16504 13124 16544
rect 13725 16541 13737 16575
rect 13771 16572 13783 16575
rect 14200 16572 14228 16612
rect 13771 16544 14228 16572
rect 14277 16575 14335 16581
rect 13771 16541 13783 16544
rect 13725 16535 13783 16541
rect 14277 16541 14289 16575
rect 14323 16572 14335 16575
rect 14476 16572 14504 16612
rect 15028 16612 15884 16640
rect 15028 16572 15056 16612
rect 14323 16544 14357 16572
rect 14476 16544 15056 16572
rect 15289 16575 15347 16581
rect 14323 16541 14335 16544
rect 14277 16535 14335 16541
rect 15289 16541 15301 16575
rect 15335 16572 15347 16575
rect 15378 16572 15384 16584
rect 15335 16544 15384 16572
rect 15335 16541 15347 16544
rect 15289 16535 15347 16541
rect 12943 16476 13124 16504
rect 12943 16473 12955 16476
rect 12897 16467 12955 16473
rect 13170 16464 13176 16516
rect 13228 16504 13234 16516
rect 13268 16507 13326 16513
rect 13268 16504 13280 16507
rect 13228 16476 13280 16504
rect 13228 16464 13234 16476
rect 13268 16473 13280 16476
rect 13314 16473 13326 16507
rect 13268 16467 13326 16473
rect 13538 16464 13544 16516
rect 13596 16504 13602 16516
rect 14292 16504 14320 16535
rect 15378 16532 15384 16544
rect 15436 16532 15442 16584
rect 15856 16581 15884 16612
rect 16022 16600 16028 16652
rect 16080 16640 16086 16652
rect 16080 16612 17172 16640
rect 16080 16600 16086 16612
rect 15841 16575 15899 16581
rect 15841 16541 15853 16575
rect 15887 16541 15899 16575
rect 16574 16572 16580 16584
rect 16514 16544 16580 16572
rect 15841 16535 15899 16541
rect 16574 16532 16580 16544
rect 16632 16572 16638 16584
rect 17144 16581 17172 16612
rect 16945 16575 17003 16581
rect 16945 16572 16957 16575
rect 16632 16544 16957 16572
rect 16632 16532 16638 16544
rect 16945 16541 16957 16544
rect 16991 16541 17003 16575
rect 16945 16535 17003 16541
rect 17129 16575 17187 16581
rect 17129 16541 17141 16575
rect 17175 16541 17187 16575
rect 17129 16535 17187 16541
rect 17405 16575 17463 16581
rect 17405 16541 17417 16575
rect 17451 16541 17463 16575
rect 17405 16535 17463 16541
rect 14369 16507 14427 16513
rect 14369 16504 14381 16507
rect 13596 16476 14381 16504
rect 13596 16464 13602 16476
rect 14369 16473 14381 16476
rect 14415 16473 14427 16507
rect 14369 16467 14427 16473
rect 14734 16464 14740 16516
rect 14792 16504 14798 16516
rect 14792 16476 15056 16504
rect 14792 16464 14798 16476
rect 12986 16436 12992 16448
rect 12452 16408 12992 16436
rect 12227 16399 12285 16405
rect 12986 16396 12992 16408
rect 13044 16396 13050 16448
rect 13078 16396 13084 16448
rect 13136 16396 13142 16448
rect 13354 16396 13360 16448
rect 13412 16396 13418 16448
rect 13446 16396 13452 16448
rect 13504 16436 13510 16448
rect 14093 16439 14151 16445
rect 14093 16436 14105 16439
rect 13504 16408 14105 16436
rect 13504 16396 13510 16408
rect 14093 16405 14105 16408
rect 14139 16405 14151 16439
rect 15028 16436 15056 16476
rect 15102 16464 15108 16516
rect 15160 16464 15166 16516
rect 15197 16507 15255 16513
rect 15197 16473 15209 16507
rect 15243 16504 15255 16507
rect 15562 16504 15568 16516
rect 15243 16476 15568 16504
rect 15243 16473 15255 16476
rect 15197 16467 15255 16473
rect 15562 16464 15568 16476
rect 15620 16464 15626 16516
rect 16666 16504 16672 16516
rect 16224 16476 16672 16504
rect 16224 16436 16252 16476
rect 16666 16464 16672 16476
rect 16724 16464 16730 16516
rect 16758 16464 16764 16516
rect 16816 16504 16822 16516
rect 16853 16507 16911 16513
rect 16853 16504 16865 16507
rect 16816 16476 16865 16504
rect 16816 16464 16822 16476
rect 16853 16473 16865 16476
rect 16899 16473 16911 16507
rect 17420 16504 17448 16535
rect 17494 16532 17500 16584
rect 17552 16572 17558 16584
rect 17681 16575 17739 16581
rect 17681 16572 17693 16575
rect 17552 16544 17693 16572
rect 17552 16532 17558 16544
rect 17681 16541 17693 16544
rect 17727 16541 17739 16575
rect 17681 16535 17739 16541
rect 17770 16532 17776 16584
rect 17828 16532 17834 16584
rect 17865 16575 17923 16581
rect 17865 16541 17877 16575
rect 17911 16572 17923 16575
rect 18049 16575 18107 16581
rect 18049 16572 18061 16575
rect 17911 16544 18061 16572
rect 17911 16541 17923 16544
rect 17865 16535 17923 16541
rect 18049 16541 18061 16544
rect 18095 16541 18107 16575
rect 18049 16535 18107 16541
rect 18322 16532 18328 16584
rect 18380 16532 18386 16584
rect 16853 16467 16911 16473
rect 16960 16476 17448 16504
rect 15028 16408 16252 16436
rect 14093 16399 14151 16405
rect 16298 16396 16304 16448
rect 16356 16436 16362 16448
rect 16960 16436 16988 16476
rect 16356 16408 16988 16436
rect 16356 16396 16362 16408
rect 17218 16396 17224 16448
rect 17276 16396 17282 16448
rect 1104 16346 18860 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 18860 16346
rect 1104 16272 18860 16294
rect 1486 16192 1492 16244
rect 1544 16232 1550 16244
rect 1857 16235 1915 16241
rect 1857 16232 1869 16235
rect 1544 16204 1869 16232
rect 1544 16192 1550 16204
rect 1857 16201 1869 16204
rect 1903 16201 1915 16235
rect 1857 16195 1915 16201
rect 5721 16235 5779 16241
rect 5721 16201 5733 16235
rect 5767 16232 5779 16235
rect 7466 16232 7472 16244
rect 5767 16204 7472 16232
rect 5767 16201 5779 16204
rect 5721 16195 5779 16201
rect 7466 16192 7472 16204
rect 7524 16192 7530 16244
rect 8754 16192 8760 16244
rect 8812 16232 8818 16244
rect 9217 16235 9275 16241
rect 9217 16232 9229 16235
rect 8812 16204 9229 16232
rect 8812 16192 8818 16204
rect 9217 16201 9229 16204
rect 9263 16201 9275 16235
rect 9217 16195 9275 16201
rect 9306 16192 9312 16244
rect 9364 16232 9370 16244
rect 9364 16204 11284 16232
rect 9364 16192 9370 16204
rect 8573 16167 8631 16173
rect 4264 16136 5396 16164
rect 1302 16056 1308 16108
rect 1360 16096 1366 16108
rect 4264 16105 4292 16136
rect 5368 16105 5396 16136
rect 8573 16133 8585 16167
rect 8619 16164 8631 16167
rect 11146 16164 11152 16176
rect 8619 16136 11152 16164
rect 8619 16133 8631 16136
rect 8573 16127 8631 16133
rect 11146 16124 11152 16136
rect 11204 16124 11210 16176
rect 11256 16164 11284 16204
rect 11698 16192 11704 16244
rect 11756 16192 11762 16244
rect 12158 16232 12164 16244
rect 11808 16204 12164 16232
rect 11808 16164 11836 16204
rect 12158 16192 12164 16204
rect 12216 16192 12222 16244
rect 12434 16192 12440 16244
rect 12492 16232 12498 16244
rect 12989 16235 13047 16241
rect 12989 16232 13001 16235
rect 12492 16204 13001 16232
rect 12492 16192 12498 16204
rect 12989 16201 13001 16204
rect 13035 16201 13047 16235
rect 12989 16195 13047 16201
rect 13262 16192 13268 16244
rect 13320 16192 13326 16244
rect 13998 16192 14004 16244
rect 14056 16192 14062 16244
rect 15102 16192 15108 16244
rect 15160 16192 15166 16244
rect 15654 16192 15660 16244
rect 15712 16241 15718 16244
rect 15712 16235 15731 16241
rect 15719 16201 15731 16235
rect 15712 16195 15731 16201
rect 15841 16235 15899 16241
rect 15841 16201 15853 16235
rect 15887 16232 15899 16235
rect 16574 16232 16580 16244
rect 15887 16204 16580 16232
rect 15887 16201 15899 16204
rect 15841 16195 15899 16201
rect 15712 16192 15718 16195
rect 16574 16192 16580 16204
rect 16632 16192 16638 16244
rect 16850 16192 16856 16244
rect 16908 16192 16914 16244
rect 17405 16235 17463 16241
rect 17405 16201 17417 16235
rect 17451 16232 17463 16235
rect 17494 16232 17500 16244
rect 17451 16204 17500 16232
rect 17451 16201 17463 16204
rect 17405 16195 17463 16201
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 17954 16192 17960 16244
rect 18012 16192 18018 16244
rect 18506 16192 18512 16244
rect 18564 16192 18570 16244
rect 11256 16136 11836 16164
rect 12069 16167 12127 16173
rect 12069 16133 12081 16167
rect 12115 16164 12127 16167
rect 12345 16167 12403 16173
rect 12345 16164 12357 16167
rect 12115 16136 12357 16164
rect 12115 16133 12127 16136
rect 12069 16127 12127 16133
rect 12345 16133 12357 16136
rect 12391 16133 12403 16167
rect 13354 16164 13360 16176
rect 12345 16127 12403 16133
rect 12544 16136 13360 16164
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 1360 16068 1409 16096
rect 1360 16056 1366 16068
rect 1397 16065 1409 16068
rect 1443 16096 1455 16099
rect 1673 16099 1731 16105
rect 1673 16096 1685 16099
rect 1443 16068 1685 16096
rect 1443 16065 1455 16068
rect 1397 16059 1455 16065
rect 1673 16065 1685 16068
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 4249 16099 4307 16105
rect 4249 16065 4261 16099
rect 4295 16065 4307 16099
rect 5169 16099 5227 16105
rect 5169 16096 5181 16099
rect 4249 16059 4307 16065
rect 4356 16068 5181 16096
rect 4157 16031 4215 16037
rect 4157 15997 4169 16031
rect 4203 16028 4215 16031
rect 4356 16028 4384 16068
rect 5169 16065 5181 16068
rect 5215 16065 5227 16099
rect 5169 16059 5227 16065
rect 5353 16099 5411 16105
rect 5353 16065 5365 16099
rect 5399 16065 5411 16099
rect 5353 16059 5411 16065
rect 4203 16000 4384 16028
rect 4203 15997 4215 16000
rect 4157 15991 4215 15997
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15960 1639 15963
rect 4172 15960 4200 15991
rect 4982 15988 4988 16040
rect 5040 15988 5046 16040
rect 5368 16028 5396 16059
rect 5626 16056 5632 16108
rect 5684 16056 5690 16108
rect 5810 16056 5816 16108
rect 5868 16056 5874 16108
rect 6914 16056 6920 16108
rect 6972 16056 6978 16108
rect 9125 16099 9183 16105
rect 9125 16065 9137 16099
rect 9171 16096 9183 16099
rect 9171 16068 9720 16096
rect 9171 16065 9183 16068
rect 9125 16059 9183 16065
rect 5828 16028 5856 16056
rect 5368 16000 5856 16028
rect 7006 15988 7012 16040
rect 7064 15988 7070 16040
rect 9214 15988 9220 16040
rect 9272 16028 9278 16040
rect 9309 16031 9367 16037
rect 9309 16028 9321 16031
rect 9272 16000 9321 16028
rect 9272 15988 9278 16000
rect 9309 15997 9321 16000
rect 9355 15997 9367 16031
rect 9692 16028 9720 16068
rect 9766 16056 9772 16108
rect 9824 16096 9830 16108
rect 10229 16099 10287 16105
rect 10229 16096 10241 16099
rect 9824 16068 10241 16096
rect 9824 16056 9830 16068
rect 10229 16065 10241 16068
rect 10275 16065 10287 16099
rect 10229 16059 10287 16065
rect 10873 16099 10931 16105
rect 10873 16065 10885 16099
rect 10919 16065 10931 16099
rect 10873 16059 10931 16065
rect 10965 16099 11023 16105
rect 10965 16065 10977 16099
rect 11011 16096 11023 16099
rect 11238 16096 11244 16108
rect 11011 16068 11244 16096
rect 11011 16065 11023 16068
rect 10965 16059 11023 16065
rect 10045 16031 10103 16037
rect 10045 16028 10057 16031
rect 9692 16000 10057 16028
rect 9309 15991 9367 15997
rect 10045 15997 10057 16000
rect 10091 16028 10103 16031
rect 10594 16028 10600 16040
rect 10091 16000 10600 16028
rect 10091 15997 10103 16000
rect 10045 15991 10103 15997
rect 10594 15988 10600 16000
rect 10652 15988 10658 16040
rect 10888 16028 10916 16059
rect 11238 16056 11244 16068
rect 11296 16056 11302 16108
rect 11882 16056 11888 16108
rect 11940 16056 11946 16108
rect 11974 16056 11980 16108
rect 12032 16056 12038 16108
rect 12233 16099 12291 16105
rect 12233 16065 12245 16099
rect 12279 16065 12291 16099
rect 12233 16059 12291 16065
rect 10888 16000 11008 16028
rect 1627 15932 4200 15960
rect 7285 15963 7343 15969
rect 1627 15929 1639 15932
rect 1581 15923 1639 15929
rect 7285 15929 7297 15963
rect 7331 15960 7343 15963
rect 8202 15960 8208 15972
rect 7331 15932 8208 15960
rect 7331 15929 7343 15932
rect 7285 15923 7343 15929
rect 8202 15920 8208 15932
rect 8260 15920 8266 15972
rect 9858 15920 9864 15972
rect 9916 15960 9922 15972
rect 10505 15963 10563 15969
rect 10505 15960 10517 15963
rect 9916 15932 10517 15960
rect 9916 15920 9922 15932
rect 10505 15929 10517 15932
rect 10551 15929 10563 15963
rect 10505 15923 10563 15929
rect 5261 15895 5319 15901
rect 5261 15861 5273 15895
rect 5307 15892 5319 15895
rect 5626 15892 5632 15904
rect 5307 15864 5632 15892
rect 5307 15861 5319 15864
rect 5261 15855 5319 15861
rect 5626 15852 5632 15864
rect 5684 15852 5690 15904
rect 8478 15852 8484 15904
rect 8536 15852 8542 15904
rect 8754 15852 8760 15904
rect 8812 15852 8818 15904
rect 10410 15852 10416 15904
rect 10468 15852 10474 15904
rect 10778 15852 10784 15904
rect 10836 15892 10842 15904
rect 10980 15892 11008 16000
rect 11054 15988 11060 16040
rect 11112 15988 11118 16040
rect 11238 15920 11244 15972
rect 11296 15960 11302 15972
rect 12242 15960 12270 16059
rect 12434 16056 12440 16108
rect 12492 16096 12498 16108
rect 12544 16105 12572 16136
rect 13354 16124 13360 16136
rect 13412 16124 13418 16176
rect 15473 16167 15531 16173
rect 15473 16164 15485 16167
rect 13464 16136 15485 16164
rect 12529 16099 12587 16105
rect 12529 16096 12541 16099
rect 12492 16068 12541 16096
rect 12492 16056 12498 16068
rect 12529 16065 12541 16068
rect 12575 16065 12587 16099
rect 12529 16059 12587 16065
rect 12618 16056 12624 16108
rect 12676 16056 12682 16108
rect 12710 16056 12716 16108
rect 12768 16096 12774 16108
rect 12897 16099 12955 16105
rect 12897 16096 12909 16099
rect 12768 16068 12909 16096
rect 12768 16056 12774 16068
rect 12897 16065 12909 16068
rect 12943 16065 12955 16099
rect 12897 16059 12955 16065
rect 13170 16056 13176 16108
rect 13228 16096 13234 16108
rect 13464 16096 13492 16136
rect 15473 16133 15485 16136
rect 15519 16164 15531 16167
rect 16022 16164 16028 16176
rect 15519 16136 16028 16164
rect 15519 16133 15531 16136
rect 15473 16127 15531 16133
rect 16022 16124 16028 16136
rect 16080 16124 16086 16176
rect 16298 16124 16304 16176
rect 16356 16164 16362 16176
rect 17037 16167 17095 16173
rect 17037 16164 17049 16167
rect 16356 16136 17049 16164
rect 16356 16124 16362 16136
rect 17037 16133 17049 16136
rect 17083 16133 17095 16167
rect 17037 16127 17095 16133
rect 13228 16068 13492 16096
rect 13817 16099 13875 16105
rect 13228 16056 13234 16068
rect 13817 16065 13829 16099
rect 13863 16096 13875 16099
rect 13906 16096 13912 16108
rect 13863 16068 13912 16096
rect 13863 16065 13875 16068
rect 13817 16059 13875 16065
rect 13906 16056 13912 16068
rect 13964 16096 13970 16108
rect 14550 16096 14556 16108
rect 13964 16068 14556 16096
rect 13964 16056 13970 16068
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 15289 16099 15347 16105
rect 15289 16065 15301 16099
rect 15335 16065 15347 16099
rect 15289 16059 15347 16065
rect 15304 16028 15332 16059
rect 16482 16056 16488 16108
rect 16540 16096 16546 16108
rect 17497 16099 17555 16105
rect 17497 16096 17509 16099
rect 16540 16068 17509 16096
rect 16540 16056 16546 16068
rect 17497 16065 17509 16068
rect 17543 16065 17555 16099
rect 17972 16096 18000 16192
rect 18233 16099 18291 16105
rect 18233 16096 18245 16099
rect 17972 16068 18245 16096
rect 17497 16059 17555 16065
rect 18233 16065 18245 16068
rect 18279 16065 18291 16099
rect 18233 16059 18291 16065
rect 15930 16028 15936 16040
rect 15304 16000 15936 16028
rect 15930 15988 15936 16000
rect 15988 16028 15994 16040
rect 17218 16028 17224 16040
rect 15988 16000 17224 16028
rect 15988 15988 15994 16000
rect 17218 15988 17224 16000
rect 17276 15988 17282 16040
rect 11296 15932 12270 15960
rect 12406 15932 12848 15960
rect 11296 15920 11302 15932
rect 12406 15892 12434 15932
rect 12820 15904 12848 15932
rect 13078 15920 13084 15972
rect 13136 15960 13142 15972
rect 15746 15960 15752 15972
rect 13136 15932 15752 15960
rect 13136 15920 13142 15932
rect 10836 15864 12434 15892
rect 10836 15852 10842 15864
rect 12802 15852 12808 15904
rect 12860 15852 12866 15904
rect 13722 15852 13728 15904
rect 13780 15852 13786 15904
rect 15672 15901 15700 15932
rect 15746 15920 15752 15932
rect 15804 15960 15810 15972
rect 16574 15960 16580 15972
rect 15804 15932 16580 15960
rect 15804 15920 15810 15932
rect 16574 15920 16580 15932
rect 16632 15920 16638 15972
rect 15657 15895 15715 15901
rect 15657 15861 15669 15895
rect 15703 15861 15715 15895
rect 15657 15855 15715 15861
rect 16022 15852 16028 15904
rect 16080 15892 16086 15904
rect 18049 15895 18107 15901
rect 18049 15892 18061 15895
rect 16080 15864 18061 15892
rect 16080 15852 16086 15864
rect 18049 15861 18061 15864
rect 18095 15861 18107 15895
rect 18049 15855 18107 15861
rect 1104 15802 18860 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 18860 15802
rect 1104 15728 18860 15750
rect 7009 15691 7067 15697
rect 7009 15657 7021 15691
rect 7055 15688 7067 15691
rect 7055 15660 11192 15688
rect 7055 15657 7067 15660
rect 7009 15651 7067 15657
rect 8205 15623 8263 15629
rect 8205 15589 8217 15623
rect 8251 15620 8263 15623
rect 9306 15620 9312 15632
rect 8251 15592 9312 15620
rect 8251 15589 8263 15592
rect 8205 15583 8263 15589
rect 9306 15580 9312 15592
rect 9364 15580 9370 15632
rect 9766 15620 9772 15632
rect 9600 15592 9772 15620
rect 4982 15512 4988 15564
rect 5040 15512 5046 15564
rect 6730 15512 6736 15564
rect 6788 15512 6794 15564
rect 9600 15561 9628 15592
rect 9766 15580 9772 15592
rect 9824 15580 9830 15632
rect 9585 15555 9643 15561
rect 9585 15521 9597 15555
rect 9631 15521 9643 15555
rect 9585 15515 9643 15521
rect 10045 15555 10103 15561
rect 10045 15521 10057 15555
rect 10091 15552 10103 15555
rect 11164 15552 11192 15660
rect 11238 15648 11244 15700
rect 11296 15648 11302 15700
rect 12986 15648 12992 15700
rect 13044 15688 13050 15700
rect 13633 15691 13691 15697
rect 13633 15688 13645 15691
rect 13044 15660 13645 15688
rect 13044 15648 13050 15660
rect 13633 15657 13645 15660
rect 13679 15688 13691 15691
rect 13722 15688 13728 15700
rect 13679 15660 13728 15688
rect 13679 15657 13691 15660
rect 13633 15651 13691 15657
rect 13722 15648 13728 15660
rect 13780 15648 13786 15700
rect 11882 15580 11888 15632
rect 11940 15620 11946 15632
rect 12069 15623 12127 15629
rect 12069 15620 12081 15623
rect 11940 15592 12081 15620
rect 11940 15580 11946 15592
rect 12069 15589 12081 15592
rect 12115 15589 12127 15623
rect 12069 15583 12127 15589
rect 13357 15623 13415 15629
rect 13357 15589 13369 15623
rect 13403 15620 13415 15623
rect 13446 15620 13452 15632
rect 13403 15592 13452 15620
rect 13403 15589 13415 15592
rect 13357 15583 13415 15589
rect 11974 15552 11980 15564
rect 10091 15524 10916 15552
rect 11164 15524 11980 15552
rect 10091 15521 10103 15524
rect 10045 15515 10103 15521
rect 5258 15444 5264 15496
rect 5316 15444 5322 15496
rect 5626 15444 5632 15496
rect 5684 15444 5690 15496
rect 6546 15444 6552 15496
rect 6604 15484 6610 15496
rect 6641 15487 6699 15493
rect 6641 15484 6653 15487
rect 6604 15456 6653 15484
rect 6604 15444 6610 15456
rect 6641 15453 6653 15456
rect 6687 15453 6699 15487
rect 6641 15447 6699 15453
rect 9401 15487 9459 15493
rect 9401 15453 9413 15487
rect 9447 15453 9459 15487
rect 9401 15447 9459 15453
rect 5905 15419 5963 15425
rect 5905 15385 5917 15419
rect 5951 15416 5963 15419
rect 6454 15416 6460 15428
rect 5951 15388 6460 15416
rect 5951 15385 5963 15388
rect 5905 15379 5963 15385
rect 6454 15376 6460 15388
rect 6512 15416 6518 15428
rect 8389 15419 8447 15425
rect 8389 15416 8401 15419
rect 6512 15388 8401 15416
rect 6512 15376 6518 15388
rect 8389 15385 8401 15388
rect 8435 15385 8447 15419
rect 8389 15379 8447 15385
rect 8757 15419 8815 15425
rect 8757 15385 8769 15419
rect 8803 15416 8815 15419
rect 8846 15416 8852 15428
rect 8803 15388 8852 15416
rect 8803 15385 8815 15388
rect 8757 15379 8815 15385
rect 8846 15376 8852 15388
rect 8904 15376 8910 15428
rect 9416 15416 9444 15447
rect 9674 15444 9680 15496
rect 9732 15444 9738 15496
rect 9766 15444 9772 15496
rect 9824 15444 9830 15496
rect 9861 15487 9919 15493
rect 9861 15453 9873 15487
rect 9907 15484 9919 15487
rect 9950 15484 9956 15496
rect 9907 15456 9956 15484
rect 9907 15453 9919 15456
rect 9861 15447 9919 15453
rect 9950 15444 9956 15456
rect 10008 15444 10014 15496
rect 10410 15444 10416 15496
rect 10468 15484 10474 15496
rect 10778 15493 10784 15496
rect 10597 15487 10655 15493
rect 10597 15484 10609 15487
rect 10468 15456 10609 15484
rect 10468 15444 10474 15456
rect 10597 15453 10609 15456
rect 10643 15453 10655 15487
rect 10597 15447 10655 15453
rect 10745 15487 10784 15493
rect 10745 15453 10757 15487
rect 10745 15447 10784 15453
rect 10778 15444 10784 15447
rect 10836 15444 10842 15496
rect 10888 15484 10916 15524
rect 11974 15512 11980 15524
rect 12032 15512 12038 15564
rect 12084 15552 12112 15583
rect 13446 15580 13452 15592
rect 13504 15580 13510 15632
rect 13814 15580 13820 15632
rect 13872 15620 13878 15632
rect 13872 15592 14412 15620
rect 13872 15580 13878 15592
rect 12618 15552 12624 15564
rect 12084 15524 12624 15552
rect 12618 15512 12624 15524
rect 12676 15552 12682 15564
rect 14384 15561 14412 15592
rect 14093 15555 14151 15561
rect 14093 15552 14105 15555
rect 12676 15524 14105 15552
rect 12676 15512 12682 15524
rect 14093 15521 14105 15524
rect 14139 15521 14151 15555
rect 14093 15515 14151 15521
rect 14369 15555 14427 15561
rect 14369 15521 14381 15555
rect 14415 15521 14427 15555
rect 14369 15515 14427 15521
rect 15194 15512 15200 15564
rect 15252 15552 15258 15564
rect 15654 15552 15660 15564
rect 15252 15524 15660 15552
rect 15252 15512 15258 15524
rect 15654 15512 15660 15524
rect 15712 15552 15718 15564
rect 15933 15555 15991 15561
rect 15712 15524 15792 15552
rect 15712 15512 15718 15524
rect 11062 15487 11120 15493
rect 11062 15484 11074 15487
rect 10888 15456 11074 15484
rect 11062 15453 11074 15456
rect 11108 15453 11120 15487
rect 11062 15447 11120 15453
rect 12345 15487 12403 15493
rect 12345 15453 12357 15487
rect 12391 15484 12403 15487
rect 12434 15484 12440 15496
rect 12391 15456 12440 15484
rect 12391 15453 12403 15456
rect 12345 15447 12403 15453
rect 12434 15444 12440 15456
rect 12492 15444 12498 15496
rect 13078 15444 13084 15496
rect 13136 15484 13142 15496
rect 13136 15456 13584 15484
rect 13136 15444 13142 15456
rect 10502 15416 10508 15428
rect 9416 15388 10508 15416
rect 10502 15376 10508 15388
rect 10560 15376 10566 15428
rect 10873 15419 10931 15425
rect 10873 15385 10885 15419
rect 10919 15385 10931 15419
rect 10873 15379 10931 15385
rect 8478 15308 8484 15360
rect 8536 15308 8542 15360
rect 8570 15308 8576 15360
rect 8628 15308 8634 15360
rect 8662 15308 8668 15360
rect 8720 15348 8726 15360
rect 10778 15348 10784 15360
rect 8720 15320 10784 15348
rect 8720 15308 8726 15320
rect 10778 15308 10784 15320
rect 10836 15308 10842 15360
rect 10888 15348 10916 15379
rect 10962 15376 10968 15428
rect 11020 15376 11026 15428
rect 12526 15416 12532 15428
rect 11348 15388 12532 15416
rect 11348 15348 11376 15388
rect 12526 15376 12532 15388
rect 12584 15376 12590 15428
rect 13354 15376 13360 15428
rect 13412 15416 13418 15428
rect 13449 15419 13507 15425
rect 13449 15416 13461 15419
rect 13412 15388 13461 15416
rect 13412 15376 13418 15388
rect 13449 15385 13461 15388
rect 13495 15385 13507 15419
rect 13556 15416 13584 15456
rect 14458 15444 14464 15496
rect 14516 15444 14522 15496
rect 15378 15444 15384 15496
rect 15436 15444 15442 15496
rect 15562 15444 15568 15496
rect 15620 15444 15626 15496
rect 15764 15493 15792 15524
rect 15933 15521 15945 15555
rect 15979 15552 15991 15555
rect 16022 15552 16028 15564
rect 15979 15524 16028 15552
rect 15979 15521 15991 15524
rect 15933 15515 15991 15521
rect 16022 15512 16028 15524
rect 16080 15552 16086 15564
rect 16669 15555 16727 15561
rect 16669 15552 16681 15555
rect 16080 15524 16681 15552
rect 16080 15512 16086 15524
rect 16669 15521 16681 15524
rect 16715 15521 16727 15555
rect 16669 15515 16727 15521
rect 15749 15487 15807 15493
rect 15749 15453 15761 15487
rect 15795 15453 15807 15487
rect 15749 15447 15807 15453
rect 16114 15444 16120 15496
rect 16172 15444 16178 15496
rect 16574 15444 16580 15496
rect 16632 15484 16638 15496
rect 16761 15487 16819 15493
rect 16761 15484 16773 15487
rect 16632 15456 16773 15484
rect 16632 15444 16638 15456
rect 16761 15453 16773 15456
rect 16807 15453 16819 15487
rect 16761 15447 16819 15453
rect 13649 15419 13707 15425
rect 13649 15416 13661 15419
rect 13556 15388 13661 15416
rect 13449 15379 13507 15385
rect 13649 15385 13661 15388
rect 13695 15385 13707 15419
rect 13649 15379 13707 15385
rect 10888 15320 11376 15348
rect 11422 15308 11428 15360
rect 11480 15348 11486 15360
rect 11885 15351 11943 15357
rect 11885 15348 11897 15351
rect 11480 15320 11897 15348
rect 11480 15308 11486 15320
rect 11885 15317 11897 15320
rect 11931 15317 11943 15351
rect 11885 15311 11943 15317
rect 12986 15308 12992 15360
rect 13044 15348 13050 15360
rect 13173 15351 13231 15357
rect 13173 15348 13185 15351
rect 13044 15320 13185 15348
rect 13044 15308 13050 15320
rect 13173 15317 13185 15320
rect 13219 15317 13231 15351
rect 13173 15311 13231 15317
rect 17126 15308 17132 15360
rect 17184 15308 17190 15360
rect 1104 15258 18860 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 18860 15258
rect 1104 15184 18860 15206
rect 1581 15147 1639 15153
rect 1581 15113 1593 15147
rect 1627 15144 1639 15147
rect 1627 15116 2774 15144
rect 1627 15113 1639 15116
rect 1581 15107 1639 15113
rect 1302 14968 1308 15020
rect 1360 15008 1366 15020
rect 1397 15011 1455 15017
rect 1397 15008 1409 15011
rect 1360 14980 1409 15008
rect 1360 14968 1366 14980
rect 1397 14977 1409 14980
rect 1443 15008 1455 15011
rect 1673 15011 1731 15017
rect 1673 15008 1685 15011
rect 1443 14980 1685 15008
rect 1443 14977 1455 14980
rect 1397 14971 1455 14977
rect 1673 14977 1685 14980
rect 1719 14977 1731 15011
rect 2746 15008 2774 15116
rect 6730 15104 6736 15156
rect 6788 15104 6794 15156
rect 8757 15147 8815 15153
rect 8757 15113 8769 15147
rect 8803 15144 8815 15147
rect 9766 15144 9772 15156
rect 8803 15116 9772 15144
rect 8803 15113 8815 15116
rect 8757 15107 8815 15113
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 12802 15104 12808 15156
rect 12860 15144 12866 15156
rect 13541 15147 13599 15153
rect 13541 15144 13553 15147
rect 12860 15116 13553 15144
rect 12860 15104 12866 15116
rect 13541 15113 13553 15116
rect 13587 15113 13599 15147
rect 13541 15107 13599 15113
rect 5534 15076 5540 15088
rect 4632 15048 5540 15076
rect 4062 15008 4068 15020
rect 2746 14980 4068 15008
rect 1673 14971 1731 14977
rect 4062 14968 4068 14980
rect 4120 15008 4126 15020
rect 4632 15017 4660 15048
rect 5534 15036 5540 15048
rect 5592 15076 5598 15088
rect 6748 15076 6776 15104
rect 8846 15076 8852 15088
rect 5592 15048 6776 15076
rect 8772 15048 8852 15076
rect 5592 15036 5598 15048
rect 4433 15011 4491 15017
rect 4433 15008 4445 15011
rect 4120 14980 4445 15008
rect 4120 14968 4126 14980
rect 4433 14977 4445 14980
rect 4479 14977 4491 15011
rect 4433 14971 4491 14977
rect 4617 15011 4675 15017
rect 4617 14977 4629 15011
rect 4663 14977 4675 15011
rect 4617 14971 4675 14977
rect 4798 14968 4804 15020
rect 4856 15008 4862 15020
rect 4985 15011 5043 15017
rect 4985 15008 4997 15011
rect 4856 14980 4997 15008
rect 4856 14968 4862 14980
rect 4985 14977 4997 14980
rect 5031 14977 5043 15011
rect 4985 14971 5043 14977
rect 6730 14968 6736 15020
rect 6788 15008 6794 15020
rect 8113 15011 8171 15017
rect 8113 15008 8125 15011
rect 6788 14980 8125 15008
rect 6788 14968 6794 14980
rect 8113 14977 8125 14980
rect 8159 15008 8171 15011
rect 8478 15008 8484 15020
rect 8159 14980 8484 15008
rect 8159 14977 8171 14980
rect 8113 14971 8171 14977
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 8772 15017 8800 15048
rect 8846 15036 8852 15048
rect 8904 15076 8910 15088
rect 15286 15076 15292 15088
rect 8904 15048 15292 15076
rect 8904 15036 8910 15048
rect 15286 15036 15292 15048
rect 15344 15076 15350 15088
rect 16114 15076 16120 15088
rect 15344 15048 16120 15076
rect 15344 15036 15350 15048
rect 8757 15011 8815 15017
rect 8757 14977 8769 15011
rect 8803 14977 8815 15011
rect 8757 14971 8815 14977
rect 9033 15011 9091 15017
rect 9033 14977 9045 15011
rect 9079 15008 9091 15011
rect 9306 15008 9312 15020
rect 9079 14980 9312 15008
rect 9079 14977 9091 14980
rect 9033 14971 9091 14977
rect 9306 14968 9312 14980
rect 9364 14968 9370 15020
rect 12621 15011 12679 15017
rect 12621 14977 12633 15011
rect 12667 15008 12679 15011
rect 12894 15008 12900 15020
rect 12667 14980 12900 15008
rect 12667 14977 12679 14980
rect 12621 14971 12679 14977
rect 12894 14968 12900 14980
rect 12952 14968 12958 15020
rect 13446 14968 13452 15020
rect 13504 14968 13510 15020
rect 13633 15011 13691 15017
rect 13633 14977 13645 15011
rect 13679 15008 13691 15011
rect 13814 15008 13820 15020
rect 13679 14980 13820 15008
rect 13679 14977 13691 14980
rect 13633 14971 13691 14977
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 15378 14968 15384 15020
rect 15436 15008 15442 15020
rect 15473 15011 15531 15017
rect 15473 15008 15485 15011
rect 15436 14980 15485 15008
rect 15436 14968 15442 14980
rect 15473 14977 15485 14980
rect 15519 14977 15531 15011
rect 15473 14971 15531 14977
rect 15654 14968 15660 15020
rect 15712 14968 15718 15020
rect 15764 15017 15792 15048
rect 16114 15036 16120 15048
rect 16172 15036 16178 15088
rect 15749 15011 15807 15017
rect 15749 14977 15761 15011
rect 15795 14977 15807 15011
rect 15749 14971 15807 14977
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14940 4583 14943
rect 5077 14943 5135 14949
rect 5077 14940 5089 14943
rect 4571 14912 5089 14940
rect 4571 14909 4583 14912
rect 4525 14903 4583 14909
rect 5077 14909 5089 14912
rect 5123 14940 5135 14943
rect 5258 14940 5264 14952
rect 5123 14912 5264 14940
rect 5123 14909 5135 14912
rect 5077 14903 5135 14909
rect 5258 14900 5264 14912
rect 5316 14900 5322 14952
rect 6454 14900 6460 14952
rect 6512 14940 6518 14952
rect 7929 14943 7987 14949
rect 7929 14940 7941 14943
rect 6512 14912 7941 14940
rect 6512 14900 6518 14912
rect 7929 14909 7941 14912
rect 7975 14909 7987 14943
rect 7929 14903 7987 14909
rect 8297 14943 8355 14949
rect 8297 14909 8309 14943
rect 8343 14940 8355 14943
rect 8570 14940 8576 14952
rect 8343 14912 8576 14940
rect 8343 14909 8355 14912
rect 8297 14903 8355 14909
rect 5353 14875 5411 14881
rect 5353 14841 5365 14875
rect 5399 14872 5411 14875
rect 5442 14872 5448 14884
rect 5399 14844 5448 14872
rect 5399 14841 5411 14844
rect 5353 14835 5411 14841
rect 5442 14832 5448 14844
rect 5500 14832 5506 14884
rect 7944 14872 7972 14903
rect 8570 14900 8576 14912
rect 8628 14940 8634 14952
rect 8849 14943 8907 14949
rect 8628 14912 8800 14940
rect 8628 14900 8634 14912
rect 8772 14884 8800 14912
rect 8849 14909 8861 14943
rect 8895 14940 8907 14943
rect 9950 14940 9956 14952
rect 8895 14912 9956 14940
rect 8895 14909 8907 14912
rect 8849 14903 8907 14909
rect 9950 14900 9956 14912
rect 10008 14900 10014 14952
rect 15562 14900 15568 14952
rect 15620 14900 15626 14952
rect 8386 14872 8392 14884
rect 7944 14844 8392 14872
rect 8386 14832 8392 14844
rect 8444 14832 8450 14884
rect 8754 14832 8760 14884
rect 8812 14832 8818 14884
rect 12342 14764 12348 14816
rect 12400 14804 12406 14816
rect 12437 14807 12495 14813
rect 12437 14804 12449 14807
rect 12400 14776 12449 14804
rect 12400 14764 12406 14776
rect 12437 14773 12449 14776
rect 12483 14773 12495 14807
rect 12437 14767 12495 14773
rect 15286 14764 15292 14816
rect 15344 14764 15350 14816
rect 1104 14714 18860 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 18860 14714
rect 1104 14640 18860 14662
rect 9950 14600 9956 14612
rect 8588 14572 9956 14600
rect 4062 14424 4068 14476
rect 4120 14464 4126 14476
rect 4249 14467 4307 14473
rect 4249 14464 4261 14467
rect 4120 14436 4261 14464
rect 4120 14424 4126 14436
rect 4249 14433 4261 14436
rect 4295 14433 4307 14467
rect 4249 14427 4307 14433
rect 4522 14424 4528 14476
rect 4580 14424 4586 14476
rect 6454 14424 6460 14476
rect 6512 14424 6518 14476
rect 4157 14399 4215 14405
rect 4157 14365 4169 14399
rect 4203 14396 4215 14399
rect 5534 14396 5540 14408
rect 4203 14368 5540 14396
rect 4203 14365 4215 14368
rect 4157 14359 4215 14365
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 6549 14399 6607 14405
rect 6549 14365 6561 14399
rect 6595 14396 6607 14399
rect 6730 14396 6736 14408
rect 6595 14368 6736 14396
rect 6595 14365 6607 14368
rect 6549 14359 6607 14365
rect 6730 14356 6736 14368
rect 6788 14356 6794 14408
rect 8588 14405 8616 14572
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 12713 14603 12771 14609
rect 12713 14569 12725 14603
rect 12759 14600 12771 14603
rect 13078 14600 13084 14612
rect 12759 14572 13084 14600
rect 12759 14569 12771 14572
rect 12713 14563 12771 14569
rect 13078 14560 13084 14572
rect 13136 14560 13142 14612
rect 9766 14532 9772 14544
rect 8772 14504 9772 14532
rect 8772 14405 8800 14504
rect 9766 14492 9772 14504
rect 9824 14492 9830 14544
rect 10594 14492 10600 14544
rect 10652 14492 10658 14544
rect 11514 14492 11520 14544
rect 11572 14532 11578 14544
rect 12161 14535 12219 14541
rect 12161 14532 12173 14535
rect 11572 14504 12173 14532
rect 11572 14492 11578 14504
rect 12161 14501 12173 14504
rect 12207 14532 12219 14535
rect 12618 14532 12624 14544
rect 12207 14504 12624 14532
rect 12207 14501 12219 14504
rect 12161 14495 12219 14501
rect 12618 14492 12624 14504
rect 12676 14492 12682 14544
rect 9214 14424 9220 14476
rect 9272 14464 9278 14476
rect 9493 14467 9551 14473
rect 9493 14464 9505 14467
rect 9272 14436 9505 14464
rect 9272 14424 9278 14436
rect 9493 14433 9505 14436
rect 9539 14433 9551 14467
rect 9784 14464 9812 14492
rect 10873 14467 10931 14473
rect 10873 14464 10885 14467
rect 9784 14436 10180 14464
rect 9493 14427 9551 14433
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14365 8631 14399
rect 8573 14359 8631 14365
rect 8757 14399 8815 14405
rect 8757 14365 8769 14399
rect 8803 14365 8815 14399
rect 8757 14359 8815 14365
rect 9309 14399 9367 14405
rect 9309 14365 9321 14399
rect 9355 14396 9367 14399
rect 9674 14396 9680 14408
rect 9355 14368 9680 14396
rect 9355 14365 9367 14368
rect 9309 14359 9367 14365
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 9950 14356 9956 14408
rect 10008 14396 10014 14408
rect 10152 14405 10180 14436
rect 10244 14436 10885 14464
rect 10244 14405 10272 14436
rect 10873 14433 10885 14436
rect 10919 14464 10931 14467
rect 11606 14464 11612 14476
rect 10919 14436 11612 14464
rect 10919 14433 10931 14436
rect 10873 14427 10931 14433
rect 11606 14424 11612 14436
rect 11664 14424 11670 14476
rect 12805 14467 12863 14473
rect 12805 14464 12817 14467
rect 11716 14436 12817 14464
rect 10045 14399 10103 14405
rect 10045 14396 10057 14399
rect 10008 14368 10057 14396
rect 10008 14356 10014 14368
rect 10045 14365 10057 14368
rect 10091 14365 10103 14399
rect 10045 14359 10103 14365
rect 10137 14399 10195 14405
rect 10137 14365 10149 14399
rect 10183 14365 10195 14399
rect 10137 14359 10195 14365
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 10410 14356 10416 14408
rect 10468 14356 10474 14408
rect 10965 14399 11023 14405
rect 10965 14365 10977 14399
rect 11011 14365 11023 14399
rect 10965 14359 11023 14365
rect 8665 14331 8723 14337
rect 8665 14297 8677 14331
rect 8711 14328 8723 14331
rect 9401 14331 9459 14337
rect 9401 14328 9413 14331
rect 8711 14300 9413 14328
rect 8711 14297 8723 14300
rect 8665 14291 8723 14297
rect 9401 14297 9413 14300
rect 9447 14297 9459 14331
rect 10980 14328 11008 14359
rect 11330 14356 11336 14408
rect 11388 14396 11394 14408
rect 11425 14399 11483 14405
rect 11425 14396 11437 14399
rect 11388 14368 11437 14396
rect 11388 14356 11394 14368
rect 11425 14365 11437 14368
rect 11471 14396 11483 14399
rect 11716 14396 11744 14436
rect 12805 14433 12817 14436
rect 12851 14433 12863 14467
rect 12805 14427 12863 14433
rect 14553 14467 14611 14473
rect 14553 14433 14565 14467
rect 14599 14464 14611 14467
rect 17494 14464 17500 14476
rect 14599 14436 17500 14464
rect 14599 14433 14611 14436
rect 14553 14427 14611 14433
rect 17494 14424 17500 14436
rect 17552 14424 17558 14476
rect 12618 14396 12624 14408
rect 11471 14368 11744 14396
rect 11808 14368 12624 14396
rect 11471 14365 11483 14368
rect 11425 14359 11483 14365
rect 11808 14328 11836 14368
rect 12618 14356 12624 14368
rect 12676 14396 12682 14408
rect 12986 14396 12992 14408
rect 12676 14368 12992 14396
rect 12676 14356 12682 14368
rect 12986 14356 12992 14368
rect 13044 14356 13050 14408
rect 13081 14399 13139 14405
rect 13081 14365 13093 14399
rect 13127 14396 13139 14399
rect 13630 14396 13636 14408
rect 13127 14368 13636 14396
rect 13127 14365 13139 14368
rect 13081 14359 13139 14365
rect 13630 14356 13636 14368
rect 13688 14356 13694 14408
rect 16390 14356 16396 14408
rect 16448 14356 16454 14408
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14365 16635 14399
rect 16577 14359 16635 14365
rect 12437 14331 12495 14337
rect 12437 14328 12449 14331
rect 10980 14300 11836 14328
rect 12268 14300 12449 14328
rect 9401 14291 9459 14297
rect 6914 14220 6920 14272
rect 6972 14220 6978 14272
rect 8938 14220 8944 14272
rect 8996 14220 9002 14272
rect 9490 14220 9496 14272
rect 9548 14260 9554 14272
rect 9769 14263 9827 14269
rect 9769 14260 9781 14263
rect 9548 14232 9781 14260
rect 9548 14220 9554 14232
rect 9769 14229 9781 14232
rect 9815 14229 9827 14263
rect 9769 14223 9827 14229
rect 11054 14220 11060 14272
rect 11112 14260 11118 14272
rect 11241 14263 11299 14269
rect 11241 14260 11253 14263
rect 11112 14232 11253 14260
rect 11112 14220 11118 14232
rect 11241 14229 11253 14232
rect 11287 14260 11299 14263
rect 12268 14260 12296 14300
rect 12437 14297 12449 14300
rect 12483 14297 12495 14331
rect 12437 14291 12495 14297
rect 14182 14288 14188 14340
rect 14240 14288 14246 14340
rect 14366 14288 14372 14340
rect 14424 14288 14430 14340
rect 16206 14288 16212 14340
rect 16264 14328 16270 14340
rect 16592 14328 16620 14359
rect 16264 14300 16620 14328
rect 16264 14288 16270 14300
rect 11287 14232 12296 14260
rect 11287 14229 11299 14232
rect 11241 14223 11299 14229
rect 12342 14220 12348 14272
rect 12400 14220 12406 14272
rect 12526 14220 12532 14272
rect 12584 14220 12590 14272
rect 16485 14263 16543 14269
rect 16485 14229 16497 14263
rect 16531 14260 16543 14263
rect 16942 14260 16948 14272
rect 16531 14232 16948 14260
rect 16531 14229 16543 14232
rect 16485 14223 16543 14229
rect 16942 14220 16948 14232
rect 17000 14220 17006 14272
rect 1104 14170 18860 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 18860 14170
rect 1104 14096 18860 14118
rect 4985 14059 5043 14065
rect 4985 14025 4997 14059
rect 5031 14056 5043 14059
rect 5718 14056 5724 14068
rect 5031 14028 5724 14056
rect 5031 14025 5043 14028
rect 4985 14019 5043 14025
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 7193 14059 7251 14065
rect 7193 14025 7205 14059
rect 7239 14056 7251 14059
rect 9585 14059 9643 14065
rect 7239 14028 8616 14056
rect 7239 14025 7251 14028
rect 7193 14019 7251 14025
rect 4522 13948 4528 14000
rect 4580 13988 4586 14000
rect 5353 13991 5411 13997
rect 5353 13988 5365 13991
rect 4580 13960 5365 13988
rect 4580 13948 4586 13960
rect 5353 13957 5365 13960
rect 5399 13957 5411 13991
rect 5353 13951 5411 13957
rect 6914 13948 6920 14000
rect 6972 13988 6978 14000
rect 7469 13991 7527 13997
rect 7469 13988 7481 13991
rect 6972 13960 7481 13988
rect 6972 13948 6978 13960
rect 7469 13957 7481 13960
rect 7515 13957 7527 13991
rect 7469 13951 7527 13957
rect 8294 13948 8300 14000
rect 8352 13988 8358 14000
rect 8588 13997 8616 14028
rect 9585 14025 9597 14059
rect 9631 14056 9643 14059
rect 9674 14056 9680 14068
rect 9631 14028 9680 14056
rect 9631 14025 9643 14028
rect 9585 14019 9643 14025
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 10410 14016 10416 14068
rect 10468 14056 10474 14068
rect 10781 14059 10839 14065
rect 10781 14056 10793 14059
rect 10468 14028 10793 14056
rect 10468 14016 10474 14028
rect 10781 14025 10793 14028
rect 10827 14025 10839 14059
rect 10781 14019 10839 14025
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 13725 14059 13783 14065
rect 13725 14056 13737 14059
rect 12492 14028 13737 14056
rect 12492 14016 12498 14028
rect 13725 14025 13737 14028
rect 13771 14025 13783 14059
rect 13725 14019 13783 14025
rect 16942 14016 16948 14068
rect 17000 14016 17006 14068
rect 17405 14059 17463 14065
rect 17405 14025 17417 14059
rect 17451 14056 17463 14059
rect 17678 14056 17684 14068
rect 17451 14028 17684 14056
rect 17451 14025 17463 14028
rect 17405 14019 17463 14025
rect 17678 14016 17684 14028
rect 17736 14016 17742 14068
rect 8481 13991 8539 13997
rect 8481 13988 8493 13991
rect 8352 13960 8493 13988
rect 8352 13948 8358 13960
rect 8481 13957 8493 13960
rect 8527 13957 8539 13991
rect 8481 13951 8539 13957
rect 8573 13991 8631 13997
rect 8573 13957 8585 13991
rect 8619 13957 8631 13991
rect 9490 13988 9496 14000
rect 8573 13951 8631 13957
rect 8772 13960 9496 13988
rect 1302 13880 1308 13932
rect 1360 13920 1366 13932
rect 1397 13923 1455 13929
rect 1397 13920 1409 13923
rect 1360 13892 1409 13920
rect 1360 13880 1366 13892
rect 1397 13889 1409 13892
rect 1443 13920 1455 13923
rect 1673 13923 1731 13929
rect 1673 13920 1685 13923
rect 1443 13892 1685 13920
rect 1443 13889 1455 13892
rect 1397 13883 1455 13889
rect 1673 13889 1685 13892
rect 1719 13889 1731 13923
rect 5445 13923 5503 13929
rect 5445 13920 5457 13923
rect 1673 13883 1731 13889
rect 5000 13892 5457 13920
rect 4890 13744 4896 13796
rect 4948 13784 4954 13796
rect 5000 13784 5028 13892
rect 5445 13889 5457 13892
rect 5491 13889 5503 13923
rect 5445 13883 5503 13889
rect 5902 13880 5908 13932
rect 5960 13920 5966 13932
rect 6641 13923 6699 13929
rect 6641 13920 6653 13923
rect 5960 13892 6653 13920
rect 5960 13880 5966 13892
rect 6641 13889 6653 13892
rect 6687 13889 6699 13923
rect 6641 13883 6699 13889
rect 6822 13880 6828 13932
rect 6880 13880 6886 13932
rect 7009 13923 7067 13929
rect 7009 13889 7021 13923
rect 7055 13920 7067 13923
rect 7190 13920 7196 13932
rect 7055 13892 7196 13920
rect 7055 13889 7067 13892
rect 7009 13883 7067 13889
rect 7190 13880 7196 13892
rect 7248 13920 7254 13932
rect 8772 13929 8800 13960
rect 9490 13948 9496 13960
rect 9548 13948 9554 14000
rect 7285 13923 7343 13929
rect 7285 13920 7297 13923
rect 7248 13892 7297 13920
rect 7248 13880 7254 13892
rect 7285 13889 7297 13892
rect 7331 13889 7343 13923
rect 7285 13883 7343 13889
rect 7653 13923 7711 13929
rect 7653 13889 7665 13923
rect 7699 13920 7711 13923
rect 8389 13923 8447 13929
rect 8389 13920 8401 13923
rect 7699 13892 8401 13920
rect 7699 13889 7711 13892
rect 7653 13883 7711 13889
rect 8389 13889 8401 13892
rect 8435 13889 8447 13923
rect 8389 13883 8447 13889
rect 8757 13923 8815 13929
rect 8757 13889 8769 13923
rect 8803 13889 8815 13923
rect 8757 13883 8815 13889
rect 8846 13880 8852 13932
rect 8904 13880 8910 13932
rect 9769 13923 9827 13929
rect 9769 13889 9781 13923
rect 9815 13920 9827 13923
rect 10428 13920 10456 14016
rect 13081 13991 13139 13997
rect 11072 13960 12664 13988
rect 11072 13932 11100 13960
rect 9815 13892 10456 13920
rect 9815 13889 9827 13892
rect 9769 13883 9827 13889
rect 11054 13880 11060 13932
rect 11112 13880 11118 13932
rect 11241 13923 11299 13929
rect 11241 13889 11253 13923
rect 11287 13920 11299 13923
rect 11514 13920 11520 13932
rect 11287 13892 11520 13920
rect 11287 13889 11299 13892
rect 11241 13883 11299 13889
rect 11514 13880 11520 13892
rect 11572 13880 11578 13932
rect 11606 13880 11612 13932
rect 11664 13880 11670 13932
rect 12084 13929 12112 13960
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13889 11943 13923
rect 11885 13883 11943 13889
rect 12069 13923 12127 13929
rect 12069 13889 12081 13923
rect 12115 13889 12127 13923
rect 12069 13883 12127 13889
rect 12345 13923 12403 13929
rect 12345 13889 12357 13923
rect 12391 13920 12403 13923
rect 12526 13920 12532 13932
rect 12391 13892 12532 13920
rect 12391 13889 12403 13892
rect 12345 13883 12403 13889
rect 5261 13855 5319 13861
rect 5261 13821 5273 13855
rect 5307 13821 5319 13855
rect 8662 13852 8668 13864
rect 5261 13815 5319 13821
rect 8220 13824 8668 13852
rect 4948 13756 5028 13784
rect 4948 13744 4954 13756
rect 1578 13676 1584 13728
rect 1636 13676 1642 13728
rect 5276 13716 5304 13815
rect 8220 13793 8248 13824
rect 8662 13812 8668 13824
rect 8720 13812 8726 13864
rect 9953 13855 10011 13861
rect 9953 13821 9965 13855
rect 9999 13852 10011 13855
rect 9999 13824 10916 13852
rect 9999 13821 10011 13824
rect 9953 13815 10011 13821
rect 8205 13787 8263 13793
rect 8205 13753 8217 13787
rect 8251 13753 8263 13787
rect 10888 13784 10916 13824
rect 10962 13812 10968 13864
rect 11020 13812 11026 13864
rect 11149 13855 11207 13861
rect 11149 13821 11161 13855
rect 11195 13852 11207 13855
rect 11900 13852 11928 13883
rect 12526 13880 12532 13892
rect 12584 13880 12590 13932
rect 12636 13929 12664 13960
rect 13081 13957 13093 13991
rect 13127 13988 13139 13991
rect 15746 13988 15752 14000
rect 13127 13960 15752 13988
rect 13127 13957 13139 13960
rect 13081 13951 13139 13957
rect 15746 13948 15752 13960
rect 15804 13988 15810 14000
rect 16390 13988 16396 14000
rect 15804 13960 16396 13988
rect 15804 13948 15810 13960
rect 12621 13923 12679 13929
rect 12621 13889 12633 13923
rect 12667 13889 12679 13923
rect 12621 13883 12679 13889
rect 12986 13880 12992 13932
rect 13044 13920 13050 13932
rect 13541 13923 13599 13929
rect 13541 13920 13553 13923
rect 13044 13892 13553 13920
rect 13044 13880 13050 13892
rect 13541 13889 13553 13892
rect 13587 13889 13599 13923
rect 13541 13883 13599 13889
rect 13630 13880 13636 13932
rect 13688 13880 13694 13932
rect 14458 13880 14464 13932
rect 14516 13880 14522 13932
rect 15286 13880 15292 13932
rect 15344 13920 15350 13932
rect 15841 13923 15899 13929
rect 15841 13920 15853 13923
rect 15344 13892 15853 13920
rect 15344 13880 15350 13892
rect 15841 13889 15853 13892
rect 15887 13889 15899 13923
rect 15841 13883 15899 13889
rect 16022 13880 16028 13932
rect 16080 13880 16086 13932
rect 16132 13929 16160 13960
rect 16390 13948 16396 13960
rect 16448 13948 16454 14000
rect 16117 13923 16175 13929
rect 16117 13889 16129 13923
rect 16163 13889 16175 13923
rect 16117 13883 16175 13889
rect 16206 13880 16212 13932
rect 16264 13880 16270 13932
rect 17034 13880 17040 13932
rect 17092 13880 17098 13932
rect 12250 13852 12256 13864
rect 11195 13824 12256 13852
rect 11195 13821 11207 13824
rect 11149 13815 11207 13821
rect 12250 13812 12256 13824
rect 12308 13812 12314 13864
rect 12434 13812 12440 13864
rect 12492 13812 12498 13864
rect 11606 13784 11612 13796
rect 10888 13756 11612 13784
rect 8205 13747 8263 13753
rect 11606 13744 11612 13756
rect 11664 13744 11670 13796
rect 12544 13784 12572 13880
rect 12710 13812 12716 13864
rect 12768 13852 12774 13864
rect 13265 13855 13323 13861
rect 13265 13852 13277 13855
rect 12768 13824 13277 13852
rect 12768 13812 12774 13824
rect 13265 13821 13277 13824
rect 13311 13852 13323 13855
rect 13357 13855 13415 13861
rect 13357 13852 13369 13855
rect 13311 13824 13369 13852
rect 13311 13821 13323 13824
rect 13265 13815 13323 13821
rect 13357 13821 13369 13824
rect 13403 13821 13415 13855
rect 13357 13815 13415 13821
rect 14366 13812 14372 13864
rect 14424 13812 14430 13864
rect 15197 13855 15255 13861
rect 15197 13821 15209 13855
rect 15243 13821 15255 13855
rect 15197 13815 15255 13821
rect 12406 13756 12572 13784
rect 5626 13716 5632 13728
rect 5276 13688 5632 13716
rect 5626 13676 5632 13688
rect 5684 13676 5690 13728
rect 5810 13676 5816 13728
rect 5868 13676 5874 13728
rect 10962 13676 10968 13728
rect 11020 13716 11026 13728
rect 12406 13716 12434 13756
rect 12618 13744 12624 13796
rect 12676 13784 12682 13796
rect 14274 13784 14280 13796
rect 12676 13756 14280 13784
rect 12676 13744 12682 13756
rect 14274 13744 14280 13756
rect 14332 13784 14338 13796
rect 15212 13784 15240 13815
rect 16482 13812 16488 13864
rect 16540 13812 16546 13864
rect 16853 13855 16911 13861
rect 16853 13821 16865 13855
rect 16899 13821 16911 13855
rect 16853 13815 16911 13821
rect 16574 13784 16580 13796
rect 14332 13756 14872 13784
rect 15212 13756 16580 13784
rect 14332 13744 14338 13756
rect 11020 13688 12434 13716
rect 13909 13719 13967 13725
rect 11020 13676 11026 13688
rect 13909 13685 13921 13719
rect 13955 13716 13967 13719
rect 13998 13716 14004 13728
rect 13955 13688 14004 13716
rect 13955 13685 13967 13688
rect 13909 13679 13967 13685
rect 13998 13676 14004 13688
rect 14056 13676 14062 13728
rect 14844 13716 14872 13756
rect 16574 13744 16580 13756
rect 16632 13744 16638 13796
rect 16868 13784 16896 13815
rect 17310 13784 17316 13796
rect 16868 13756 17316 13784
rect 17310 13744 17316 13756
rect 17368 13784 17374 13796
rect 17770 13784 17776 13796
rect 17368 13756 17776 13784
rect 17368 13744 17374 13756
rect 17770 13744 17776 13756
rect 17828 13744 17834 13796
rect 17862 13716 17868 13728
rect 14844 13688 17868 13716
rect 17862 13676 17868 13688
rect 17920 13676 17926 13728
rect 1104 13626 18860 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 18860 13626
rect 1104 13552 18860 13574
rect 4341 13515 4399 13521
rect 4341 13481 4353 13515
rect 4387 13512 4399 13515
rect 4890 13512 4896 13524
rect 4387 13484 4896 13512
rect 4387 13481 4399 13484
rect 4341 13475 4399 13481
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 5902 13472 5908 13524
rect 5960 13472 5966 13524
rect 6457 13515 6515 13521
rect 6457 13481 6469 13515
rect 6503 13512 6515 13515
rect 6822 13512 6828 13524
rect 6503 13484 6828 13512
rect 6503 13481 6515 13484
rect 6457 13475 6515 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 13633 13515 13691 13521
rect 13633 13481 13645 13515
rect 13679 13512 13691 13515
rect 14182 13512 14188 13524
rect 13679 13484 14188 13512
rect 13679 13481 13691 13484
rect 13633 13475 13691 13481
rect 14182 13472 14188 13484
rect 14240 13472 14246 13524
rect 14274 13472 14280 13524
rect 14332 13472 14338 13524
rect 14366 13472 14372 13524
rect 14424 13512 14430 13524
rect 14461 13515 14519 13521
rect 14461 13512 14473 13515
rect 14424 13484 14473 13512
rect 14424 13472 14430 13484
rect 14461 13481 14473 13484
rect 14507 13481 14519 13515
rect 14461 13475 14519 13481
rect 14645 13515 14703 13521
rect 14645 13481 14657 13515
rect 14691 13512 14703 13515
rect 15654 13512 15660 13524
rect 14691 13484 15660 13512
rect 14691 13481 14703 13484
rect 14645 13475 14703 13481
rect 8662 13404 8668 13456
rect 8720 13444 8726 13456
rect 8938 13444 8944 13456
rect 8720 13416 8944 13444
rect 8720 13404 8726 13416
rect 8938 13404 8944 13416
rect 8996 13444 9002 13456
rect 9398 13444 9404 13456
rect 8996 13416 9404 13444
rect 8996 13404 9002 13416
rect 9398 13404 9404 13416
rect 9456 13404 9462 13456
rect 14660 13444 14688 13475
rect 15654 13472 15660 13484
rect 15712 13512 15718 13524
rect 16577 13515 16635 13521
rect 15712 13484 16252 13512
rect 15712 13472 15718 13484
rect 16224 13456 16252 13484
rect 16577 13481 16589 13515
rect 16623 13512 16635 13515
rect 17034 13512 17040 13524
rect 16623 13484 17040 13512
rect 16623 13481 16635 13484
rect 16577 13475 16635 13481
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 13924 13416 14688 13444
rect 4062 13336 4068 13388
rect 4120 13336 4126 13388
rect 12713 13379 12771 13385
rect 12713 13345 12725 13379
rect 12759 13376 12771 13379
rect 12894 13376 12900 13388
rect 12759 13348 12900 13376
rect 12759 13345 12771 13348
rect 12713 13339 12771 13345
rect 12894 13336 12900 13348
rect 12952 13336 12958 13388
rect 12986 13336 12992 13388
rect 13044 13336 13050 13388
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13308 4031 13311
rect 4798 13308 4804 13320
rect 4019 13280 4804 13308
rect 4019 13277 4031 13280
rect 3973 13271 4031 13277
rect 4798 13268 4804 13280
rect 4856 13268 4862 13320
rect 5442 13268 5448 13320
rect 5500 13268 5506 13320
rect 5718 13268 5724 13320
rect 5776 13268 5782 13320
rect 8386 13268 8392 13320
rect 8444 13308 8450 13320
rect 8570 13308 8576 13320
rect 8444 13280 8576 13308
rect 8444 13268 8450 13280
rect 8570 13268 8576 13280
rect 8628 13268 8634 13320
rect 13354 13268 13360 13320
rect 13412 13308 13418 13320
rect 13924 13317 13952 13416
rect 15470 13404 15476 13456
rect 15528 13444 15534 13456
rect 16022 13444 16028 13456
rect 15528 13416 16028 13444
rect 15528 13404 15534 13416
rect 16022 13404 16028 13416
rect 16080 13404 16086 13456
rect 16206 13404 16212 13456
rect 16264 13444 16270 13456
rect 16264 13416 17816 13444
rect 16264 13404 16270 13416
rect 13998 13336 14004 13388
rect 14056 13376 14062 13388
rect 17788 13385 17816 13416
rect 17129 13379 17187 13385
rect 17129 13376 17141 13379
rect 14056 13348 17141 13376
rect 14056 13336 14062 13348
rect 14752 13317 14780 13348
rect 17129 13345 17141 13348
rect 17175 13345 17187 13379
rect 17129 13339 17187 13345
rect 17773 13379 17831 13385
rect 17773 13345 17785 13379
rect 17819 13345 17831 13379
rect 17773 13339 17831 13345
rect 18046 13336 18052 13388
rect 18104 13376 18110 13388
rect 18233 13379 18291 13385
rect 18233 13376 18245 13379
rect 18104 13348 18245 13376
rect 18104 13336 18110 13348
rect 18233 13345 18245 13348
rect 18279 13345 18291 13379
rect 18233 13339 18291 13345
rect 13633 13311 13691 13317
rect 13633 13308 13645 13311
rect 13412 13280 13645 13308
rect 13412 13268 13418 13280
rect 13633 13277 13645 13280
rect 13679 13277 13691 13311
rect 13633 13271 13691 13277
rect 13909 13311 13967 13317
rect 13909 13277 13921 13311
rect 13955 13308 13967 13311
rect 14737 13311 14795 13317
rect 13955 13280 14320 13308
rect 13955 13277 13967 13280
rect 13909 13271 13967 13277
rect 5460 13240 5488 13268
rect 6089 13243 6147 13249
rect 6089 13240 6101 13243
rect 5460 13212 6101 13240
rect 6089 13209 6101 13212
rect 6135 13209 6147 13243
rect 6089 13203 6147 13209
rect 6273 13243 6331 13249
rect 6273 13209 6285 13243
rect 6319 13209 6331 13243
rect 6273 13203 6331 13209
rect 8665 13243 8723 13249
rect 8665 13209 8677 13243
rect 8711 13209 8723 13243
rect 13648 13240 13676 13271
rect 14093 13243 14151 13249
rect 14093 13240 14105 13243
rect 13648 13212 14105 13240
rect 8665 13203 8723 13209
rect 14093 13209 14105 13212
rect 14139 13209 14151 13243
rect 14093 13203 14151 13209
rect 5534 13132 5540 13184
rect 5592 13172 5598 13184
rect 6288 13172 6316 13203
rect 5592 13144 6316 13172
rect 5592 13132 5598 13144
rect 8478 13132 8484 13184
rect 8536 13132 8542 13184
rect 8680 13172 8708 13203
rect 14182 13200 14188 13252
rect 14240 13200 14246 13252
rect 14292 13249 14320 13280
rect 14737 13277 14749 13311
rect 14783 13277 14795 13311
rect 14737 13271 14795 13277
rect 15286 13268 15292 13320
rect 15344 13308 15350 13320
rect 15381 13311 15439 13317
rect 15381 13308 15393 13311
rect 15344 13280 15393 13308
rect 15344 13268 15350 13280
rect 15381 13277 15393 13280
rect 15427 13277 15439 13311
rect 15381 13271 15439 13277
rect 14292 13243 14351 13249
rect 14292 13212 14305 13243
rect 14293 13209 14305 13212
rect 14339 13209 14351 13243
rect 14293 13203 14351 13209
rect 14550 13200 14556 13252
rect 14608 13240 14614 13252
rect 15396 13240 15424 13271
rect 15470 13268 15476 13320
rect 15528 13268 15534 13320
rect 15654 13268 15660 13320
rect 15712 13268 15718 13320
rect 15746 13268 15752 13320
rect 15804 13268 15810 13320
rect 16022 13268 16028 13320
rect 16080 13308 16086 13320
rect 16209 13311 16267 13317
rect 16209 13308 16221 13311
rect 16080 13280 16221 13308
rect 16080 13268 16086 13280
rect 16209 13277 16221 13280
rect 16255 13277 16267 13311
rect 16209 13271 16267 13277
rect 16393 13311 16451 13317
rect 16393 13277 16405 13311
rect 16439 13277 16451 13311
rect 16393 13271 16451 13277
rect 17221 13311 17279 13317
rect 17221 13277 17233 13311
rect 17267 13277 17279 13311
rect 17221 13271 17279 13277
rect 16408 13240 16436 13271
rect 14608 13212 15332 13240
rect 15396 13212 16436 13240
rect 14608 13200 14614 13212
rect 8754 13172 8760 13184
rect 8680 13144 8760 13172
rect 8754 13132 8760 13144
rect 8812 13172 8818 13184
rect 11330 13172 11336 13184
rect 8812 13144 11336 13172
rect 8812 13132 8818 13144
rect 11330 13132 11336 13144
rect 11388 13132 11394 13184
rect 13817 13175 13875 13181
rect 13817 13141 13829 13175
rect 13863 13172 13875 13175
rect 14200 13172 14228 13200
rect 13863 13144 14228 13172
rect 13863 13141 13875 13144
rect 13817 13135 13875 13141
rect 15194 13132 15200 13184
rect 15252 13132 15258 13184
rect 15304 13172 15332 13212
rect 17236 13172 17264 13271
rect 17862 13268 17868 13320
rect 17920 13268 17926 13320
rect 15304 13144 17264 13172
rect 17586 13132 17592 13184
rect 17644 13132 17650 13184
rect 1104 13082 18860 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 18860 13082
rect 1104 13008 18860 13030
rect 7929 12971 7987 12977
rect 7929 12937 7941 12971
rect 7975 12968 7987 12971
rect 8294 12968 8300 12980
rect 7975 12940 8300 12968
rect 7975 12937 7987 12940
rect 7929 12931 7987 12937
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 8573 12971 8631 12977
rect 8573 12937 8585 12971
rect 8619 12968 8631 12971
rect 8846 12968 8852 12980
rect 8619 12940 8852 12968
rect 8619 12937 8631 12940
rect 8573 12931 8631 12937
rect 8846 12928 8852 12940
rect 8904 12928 8910 12980
rect 14918 12928 14924 12980
rect 14976 12968 14982 12980
rect 15378 12968 15384 12980
rect 14976 12940 15384 12968
rect 14976 12928 14982 12940
rect 15378 12928 15384 12940
rect 15436 12928 15442 12980
rect 9122 12900 9128 12912
rect 8128 12872 9128 12900
rect 1302 12792 1308 12844
rect 1360 12832 1366 12844
rect 1397 12835 1455 12841
rect 1397 12832 1409 12835
rect 1360 12804 1409 12832
rect 1360 12792 1366 12804
rect 1397 12801 1409 12804
rect 1443 12832 1455 12835
rect 1673 12835 1731 12841
rect 1673 12832 1685 12835
rect 1443 12804 1685 12832
rect 1443 12801 1455 12804
rect 1397 12795 1455 12801
rect 1673 12801 1685 12804
rect 1719 12801 1731 12835
rect 1673 12795 1731 12801
rect 5442 12792 5448 12844
rect 5500 12832 5506 12844
rect 8128 12841 8156 12872
rect 9122 12860 9128 12872
rect 9180 12900 9186 12912
rect 12986 12900 12992 12912
rect 9180 12872 9260 12900
rect 9180 12860 9186 12872
rect 5997 12835 6055 12841
rect 5997 12832 6009 12835
rect 5500 12804 6009 12832
rect 5500 12792 5506 12804
rect 5997 12801 6009 12804
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 8113 12835 8171 12841
rect 8113 12801 8125 12835
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 8205 12835 8263 12841
rect 8205 12801 8217 12835
rect 8251 12801 8263 12835
rect 8205 12795 8263 12801
rect 1581 12699 1639 12705
rect 1581 12665 1593 12699
rect 1627 12696 1639 12699
rect 8220 12696 8248 12795
rect 8294 12792 8300 12844
rect 8352 12841 8358 12844
rect 8846 12841 8852 12844
rect 8352 12836 8406 12841
rect 8352 12835 8432 12836
rect 8352 12801 8360 12835
rect 8394 12804 8432 12835
rect 8829 12835 8852 12841
rect 8481 12825 8539 12831
rect 8394 12801 8406 12804
rect 8352 12795 8406 12801
rect 8352 12792 8358 12795
rect 8481 12791 8493 12825
rect 8527 12822 8539 12825
rect 8527 12794 8600 12822
rect 8829 12801 8841 12835
rect 8829 12795 8852 12801
rect 8527 12791 8539 12794
rect 8481 12785 8539 12791
rect 8572 12764 8600 12794
rect 8846 12792 8852 12795
rect 8904 12792 8910 12844
rect 8938 12835 8996 12841
rect 8938 12828 8950 12835
rect 8984 12828 8996 12835
rect 9038 12838 9096 12844
rect 9232 12841 9260 12872
rect 10612 12872 12992 12900
rect 10612 12841 10640 12872
rect 8938 12776 8944 12828
rect 8996 12776 9002 12828
rect 9038 12804 9050 12838
rect 9084 12804 9096 12838
rect 9038 12798 9096 12804
rect 9217 12835 9275 12841
rect 9217 12801 9229 12835
rect 9263 12832 9275 12835
rect 10413 12835 10471 12841
rect 10413 12832 10425 12835
rect 9263 12804 10425 12832
rect 9263 12801 9275 12804
rect 8662 12764 8668 12776
rect 8572 12736 8668 12764
rect 8662 12724 8668 12736
rect 8720 12724 8726 12776
rect 9048 12764 9076 12798
rect 9217 12795 9275 12801
rect 10413 12801 10425 12804
rect 10459 12801 10471 12835
rect 10413 12795 10471 12801
rect 10597 12835 10655 12841
rect 10597 12801 10609 12835
rect 10643 12801 10655 12835
rect 10597 12795 10655 12801
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 10796 12764 10824 12795
rect 10870 12792 10876 12844
rect 10928 12792 10934 12844
rect 10980 12841 11008 12872
rect 12986 12860 12992 12872
rect 13044 12860 13050 12912
rect 14366 12860 14372 12912
rect 14424 12900 14430 12912
rect 15013 12903 15071 12909
rect 15013 12900 15025 12903
rect 14424 12872 15025 12900
rect 14424 12860 14430 12872
rect 15013 12869 15025 12872
rect 15059 12900 15071 12903
rect 15562 12900 15568 12912
rect 15059 12872 15568 12900
rect 15059 12869 15071 12872
rect 15013 12863 15071 12869
rect 15562 12860 15568 12872
rect 15620 12900 15626 12912
rect 15657 12903 15715 12909
rect 15657 12900 15669 12903
rect 15620 12872 15669 12900
rect 15620 12860 15626 12872
rect 15657 12869 15669 12872
rect 15703 12869 15715 12903
rect 15657 12863 15715 12869
rect 15930 12860 15936 12912
rect 15988 12900 15994 12912
rect 16025 12903 16083 12909
rect 16025 12900 16037 12903
rect 15988 12872 16037 12900
rect 15988 12860 15994 12872
rect 16025 12869 16037 12872
rect 16071 12869 16083 12903
rect 16025 12863 16083 12869
rect 10965 12835 11023 12841
rect 10965 12801 10977 12835
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 11057 12835 11115 12841
rect 11057 12801 11069 12835
rect 11103 12801 11115 12835
rect 11057 12795 11115 12801
rect 11072 12764 11100 12795
rect 11146 12792 11152 12844
rect 11204 12832 11210 12844
rect 11241 12835 11299 12841
rect 11241 12832 11253 12835
rect 11204 12804 11253 12832
rect 11204 12792 11210 12804
rect 11241 12801 11253 12804
rect 11287 12801 11299 12835
rect 11241 12795 11299 12801
rect 14918 12792 14924 12844
rect 14976 12792 14982 12844
rect 15177 12838 15235 12841
rect 15120 12835 15240 12838
rect 15120 12810 15189 12835
rect 9048 12736 9142 12764
rect 10796 12736 11100 12764
rect 9114 12696 9142 12736
rect 9306 12696 9312 12708
rect 1627 12668 6592 12696
rect 8220 12668 9312 12696
rect 1627 12665 1639 12668
rect 1581 12659 1639 12665
rect 6086 12588 6092 12640
rect 6144 12588 6150 12640
rect 6564 12628 6592 12668
rect 9306 12656 9312 12668
rect 9364 12696 9370 12708
rect 10965 12699 11023 12705
rect 10965 12696 10977 12699
rect 9364 12668 10977 12696
rect 9364 12656 9370 12668
rect 10965 12665 10977 12668
rect 11011 12665 11023 12699
rect 10965 12659 11023 12665
rect 10318 12628 10324 12640
rect 6564 12600 10324 12628
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 11072 12628 11100 12736
rect 11330 12724 11336 12776
rect 11388 12764 11394 12776
rect 15120 12764 15148 12810
rect 15177 12801 15189 12810
rect 15223 12804 15240 12835
rect 15223 12801 15235 12804
rect 15177 12795 15235 12801
rect 15378 12792 15384 12844
rect 15436 12832 15442 12844
rect 15473 12835 15531 12841
rect 15473 12832 15485 12835
rect 15436 12804 15485 12832
rect 15436 12792 15442 12804
rect 15473 12801 15485 12804
rect 15519 12801 15531 12835
rect 15473 12795 15531 12801
rect 15749 12835 15807 12841
rect 15749 12801 15761 12835
rect 15795 12801 15807 12835
rect 15749 12795 15807 12801
rect 18049 12835 18107 12841
rect 18049 12801 18061 12835
rect 18095 12832 18107 12835
rect 18138 12832 18144 12844
rect 18095 12804 18144 12832
rect 18095 12801 18107 12804
rect 18049 12795 18107 12801
rect 15764 12764 15792 12795
rect 18138 12792 18144 12804
rect 18196 12792 18202 12844
rect 15841 12767 15899 12773
rect 15841 12764 15853 12767
rect 11388 12736 15853 12764
rect 11388 12724 11394 12736
rect 15841 12733 15853 12736
rect 15887 12733 15899 12767
rect 15841 12727 15899 12733
rect 18322 12724 18328 12776
rect 18380 12724 18386 12776
rect 12250 12628 12256 12640
rect 11072 12600 12256 12628
rect 12250 12588 12256 12600
rect 12308 12628 12314 12640
rect 13630 12628 13636 12640
rect 12308 12600 13636 12628
rect 12308 12588 12314 12600
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 15381 12631 15439 12637
rect 15381 12597 15393 12631
rect 15427 12628 15439 12631
rect 15654 12628 15660 12640
rect 15427 12600 15660 12628
rect 15427 12597 15439 12600
rect 15381 12591 15439 12597
rect 15654 12588 15660 12600
rect 15712 12588 15718 12640
rect 15746 12588 15752 12640
rect 15804 12588 15810 12640
rect 1104 12538 18860 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 18860 12538
rect 1104 12464 18860 12486
rect 6730 12384 6736 12436
rect 6788 12424 6794 12436
rect 8478 12424 8484 12436
rect 6788 12396 8484 12424
rect 6788 12384 6794 12396
rect 8478 12384 8484 12396
rect 8536 12424 8542 12436
rect 8573 12427 8631 12433
rect 8573 12424 8585 12427
rect 8536 12396 8585 12424
rect 8536 12384 8542 12396
rect 8573 12393 8585 12396
rect 8619 12393 8631 12427
rect 8573 12387 8631 12393
rect 8662 12384 8668 12436
rect 8720 12424 8726 12436
rect 10870 12424 10876 12436
rect 8720 12396 10876 12424
rect 8720 12384 8726 12396
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 12437 12427 12495 12433
rect 12437 12393 12449 12427
rect 12483 12424 12495 12427
rect 13262 12424 13268 12436
rect 12483 12396 13268 12424
rect 12483 12393 12495 12396
rect 12437 12387 12495 12393
rect 13262 12384 13268 12396
rect 13320 12384 13326 12436
rect 13357 12427 13415 12433
rect 13357 12393 13369 12427
rect 13403 12424 13415 12427
rect 13630 12424 13636 12436
rect 13403 12396 13636 12424
rect 13403 12393 13415 12396
rect 13357 12387 13415 12393
rect 13630 12384 13636 12396
rect 13688 12384 13694 12436
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 5074 12356 5080 12368
rect 4120 12328 5080 12356
rect 4120 12316 4126 12328
rect 5074 12316 5080 12328
rect 5132 12316 5138 12368
rect 5353 12359 5411 12365
rect 5353 12325 5365 12359
rect 5399 12356 5411 12359
rect 5399 12328 6960 12356
rect 5399 12325 5411 12328
rect 5353 12319 5411 12325
rect 4430 12248 4436 12300
rect 4488 12248 4494 12300
rect 5626 12248 5632 12300
rect 5684 12288 5690 12300
rect 5994 12288 6000 12300
rect 5684 12260 6000 12288
rect 5684 12248 5690 12260
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 6086 12248 6092 12300
rect 6144 12248 6150 12300
rect 6932 12297 6960 12328
rect 8294 12316 8300 12368
rect 8352 12356 8358 12368
rect 8389 12359 8447 12365
rect 8389 12356 8401 12359
rect 8352 12328 8401 12356
rect 8352 12316 8358 12328
rect 8389 12325 8401 12328
rect 8435 12356 8447 12359
rect 8846 12356 8852 12368
rect 8435 12328 8852 12356
rect 8435 12325 8447 12328
rect 8389 12319 8447 12325
rect 8846 12316 8852 12328
rect 8904 12356 8910 12368
rect 13081 12359 13139 12365
rect 8904 12328 9628 12356
rect 8904 12316 8910 12328
rect 6917 12291 6975 12297
rect 6917 12257 6929 12291
rect 6963 12288 6975 12291
rect 8662 12288 8668 12300
rect 6963 12260 8668 12288
rect 6963 12257 6975 12260
rect 6917 12251 6975 12257
rect 8662 12248 8668 12260
rect 8720 12248 8726 12300
rect 9306 12248 9312 12300
rect 9364 12248 9370 12300
rect 3786 12180 3792 12232
rect 3844 12220 3850 12232
rect 4341 12223 4399 12229
rect 4341 12220 4353 12223
rect 3844 12192 4353 12220
rect 3844 12180 3850 12192
rect 4341 12189 4353 12192
rect 4387 12220 4399 12223
rect 5169 12223 5227 12229
rect 5169 12220 5181 12223
rect 4387 12192 5181 12220
rect 4387 12189 4399 12192
rect 4341 12183 4399 12189
rect 5169 12189 5181 12192
rect 5215 12189 5227 12223
rect 5169 12183 5227 12189
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12220 6883 12223
rect 6871 12192 9076 12220
rect 6871 12189 6883 12192
rect 6825 12183 6883 12189
rect 4246 12112 4252 12164
rect 4304 12152 4310 12164
rect 4801 12155 4859 12161
rect 4801 12152 4813 12155
rect 4304 12124 4813 12152
rect 4304 12112 4310 12124
rect 4801 12121 4813 12124
rect 4847 12121 4859 12155
rect 5534 12152 5540 12164
rect 4801 12115 4859 12121
rect 4908 12124 5540 12152
rect 4709 12087 4767 12093
rect 4709 12053 4721 12087
rect 4755 12084 4767 12087
rect 4908 12084 4936 12124
rect 5534 12112 5540 12124
rect 5592 12152 5598 12164
rect 6181 12155 6239 12161
rect 6181 12152 6193 12155
rect 5592 12124 6193 12152
rect 5592 12112 5598 12124
rect 6181 12121 6193 12124
rect 6227 12121 6239 12155
rect 6181 12115 6239 12121
rect 8754 12112 8760 12164
rect 8812 12112 8818 12164
rect 9048 12152 9076 12192
rect 9122 12180 9128 12232
rect 9180 12180 9186 12232
rect 9398 12180 9404 12232
rect 9456 12180 9462 12232
rect 9600 12229 9628 12328
rect 13081 12325 13093 12359
rect 13127 12356 13139 12359
rect 13998 12356 14004 12368
rect 13127 12328 14004 12356
rect 13127 12325 13139 12328
rect 13081 12319 13139 12325
rect 13998 12316 14004 12328
rect 14056 12316 14062 12368
rect 11333 12291 11391 12297
rect 11333 12257 11345 12291
rect 11379 12288 11391 12291
rect 12805 12291 12863 12297
rect 11379 12260 12204 12288
rect 11379 12257 11391 12260
rect 11333 12251 11391 12257
rect 12176 12229 12204 12260
rect 12805 12257 12817 12291
rect 12851 12288 12863 12291
rect 14918 12288 14924 12300
rect 12851 12260 14924 12288
rect 12851 12257 12863 12260
rect 12805 12251 12863 12257
rect 14918 12248 14924 12260
rect 14976 12248 14982 12300
rect 16482 12248 16488 12300
rect 16540 12288 16546 12300
rect 16540 12260 17448 12288
rect 16540 12248 16546 12260
rect 9585 12223 9643 12229
rect 9585 12189 9597 12223
rect 9631 12189 9643 12223
rect 9585 12183 9643 12189
rect 11241 12223 11299 12229
rect 11241 12189 11253 12223
rect 11287 12189 11299 12223
rect 11241 12183 11299 12189
rect 11885 12223 11943 12229
rect 11885 12189 11897 12223
rect 11931 12189 11943 12223
rect 11885 12183 11943 12189
rect 12161 12223 12219 12229
rect 12161 12189 12173 12223
rect 12207 12220 12219 12223
rect 12526 12220 12532 12232
rect 12207 12192 12532 12220
rect 12207 12189 12219 12192
rect 12161 12183 12219 12189
rect 11256 12152 11284 12183
rect 11793 12155 11851 12161
rect 11793 12152 11805 12155
rect 9048 12124 11805 12152
rect 11793 12121 11805 12124
rect 11839 12121 11851 12155
rect 11900 12152 11928 12183
rect 12526 12180 12532 12192
rect 12584 12180 12590 12232
rect 12713 12223 12771 12229
rect 12713 12189 12725 12223
rect 12759 12220 12771 12223
rect 14366 12220 14372 12232
rect 12759 12192 14372 12220
rect 12759 12189 12771 12192
rect 12713 12183 12771 12189
rect 14366 12180 14372 12192
rect 14424 12180 14430 12232
rect 17126 12180 17132 12232
rect 17184 12180 17190 12232
rect 17420 12229 17448 12260
rect 17405 12223 17463 12229
rect 17405 12189 17417 12223
rect 17451 12189 17463 12223
rect 17405 12183 17463 12189
rect 17586 12180 17592 12232
rect 17644 12220 17650 12232
rect 17865 12223 17923 12229
rect 17865 12220 17877 12223
rect 17644 12192 17877 12220
rect 17644 12180 17650 12192
rect 17865 12189 17877 12192
rect 17911 12189 17923 12223
rect 17865 12183 17923 12189
rect 12250 12152 12256 12164
rect 11900 12124 12256 12152
rect 11793 12115 11851 12121
rect 12250 12112 12256 12124
rect 12308 12112 12314 12164
rect 12437 12155 12495 12161
rect 12437 12121 12449 12155
rect 12483 12121 12495 12155
rect 12437 12115 12495 12121
rect 13173 12155 13231 12161
rect 13173 12121 13185 12155
rect 13219 12121 13231 12155
rect 13173 12115 13231 12121
rect 4755 12056 4936 12084
rect 4755 12053 4767 12056
rect 4709 12047 4767 12053
rect 4982 12044 4988 12096
rect 5040 12044 5046 12096
rect 5074 12044 5080 12096
rect 5132 12044 5138 12096
rect 6546 12044 6552 12096
rect 6604 12044 6610 12096
rect 7190 12044 7196 12096
rect 7248 12044 7254 12096
rect 8570 12093 8576 12096
rect 8557 12087 8576 12093
rect 8557 12053 8569 12087
rect 8557 12047 8576 12053
rect 8570 12044 8576 12047
rect 8628 12044 8634 12096
rect 8938 12044 8944 12096
rect 8996 12044 9002 12096
rect 9490 12044 9496 12096
rect 9548 12044 9554 12096
rect 11606 12044 11612 12096
rect 11664 12044 11670 12096
rect 12452 12084 12480 12115
rect 12986 12084 12992 12096
rect 12452 12056 12992 12084
rect 12986 12044 12992 12056
rect 13044 12084 13050 12096
rect 13188 12084 13216 12115
rect 13262 12112 13268 12164
rect 13320 12152 13326 12164
rect 15378 12152 15384 12164
rect 13320 12124 15384 12152
rect 13320 12112 13326 12124
rect 15378 12112 15384 12124
rect 15436 12112 15442 12164
rect 17221 12155 17279 12161
rect 17221 12121 17233 12155
rect 17267 12152 17279 12155
rect 17604 12152 17632 12180
rect 17267 12124 17632 12152
rect 17681 12155 17739 12161
rect 17267 12121 17279 12124
rect 17221 12115 17279 12121
rect 17681 12121 17693 12155
rect 17727 12152 17739 12155
rect 17727 12124 17908 12152
rect 17727 12121 17739 12124
rect 17681 12115 17739 12121
rect 17880 12096 17908 12124
rect 13044 12056 13216 12084
rect 13044 12044 13050 12056
rect 13354 12044 13360 12096
rect 13412 12093 13418 12096
rect 13412 12087 13431 12093
rect 13419 12053 13431 12087
rect 13412 12047 13431 12053
rect 13541 12087 13599 12093
rect 13541 12053 13553 12087
rect 13587 12084 13599 12087
rect 15286 12084 15292 12096
rect 13587 12056 15292 12084
rect 13587 12053 13599 12056
rect 13541 12047 13599 12053
rect 13412 12044 13418 12047
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 17589 12087 17647 12093
rect 17589 12053 17601 12087
rect 17635 12084 17647 12087
rect 17770 12084 17776 12096
rect 17635 12056 17776 12084
rect 17635 12053 17647 12056
rect 17589 12047 17647 12053
rect 17770 12044 17776 12056
rect 17828 12044 17834 12096
rect 17862 12044 17868 12096
rect 17920 12044 17926 12096
rect 18049 12087 18107 12093
rect 18049 12053 18061 12087
rect 18095 12084 18107 12087
rect 18230 12084 18236 12096
rect 18095 12056 18236 12084
rect 18095 12053 18107 12056
rect 18049 12047 18107 12053
rect 18230 12044 18236 12056
rect 18288 12044 18294 12096
rect 1104 11994 18860 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 18860 11994
rect 1104 11920 18860 11942
rect 4246 11840 4252 11892
rect 4304 11840 4310 11892
rect 4430 11840 4436 11892
rect 4488 11840 4494 11892
rect 8481 11883 8539 11889
rect 8481 11849 8493 11883
rect 8527 11880 8539 11883
rect 8938 11880 8944 11892
rect 8527 11852 8944 11880
rect 8527 11849 8539 11852
rect 8481 11843 8539 11849
rect 8938 11840 8944 11852
rect 8996 11840 9002 11892
rect 10689 11883 10747 11889
rect 10689 11849 10701 11883
rect 10735 11880 10747 11883
rect 12526 11880 12532 11892
rect 10735 11852 12532 11880
rect 10735 11849 10747 11852
rect 10689 11843 10747 11849
rect 12526 11840 12532 11852
rect 12584 11880 12590 11892
rect 13354 11880 13360 11892
rect 12584 11852 13360 11880
rect 12584 11840 12590 11852
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 15194 11880 15200 11892
rect 14476 11852 15200 11880
rect 4798 11812 4804 11824
rect 3344 11784 4108 11812
rect 1302 11704 1308 11756
rect 1360 11744 1366 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 1360 11716 1409 11744
rect 1360 11704 1366 11716
rect 1397 11713 1409 11716
rect 1443 11744 1455 11747
rect 1673 11747 1731 11753
rect 1673 11744 1685 11747
rect 1443 11716 1685 11744
rect 1443 11713 1455 11716
rect 1397 11707 1455 11713
rect 1673 11713 1685 11716
rect 1719 11713 1731 11747
rect 1673 11707 1731 11713
rect 3344 11685 3372 11784
rect 4080 11753 4108 11784
rect 4356 11784 4804 11812
rect 4356 11753 4384 11784
rect 4798 11772 4804 11784
rect 4856 11812 4862 11824
rect 8573 11815 8631 11821
rect 4856 11784 8156 11812
rect 4856 11772 4862 11784
rect 3421 11747 3479 11753
rect 3421 11713 3433 11747
rect 3467 11713 3479 11747
rect 3421 11707 3479 11713
rect 4065 11747 4123 11753
rect 4065 11713 4077 11747
rect 4111 11713 4123 11747
rect 4065 11707 4123 11713
rect 4341 11747 4399 11753
rect 4341 11713 4353 11747
rect 4387 11713 4399 11747
rect 4341 11707 4399 11713
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11713 4583 11747
rect 4525 11707 4583 11713
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11744 6607 11747
rect 6730 11744 6736 11756
rect 6595 11716 6736 11744
rect 6595 11713 6607 11716
rect 6549 11707 6607 11713
rect 3329 11679 3387 11685
rect 3329 11645 3341 11679
rect 3375 11645 3387 11679
rect 3329 11639 3387 11645
rect 1581 11611 1639 11617
rect 1581 11577 1593 11611
rect 1627 11608 1639 11611
rect 3344 11608 3372 11639
rect 1627 11580 3372 11608
rect 3436 11608 3464 11707
rect 3786 11636 3792 11688
rect 3844 11636 3850 11688
rect 3881 11679 3939 11685
rect 3881 11645 3893 11679
rect 3927 11645 3939 11679
rect 3881 11639 3939 11645
rect 3896 11608 3924 11639
rect 3970 11636 3976 11688
rect 4028 11676 4034 11688
rect 4540 11676 4568 11707
rect 6730 11704 6736 11716
rect 6788 11704 6794 11756
rect 8128 11744 8156 11784
rect 8573 11781 8585 11815
rect 8619 11812 8631 11815
rect 9490 11812 9496 11824
rect 8619 11784 9496 11812
rect 8619 11781 8631 11784
rect 8573 11775 8631 11781
rect 9490 11772 9496 11784
rect 9548 11772 9554 11824
rect 9784 11784 10456 11812
rect 9784 11744 9812 11784
rect 8128 11716 9812 11744
rect 9861 11747 9919 11753
rect 9861 11713 9873 11747
rect 9907 11713 9919 11747
rect 9861 11707 9919 11713
rect 4028 11648 4568 11676
rect 6641 11679 6699 11685
rect 4028 11636 4034 11648
rect 6641 11645 6653 11679
rect 6687 11676 6699 11679
rect 8570 11676 8576 11688
rect 6687 11648 8576 11676
rect 6687 11645 6699 11648
rect 6641 11639 6699 11645
rect 8570 11636 8576 11648
rect 8628 11636 8634 11688
rect 8754 11636 8760 11688
rect 8812 11676 8818 11688
rect 9214 11676 9220 11688
rect 8812 11648 9220 11676
rect 8812 11636 8818 11648
rect 9214 11636 9220 11648
rect 9272 11636 9278 11688
rect 9674 11636 9680 11688
rect 9732 11636 9738 11688
rect 9306 11608 9312 11620
rect 3436 11580 9312 11608
rect 1627 11577 1639 11580
rect 1581 11571 1639 11577
rect 9306 11568 9312 11580
rect 9364 11608 9370 11620
rect 9876 11608 9904 11707
rect 10318 11704 10324 11756
rect 10376 11704 10382 11756
rect 10428 11753 10456 11784
rect 11606 11772 11612 11824
rect 11664 11812 11670 11824
rect 11664 11784 14228 11812
rect 11664 11772 11670 11784
rect 14200 11756 14228 11784
rect 10413 11747 10471 11753
rect 10413 11713 10425 11747
rect 10459 11744 10471 11747
rect 10686 11744 10692 11756
rect 10459 11716 10692 11744
rect 10459 11713 10471 11716
rect 10413 11707 10471 11713
rect 10686 11704 10692 11716
rect 10744 11704 10750 11756
rect 13998 11704 14004 11756
rect 14056 11704 14062 11756
rect 14182 11704 14188 11756
rect 14240 11704 14246 11756
rect 14476 11753 14504 11852
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 15286 11840 15292 11892
rect 15344 11880 15350 11892
rect 16117 11883 16175 11889
rect 15344 11852 16068 11880
rect 15344 11840 15350 11852
rect 15013 11815 15071 11821
rect 15013 11812 15025 11815
rect 14752 11784 15025 11812
rect 14752 11753 14780 11784
rect 15013 11781 15025 11784
rect 15059 11781 15071 11815
rect 15013 11775 15071 11781
rect 15488 11784 15792 11812
rect 14277 11747 14335 11753
rect 14277 11713 14289 11747
rect 14323 11713 14335 11747
rect 14277 11707 14335 11713
rect 14461 11747 14519 11753
rect 14461 11713 14473 11747
rect 14507 11713 14519 11747
rect 14461 11707 14519 11713
rect 14737 11747 14795 11753
rect 14737 11713 14749 11747
rect 14783 11713 14795 11747
rect 14737 11707 14795 11713
rect 10045 11679 10103 11685
rect 10045 11645 10057 11679
rect 10091 11676 10103 11679
rect 10229 11679 10287 11685
rect 10229 11676 10241 11679
rect 10091 11648 10241 11676
rect 10091 11645 10103 11648
rect 10045 11639 10103 11645
rect 10229 11645 10241 11648
rect 10275 11645 10287 11679
rect 10229 11639 10287 11645
rect 10502 11636 10508 11688
rect 10560 11636 10566 11688
rect 14292 11676 14320 11707
rect 15286 11704 15292 11756
rect 15344 11704 15350 11756
rect 15378 11704 15384 11756
rect 15436 11704 15442 11756
rect 15488 11753 15516 11784
rect 15764 11756 15792 11784
rect 15473 11747 15531 11753
rect 15473 11713 15485 11747
rect 15519 11713 15531 11747
rect 15473 11707 15531 11713
rect 15654 11704 15660 11756
rect 15712 11704 15718 11756
rect 15746 11704 15752 11756
rect 15804 11704 15810 11756
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11713 15991 11747
rect 16040 11744 16068 11852
rect 16117 11849 16129 11883
rect 16163 11880 16175 11883
rect 17037 11883 17095 11889
rect 17037 11880 17049 11883
rect 16163 11852 17049 11880
rect 16163 11849 16175 11852
rect 16117 11843 16175 11849
rect 17037 11849 17049 11852
rect 17083 11849 17095 11883
rect 17037 11843 17095 11849
rect 17126 11840 17132 11892
rect 17184 11880 17190 11892
rect 17862 11880 17868 11892
rect 17184 11852 17868 11880
rect 17184 11840 17190 11852
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 16301 11815 16359 11821
rect 16301 11781 16313 11815
rect 16347 11812 16359 11815
rect 16945 11815 17003 11821
rect 16945 11812 16957 11815
rect 16347 11784 16957 11812
rect 16347 11781 16359 11784
rect 16301 11775 16359 11781
rect 16945 11781 16957 11784
rect 16991 11781 17003 11815
rect 16945 11775 17003 11781
rect 17954 11772 17960 11824
rect 18012 11772 18018 11824
rect 16390 11753 16396 11756
rect 16209 11747 16267 11753
rect 16209 11744 16221 11747
rect 16040 11716 16221 11744
rect 15933 11707 15991 11713
rect 16209 11713 16221 11716
rect 16255 11713 16267 11747
rect 16387 11744 16396 11753
rect 16351 11716 16396 11744
rect 16209 11707 16267 11713
rect 16387 11707 16396 11716
rect 14826 11676 14832 11688
rect 14292 11648 14832 11676
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 15672 11676 15700 11704
rect 15948 11676 15976 11707
rect 16390 11704 16396 11707
rect 16448 11704 16454 11756
rect 17681 11747 17739 11753
rect 17681 11744 17693 11747
rect 16500 11716 17693 11744
rect 15672 11648 15976 11676
rect 11790 11608 11796 11620
rect 9364 11580 11796 11608
rect 9364 11568 9370 11580
rect 11790 11568 11796 11580
rect 11848 11568 11854 11620
rect 14185 11611 14243 11617
rect 14185 11577 14197 11611
rect 14231 11608 14243 11611
rect 14553 11611 14611 11617
rect 14553 11608 14565 11611
rect 14231 11580 14565 11608
rect 14231 11577 14243 11580
rect 14185 11571 14243 11577
rect 14553 11577 14565 11580
rect 14599 11577 14611 11611
rect 14553 11571 14611 11577
rect 14642 11568 14648 11620
rect 14700 11568 14706 11620
rect 14921 11611 14979 11617
rect 14921 11577 14933 11611
rect 14967 11608 14979 11611
rect 16500 11608 16528 11716
rect 17681 11713 17693 11716
rect 17727 11713 17739 11747
rect 17681 11707 17739 11713
rect 17770 11704 17776 11756
rect 17828 11744 17834 11756
rect 17865 11747 17923 11753
rect 17865 11744 17877 11747
rect 17828 11716 17877 11744
rect 17828 11704 17834 11716
rect 17865 11713 17877 11716
rect 17911 11713 17923 11747
rect 17972 11744 18000 11772
rect 18049 11747 18107 11753
rect 18049 11744 18061 11747
rect 17972 11716 18061 11744
rect 17865 11707 17923 11713
rect 18049 11713 18061 11716
rect 18095 11713 18107 11747
rect 18049 11707 18107 11713
rect 18230 11704 18236 11756
rect 18288 11704 18294 11756
rect 16850 11636 16856 11688
rect 16908 11636 16914 11688
rect 17402 11636 17408 11688
rect 17460 11676 17466 11688
rect 17957 11679 18015 11685
rect 17957 11676 17969 11679
rect 17460 11648 17969 11676
rect 17460 11636 17466 11648
rect 17957 11645 17969 11648
rect 18003 11645 18015 11679
rect 17957 11639 18015 11645
rect 14967 11580 16528 11608
rect 14967 11577 14979 11580
rect 14921 11571 14979 11577
rect 16942 11568 16948 11620
rect 17000 11608 17006 11620
rect 17497 11611 17555 11617
rect 17497 11608 17509 11611
rect 17000 11580 17509 11608
rect 17000 11568 17006 11580
rect 17497 11577 17509 11580
rect 17543 11577 17555 11611
rect 17497 11571 17555 11577
rect 6917 11543 6975 11549
rect 6917 11509 6929 11543
rect 6963 11540 6975 11543
rect 7282 11540 7288 11552
rect 6963 11512 7288 11540
rect 6963 11509 6975 11512
rect 6917 11503 6975 11509
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 7650 11500 7656 11552
rect 7708 11540 7714 11552
rect 8113 11543 8171 11549
rect 8113 11540 8125 11543
rect 7708 11512 8125 11540
rect 7708 11500 7714 11512
rect 8113 11509 8125 11512
rect 8159 11509 8171 11543
rect 8113 11503 8171 11509
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 16390 11540 16396 11552
rect 15436 11512 16396 11540
rect 15436 11500 15442 11512
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 17218 11500 17224 11552
rect 17276 11540 17282 11552
rect 17405 11543 17463 11549
rect 17405 11540 17417 11543
rect 17276 11512 17417 11540
rect 17276 11500 17282 11512
rect 17405 11509 17417 11512
rect 17451 11509 17463 11543
rect 17405 11503 17463 11509
rect 1104 11450 18860 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 18860 11450
rect 1104 11376 18860 11398
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 6825 11339 6883 11345
rect 6825 11336 6837 11339
rect 5868 11308 6837 11336
rect 5868 11296 5874 11308
rect 6825 11305 6837 11308
rect 6871 11305 6883 11339
rect 6825 11299 6883 11305
rect 13449 11339 13507 11345
rect 13449 11305 13461 11339
rect 13495 11336 13507 11339
rect 14642 11336 14648 11348
rect 13495 11308 14648 11336
rect 13495 11305 13507 11308
rect 13449 11299 13507 11305
rect 14642 11296 14648 11308
rect 14700 11296 14706 11348
rect 14826 11296 14832 11348
rect 14884 11296 14890 11348
rect 5994 11228 6000 11280
rect 6052 11268 6058 11280
rect 15654 11268 15660 11280
rect 6052 11240 7512 11268
rect 6052 11228 6058 11240
rect 7282 11160 7288 11212
rect 7340 11160 7346 11212
rect 7484 11209 7512 11240
rect 15028 11240 15660 11268
rect 7469 11203 7527 11209
rect 7469 11169 7481 11203
rect 7515 11200 7527 11203
rect 8754 11200 8760 11212
rect 7515 11172 8760 11200
rect 7515 11169 7527 11172
rect 7469 11163 7527 11169
rect 8754 11160 8760 11172
rect 8812 11160 8818 11212
rect 9217 11203 9275 11209
rect 9217 11169 9229 11203
rect 9263 11200 9275 11203
rect 9306 11200 9312 11212
rect 9263 11172 9312 11200
rect 9263 11169 9275 11172
rect 9217 11163 9275 11169
rect 9306 11160 9312 11172
rect 9364 11160 9370 11212
rect 9493 11203 9551 11209
rect 9493 11169 9505 11203
rect 9539 11200 9551 11203
rect 10502 11200 10508 11212
rect 9539 11172 10508 11200
rect 9539 11169 9551 11172
rect 9493 11163 9551 11169
rect 10502 11160 10508 11172
rect 10560 11160 10566 11212
rect 7190 11092 7196 11144
rect 7248 11092 7254 11144
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11132 9183 11135
rect 9674 11132 9680 11144
rect 9171 11104 9680 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 1578 11024 1584 11076
rect 1636 11064 1642 11076
rect 9140 11064 9168 11095
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11132 13783 11135
rect 14182 11132 14188 11144
rect 13771 11104 14188 11132
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 1636 11036 9168 11064
rect 1636 11024 1642 11036
rect 13446 11024 13452 11076
rect 13504 11024 13510 11076
rect 13633 11067 13691 11073
rect 13633 11033 13645 11067
rect 13679 11064 13691 11067
rect 13998 11064 14004 11076
rect 13679 11036 14004 11064
rect 13679 11033 13691 11036
rect 13633 11027 13691 11033
rect 13998 11024 14004 11036
rect 14056 11024 14062 11076
rect 14108 11064 14136 11104
rect 14182 11092 14188 11104
rect 14240 11092 14246 11144
rect 15028 11141 15056 11240
rect 15654 11228 15660 11240
rect 15712 11228 15718 11280
rect 16850 11228 16856 11280
rect 16908 11268 16914 11280
rect 16908 11240 18184 11268
rect 16908 11228 16914 11240
rect 18156 11212 18184 11240
rect 15746 11200 15752 11212
rect 15120 11172 15752 11200
rect 15120 11141 15148 11172
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 18046 11160 18052 11212
rect 18104 11160 18110 11212
rect 18138 11160 18144 11212
rect 18196 11160 18202 11212
rect 15013 11135 15071 11141
rect 15013 11101 15025 11135
rect 15059 11101 15071 11135
rect 15013 11095 15071 11101
rect 15105 11135 15163 11141
rect 15105 11101 15117 11135
rect 15151 11101 15163 11135
rect 15105 11095 15163 11101
rect 15286 11092 15292 11144
rect 15344 11092 15350 11144
rect 15378 11092 15384 11144
rect 15436 11092 15442 11144
rect 17862 11092 17868 11144
rect 17920 11132 17926 11144
rect 17957 11135 18015 11141
rect 17957 11132 17969 11135
rect 17920 11104 17969 11132
rect 17920 11092 17926 11104
rect 17957 11101 17969 11104
rect 18003 11101 18015 11135
rect 17957 11095 18015 11101
rect 15194 11064 15200 11076
rect 14108 11036 15200 11064
rect 15194 11024 15200 11036
rect 15252 11024 15258 11076
rect 8202 10956 8208 11008
rect 8260 10996 8266 11008
rect 12802 10996 12808 11008
rect 8260 10968 12808 10996
rect 8260 10956 8266 10968
rect 12802 10956 12808 10968
rect 12860 10956 12866 11008
rect 17586 10956 17592 11008
rect 17644 10956 17650 11008
rect 1104 10906 18860 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 18860 10906
rect 1104 10832 18860 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 3970 10792 3976 10804
rect 1627 10764 3976 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 10502 10752 10508 10804
rect 10560 10792 10566 10804
rect 13357 10795 13415 10801
rect 10560 10764 11836 10792
rect 10560 10752 10566 10764
rect 5902 10724 5908 10736
rect 5276 10696 5908 10724
rect 1302 10616 1308 10668
rect 1360 10656 1366 10668
rect 5276 10665 5304 10696
rect 5902 10684 5908 10696
rect 5960 10724 5966 10736
rect 9674 10724 9680 10736
rect 5960 10696 9680 10724
rect 5960 10684 5966 10696
rect 9674 10684 9680 10696
rect 9732 10684 9738 10736
rect 10686 10684 10692 10736
rect 10744 10724 10750 10736
rect 10965 10727 11023 10733
rect 10744 10696 10916 10724
rect 10744 10684 10750 10696
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 1360 10628 1409 10656
rect 1360 10616 1366 10628
rect 1397 10625 1409 10628
rect 1443 10656 1455 10659
rect 1673 10659 1731 10665
rect 1673 10656 1685 10659
rect 1443 10628 1685 10656
rect 1443 10625 1455 10628
rect 1397 10619 1455 10625
rect 1673 10625 1685 10628
rect 1719 10625 1731 10659
rect 1673 10619 1731 10625
rect 5261 10659 5319 10665
rect 5261 10625 5273 10659
rect 5307 10625 5319 10659
rect 5261 10619 5319 10625
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 5350 10548 5356 10600
rect 5408 10548 5414 10600
rect 8386 10480 8392 10532
rect 8444 10520 8450 10532
rect 8481 10523 8539 10529
rect 8481 10520 8493 10523
rect 8444 10492 8493 10520
rect 8444 10480 8450 10492
rect 8481 10489 8493 10492
rect 8527 10489 8539 10523
rect 8481 10483 8539 10489
rect 5629 10455 5687 10461
rect 5629 10421 5641 10455
rect 5675 10452 5687 10455
rect 6822 10452 6828 10464
rect 5675 10424 6828 10452
rect 5675 10421 5687 10424
rect 5629 10415 5687 10421
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 8680 10452 8708 10619
rect 10318 10616 10324 10668
rect 10376 10656 10382 10668
rect 10888 10665 10916 10696
rect 10965 10693 10977 10727
rect 11011 10724 11023 10727
rect 11808 10724 11836 10764
rect 13357 10761 13369 10795
rect 13403 10792 13415 10795
rect 13446 10792 13452 10804
rect 13403 10764 13452 10792
rect 13403 10761 13415 10764
rect 13357 10755 13415 10761
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 17221 10795 17279 10801
rect 17221 10761 17233 10795
rect 17267 10792 17279 10795
rect 17310 10792 17316 10804
rect 17267 10764 17316 10792
rect 17267 10761 17279 10764
rect 17221 10755 17279 10761
rect 17310 10752 17316 10764
rect 17368 10792 17374 10804
rect 17368 10764 18184 10792
rect 17368 10752 17374 10764
rect 18156 10733 18184 10764
rect 12529 10727 12587 10733
rect 12529 10724 12541 10727
rect 11011 10696 11744 10724
rect 11011 10693 11023 10696
rect 10965 10687 11023 10693
rect 11716 10665 11744 10696
rect 11808 10696 12541 10724
rect 10413 10659 10471 10665
rect 10413 10656 10425 10659
rect 10376 10628 10425 10656
rect 10376 10616 10382 10628
rect 10413 10625 10425 10628
rect 10459 10656 10471 10659
rect 10873 10659 10931 10665
rect 10459 10628 10824 10656
rect 10459 10625 10471 10628
rect 10413 10619 10471 10625
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10588 10563 10591
rect 10686 10588 10692 10600
rect 10551 10560 10692 10588
rect 10551 10557 10563 10560
rect 10505 10551 10563 10557
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 10796 10588 10824 10628
rect 10873 10625 10885 10659
rect 10919 10625 10931 10659
rect 10873 10619 10931 10625
rect 11057 10659 11115 10665
rect 11057 10625 11069 10659
rect 11103 10625 11115 10659
rect 11057 10619 11115 10625
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 11072 10588 11100 10619
rect 11808 10597 11836 10696
rect 12529 10693 12541 10696
rect 12575 10693 12587 10727
rect 12529 10687 12587 10693
rect 18141 10727 18199 10733
rect 18141 10693 18153 10727
rect 18187 10693 18199 10727
rect 18141 10687 18199 10693
rect 12802 10616 12808 10668
rect 12860 10616 12866 10668
rect 12986 10616 12992 10668
rect 13044 10656 13050 10668
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 13044 10628 13093 10656
rect 13044 10616 13050 10628
rect 13081 10625 13093 10628
rect 13127 10625 13139 10659
rect 13081 10619 13139 10625
rect 13170 10616 13176 10668
rect 13228 10616 13234 10668
rect 13998 10616 14004 10668
rect 14056 10656 14062 10668
rect 14185 10659 14243 10665
rect 14185 10656 14197 10659
rect 14056 10628 14197 10656
rect 14056 10616 14062 10628
rect 14185 10625 14197 10628
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 16669 10659 16727 10665
rect 16669 10625 16681 10659
rect 16715 10656 16727 10659
rect 16758 10656 16764 10668
rect 16715 10628 16764 10656
rect 16715 10625 16727 10628
rect 16669 10619 16727 10625
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 16942 10616 16948 10668
rect 17000 10616 17006 10668
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 10796 10560 11100 10588
rect 11793 10591 11851 10597
rect 11793 10557 11805 10591
rect 11839 10557 11851 10591
rect 11793 10551 11851 10557
rect 11974 10548 11980 10600
rect 12032 10588 12038 10600
rect 12161 10591 12219 10597
rect 12161 10588 12173 10591
rect 12032 10560 12173 10588
rect 12032 10548 12038 10560
rect 12161 10557 12173 10560
rect 12207 10557 12219 10591
rect 12820 10588 12848 10616
rect 15746 10588 15752 10600
rect 12820 10560 15752 10588
rect 12161 10551 12219 10557
rect 15746 10548 15752 10560
rect 15804 10548 15810 10600
rect 16850 10548 16856 10600
rect 16908 10588 16914 10600
rect 17052 10588 17080 10619
rect 16908 10560 17080 10588
rect 16908 10548 16914 10560
rect 10781 10523 10839 10529
rect 10781 10489 10793 10523
rect 10827 10520 10839 10523
rect 12069 10523 12127 10529
rect 10827 10492 11652 10520
rect 10827 10489 10839 10492
rect 10781 10483 10839 10489
rect 9030 10452 9036 10464
rect 8680 10424 9036 10452
rect 9030 10412 9036 10424
rect 9088 10452 9094 10464
rect 11146 10452 11152 10464
rect 9088 10424 11152 10452
rect 9088 10412 9094 10424
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 11624 10452 11652 10492
rect 12069 10489 12081 10523
rect 12115 10520 12127 10523
rect 13170 10520 13176 10532
rect 12115 10492 13176 10520
rect 12115 10489 12127 10492
rect 12069 10483 12127 10489
rect 13170 10480 13176 10492
rect 13228 10480 13234 10532
rect 16574 10480 16580 10532
rect 16632 10520 16638 10532
rect 16761 10523 16819 10529
rect 16761 10520 16773 10523
rect 16632 10492 16773 10520
rect 16632 10480 16638 10492
rect 16761 10489 16773 10492
rect 16807 10520 16819 10523
rect 17126 10520 17132 10532
rect 16807 10492 17132 10520
rect 16807 10489 16819 10492
rect 16761 10483 16819 10489
rect 17126 10480 17132 10492
rect 17184 10480 17190 10532
rect 12526 10452 12532 10464
rect 11624 10424 12532 10452
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 12713 10455 12771 10461
rect 12713 10421 12725 10455
rect 12759 10452 12771 10455
rect 12897 10455 12955 10461
rect 12897 10452 12909 10455
rect 12759 10424 12909 10452
rect 12759 10421 12771 10424
rect 12713 10415 12771 10421
rect 12897 10421 12909 10424
rect 12943 10421 12955 10455
rect 12897 10415 12955 10421
rect 14277 10455 14335 10461
rect 14277 10421 14289 10455
rect 14323 10452 14335 10455
rect 15286 10452 15292 10464
rect 14323 10424 15292 10452
rect 14323 10421 14335 10424
rect 14277 10415 14335 10421
rect 15286 10412 15292 10424
rect 15344 10412 15350 10464
rect 18049 10455 18107 10461
rect 18049 10421 18061 10455
rect 18095 10452 18107 10455
rect 18138 10452 18144 10464
rect 18095 10424 18144 10452
rect 18095 10421 18107 10424
rect 18049 10415 18107 10421
rect 18138 10412 18144 10424
rect 18196 10412 18202 10464
rect 1104 10362 18860 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 18860 10362
rect 1104 10288 18860 10310
rect 4614 10208 4620 10260
rect 4672 10208 4678 10260
rect 4801 10251 4859 10257
rect 4801 10217 4813 10251
rect 4847 10248 4859 10251
rect 5350 10248 5356 10260
rect 4847 10220 5356 10248
rect 4847 10217 4859 10220
rect 4801 10211 4859 10217
rect 5350 10208 5356 10220
rect 5408 10208 5414 10260
rect 7745 10251 7803 10257
rect 7745 10248 7757 10251
rect 6564 10220 7757 10248
rect 4632 10180 4660 10208
rect 4890 10180 4896 10192
rect 4632 10152 4896 10180
rect 4890 10140 4896 10152
rect 4948 10140 4954 10192
rect 5169 10183 5227 10189
rect 5169 10149 5181 10183
rect 5215 10149 5227 10183
rect 5169 10143 5227 10149
rect 4816 10084 5028 10112
rect 1302 10004 1308 10056
rect 1360 10044 1366 10056
rect 1397 10047 1455 10053
rect 1397 10044 1409 10047
rect 1360 10016 1409 10044
rect 1360 10004 1366 10016
rect 1397 10013 1409 10016
rect 1443 10044 1455 10047
rect 1673 10047 1731 10053
rect 1673 10044 1685 10047
rect 1443 10016 1685 10044
rect 1443 10013 1455 10016
rect 1397 10007 1455 10013
rect 1673 10013 1685 10016
rect 1719 10013 1731 10047
rect 1673 10007 1731 10013
rect 4433 9979 4491 9985
rect 4433 9945 4445 9979
rect 4479 9976 4491 9979
rect 4816 9976 4844 10084
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10013 4951 10047
rect 4893 10007 4951 10013
rect 4479 9948 4844 9976
rect 4479 9945 4491 9948
rect 4433 9939 4491 9945
rect 1578 9868 1584 9920
rect 1636 9868 1642 9920
rect 4614 9868 4620 9920
rect 4672 9917 4678 9920
rect 4672 9911 4691 9917
rect 4679 9908 4691 9911
rect 4908 9908 4936 10007
rect 5000 9976 5028 10084
rect 5184 10044 5212 10143
rect 5261 10047 5319 10053
rect 5261 10044 5273 10047
rect 5184 10016 5273 10044
rect 5261 10013 5273 10016
rect 5307 10013 5319 10047
rect 5368 10044 5396 10208
rect 5445 10047 5503 10053
rect 5445 10044 5457 10047
rect 5368 10016 5457 10044
rect 5261 10007 5319 10013
rect 5445 10013 5457 10016
rect 5491 10013 5503 10047
rect 5445 10007 5503 10013
rect 6178 10004 6184 10056
rect 6236 10044 6242 10056
rect 6457 10047 6515 10053
rect 6457 10044 6469 10047
rect 6236 10016 6469 10044
rect 6236 10004 6242 10016
rect 6457 10013 6469 10016
rect 6503 10044 6515 10047
rect 6564 10044 6592 10220
rect 7745 10217 7757 10220
rect 7791 10217 7803 10251
rect 7745 10211 7803 10217
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 9125 10251 9183 10257
rect 9125 10248 9137 10251
rect 8444 10220 9137 10248
rect 8444 10208 8450 10220
rect 9125 10217 9137 10220
rect 9171 10217 9183 10251
rect 9125 10211 9183 10217
rect 12986 10208 12992 10260
rect 13044 10208 13050 10260
rect 13170 10208 13176 10260
rect 13228 10248 13234 10260
rect 13228 10220 17080 10248
rect 13228 10208 13234 10220
rect 6822 10140 6828 10192
rect 6880 10180 6886 10192
rect 7009 10183 7067 10189
rect 7009 10180 7021 10183
rect 6880 10152 7021 10180
rect 6880 10140 6886 10152
rect 7009 10149 7021 10152
rect 7055 10149 7067 10183
rect 8205 10183 8263 10189
rect 8205 10180 8217 10183
rect 7009 10143 7067 10149
rect 7392 10152 8217 10180
rect 6914 10112 6920 10124
rect 6656 10084 6920 10112
rect 6656 10053 6684 10084
rect 6914 10072 6920 10084
rect 6972 10112 6978 10124
rect 7392 10121 7420 10152
rect 8205 10149 8217 10152
rect 8251 10149 8263 10183
rect 8941 10183 8999 10189
rect 8941 10180 8953 10183
rect 8205 10143 8263 10149
rect 8680 10152 8953 10180
rect 8680 10121 8708 10152
rect 8941 10149 8953 10152
rect 8987 10149 8999 10183
rect 8941 10143 8999 10149
rect 12526 10140 12532 10192
rect 12584 10180 12590 10192
rect 12897 10183 12955 10189
rect 12897 10180 12909 10183
rect 12584 10152 12909 10180
rect 12584 10140 12590 10152
rect 12897 10149 12909 10152
rect 12943 10180 12955 10183
rect 14829 10183 14887 10189
rect 12943 10152 14412 10180
rect 12943 10149 12955 10152
rect 12897 10143 12955 10149
rect 14384 10121 14412 10152
rect 14829 10149 14841 10183
rect 14875 10180 14887 10183
rect 15562 10180 15568 10192
rect 14875 10152 15568 10180
rect 14875 10149 14887 10152
rect 14829 10143 14887 10149
rect 15562 10140 15568 10152
rect 15620 10140 15626 10192
rect 15657 10183 15715 10189
rect 15657 10149 15669 10183
rect 15703 10180 15715 10183
rect 16666 10180 16672 10192
rect 15703 10152 16672 10180
rect 15703 10149 15715 10152
rect 15657 10143 15715 10149
rect 16666 10140 16672 10152
rect 16724 10140 16730 10192
rect 7377 10115 7435 10121
rect 7377 10112 7389 10115
rect 6972 10084 7389 10112
rect 6972 10072 6978 10084
rect 7377 10081 7389 10084
rect 7423 10081 7435 10115
rect 8665 10115 8723 10121
rect 8665 10112 8677 10115
rect 7377 10075 7435 10081
rect 7944 10084 8677 10112
rect 6503 10016 6592 10044
rect 6641 10047 6699 10053
rect 6503 10013 6515 10016
rect 6457 10007 6515 10013
rect 6641 10013 6653 10047
rect 6687 10013 6699 10047
rect 6641 10007 6699 10013
rect 6822 10004 6828 10056
rect 6880 10004 6886 10056
rect 7944 10053 7972 10084
rect 8665 10081 8677 10084
rect 8711 10081 8723 10115
rect 8665 10075 8723 10081
rect 14277 10115 14335 10121
rect 14277 10081 14289 10115
rect 14323 10081 14335 10115
rect 14277 10075 14335 10081
rect 14369 10115 14427 10121
rect 14369 10081 14381 10115
rect 14415 10081 14427 10115
rect 14369 10075 14427 10081
rect 15013 10115 15071 10121
rect 15013 10081 15025 10115
rect 15059 10081 15071 10115
rect 15013 10075 15071 10081
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10044 8631 10047
rect 10226 10044 10232 10056
rect 8619 10016 10232 10044
rect 8619 10013 8631 10016
rect 8573 10007 8631 10013
rect 10226 10004 10232 10016
rect 10284 10044 10290 10056
rect 14292 10044 14320 10075
rect 15028 10044 15056 10075
rect 15194 10072 15200 10124
rect 15252 10072 15258 10124
rect 16761 10115 16819 10121
rect 16761 10081 16773 10115
rect 16807 10112 16819 10115
rect 16942 10112 16948 10124
rect 16807 10084 16948 10112
rect 16807 10081 16819 10084
rect 16761 10075 16819 10081
rect 16942 10072 16948 10084
rect 17000 10072 17006 10124
rect 10284 10016 10456 10044
rect 14292 10016 15056 10044
rect 10284 10004 10290 10016
rect 5169 9979 5227 9985
rect 5169 9976 5181 9979
rect 5000 9948 5181 9976
rect 5169 9945 5181 9948
rect 5215 9945 5227 9979
rect 5169 9939 5227 9945
rect 5353 9979 5411 9985
rect 5353 9945 5365 9979
rect 5399 9976 5411 9979
rect 5534 9976 5540 9988
rect 5399 9948 5540 9976
rect 5399 9945 5411 9948
rect 5353 9939 5411 9945
rect 4679 9880 4936 9908
rect 4679 9877 4691 9880
rect 4672 9871 4691 9877
rect 4672 9868 4678 9871
rect 4982 9868 4988 9920
rect 5040 9868 5046 9920
rect 5184 9908 5212 9939
rect 5534 9936 5540 9948
rect 5592 9976 5598 9988
rect 6086 9976 6092 9988
rect 5592 9948 6092 9976
rect 5592 9936 5598 9948
rect 6086 9936 6092 9948
rect 6144 9976 6150 9988
rect 6549 9979 6607 9985
rect 6549 9976 6561 9979
rect 6144 9948 6561 9976
rect 6144 9936 6150 9948
rect 6549 9945 6561 9948
rect 6595 9945 6607 9979
rect 6549 9939 6607 9945
rect 8113 9979 8171 9985
rect 8113 9945 8125 9979
rect 8159 9976 8171 9979
rect 8294 9976 8300 9988
rect 8159 9948 8300 9976
rect 8159 9945 8171 9948
rect 8113 9939 8171 9945
rect 8294 9936 8300 9948
rect 8352 9936 8358 9988
rect 9309 9979 9367 9985
rect 9309 9945 9321 9979
rect 9355 9976 9367 9979
rect 9582 9976 9588 9988
rect 9355 9948 9588 9976
rect 9355 9945 9367 9948
rect 9309 9939 9367 9945
rect 9582 9936 9588 9948
rect 9640 9936 9646 9988
rect 5258 9908 5264 9920
rect 5184 9880 5264 9908
rect 5258 9868 5264 9880
rect 5316 9908 5322 9920
rect 5626 9908 5632 9920
rect 5316 9880 5632 9908
rect 5316 9868 5322 9880
rect 5626 9868 5632 9880
rect 5684 9868 5690 9920
rect 5994 9868 6000 9920
rect 6052 9868 6058 9920
rect 6270 9868 6276 9920
rect 6328 9868 6334 9920
rect 6917 9911 6975 9917
rect 6917 9877 6929 9911
rect 6963 9908 6975 9911
rect 7926 9908 7932 9920
rect 6963 9880 7932 9908
rect 6963 9877 6975 9880
rect 6917 9871 6975 9877
rect 7926 9868 7932 9880
rect 7984 9868 7990 9920
rect 8018 9868 8024 9920
rect 8076 9908 8082 9920
rect 9099 9911 9157 9917
rect 9099 9908 9111 9911
rect 8076 9880 9111 9908
rect 8076 9868 8082 9880
rect 9099 9877 9111 9880
rect 9145 9877 9157 9911
rect 10428 9908 10456 10016
rect 11974 9936 11980 9988
rect 12032 9976 12038 9988
rect 12529 9979 12587 9985
rect 12529 9976 12541 9979
rect 12032 9948 12541 9976
rect 12032 9936 12038 9948
rect 12529 9945 12541 9948
rect 12575 9976 12587 9979
rect 14461 9979 14519 9985
rect 14461 9976 14473 9979
rect 12575 9948 14473 9976
rect 12575 9945 12587 9948
rect 12529 9939 12587 9945
rect 14461 9945 14473 9948
rect 14507 9945 14519 9979
rect 15028 9976 15056 10016
rect 15286 10004 15292 10056
rect 15344 10004 15350 10056
rect 15746 10004 15752 10056
rect 15804 10004 15810 10056
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10013 15991 10047
rect 15933 10007 15991 10013
rect 16209 10047 16267 10053
rect 16209 10013 16221 10047
rect 16255 10044 16267 10047
rect 16301 10047 16359 10053
rect 16301 10044 16313 10047
rect 16255 10016 16313 10044
rect 16255 10013 16267 10016
rect 16209 10007 16267 10013
rect 16301 10013 16313 10016
rect 16347 10013 16359 10047
rect 16301 10007 16359 10013
rect 16485 10047 16543 10053
rect 16485 10013 16497 10047
rect 16531 10013 16543 10047
rect 16485 10007 16543 10013
rect 15948 9976 15976 10007
rect 16500 9976 16528 10007
rect 16574 10004 16580 10056
rect 16632 10044 16638 10056
rect 16669 10047 16727 10053
rect 16669 10044 16681 10047
rect 16632 10016 16681 10044
rect 16632 10004 16638 10016
rect 16669 10013 16681 10016
rect 16715 10013 16727 10047
rect 16669 10007 16727 10013
rect 16850 10004 16856 10056
rect 16908 10004 16914 10056
rect 17052 10053 17080 10220
rect 17405 10183 17463 10189
rect 17405 10149 17417 10183
rect 17451 10180 17463 10183
rect 17451 10152 17908 10180
rect 17451 10149 17463 10152
rect 17405 10143 17463 10149
rect 17681 10115 17739 10121
rect 17681 10112 17693 10115
rect 17512 10084 17693 10112
rect 17037 10047 17095 10053
rect 17037 10013 17049 10047
rect 17083 10013 17095 10047
rect 17037 10007 17095 10013
rect 17313 10047 17371 10053
rect 17313 10013 17325 10047
rect 17359 10044 17371 10047
rect 17402 10044 17408 10056
rect 17359 10016 17408 10044
rect 17359 10013 17371 10016
rect 17313 10007 17371 10013
rect 16758 9976 16764 9988
rect 15028 9948 16436 9976
rect 16500 9948 16764 9976
rect 14461 9939 14519 9945
rect 13538 9908 13544 9920
rect 10428 9880 13544 9908
rect 9099 9871 9157 9877
rect 13538 9868 13544 9880
rect 13596 9868 13602 9920
rect 16025 9911 16083 9917
rect 16025 9877 16037 9911
rect 16071 9908 16083 9911
rect 16206 9908 16212 9920
rect 16071 9880 16212 9908
rect 16071 9877 16083 9880
rect 16025 9871 16083 9877
rect 16206 9868 16212 9880
rect 16264 9868 16270 9920
rect 16408 9908 16436 9948
rect 16758 9936 16764 9948
rect 16816 9936 16822 9988
rect 16942 9936 16948 9988
rect 17000 9976 17006 9988
rect 17328 9976 17356 10007
rect 17402 10004 17408 10016
rect 17460 10004 17466 10056
rect 17000 9948 17356 9976
rect 17512 9976 17540 10084
rect 17681 10081 17693 10084
rect 17727 10081 17739 10115
rect 17681 10075 17739 10081
rect 17880 10053 17908 10152
rect 17865 10047 17923 10053
rect 17865 10013 17877 10047
rect 17911 10013 17923 10047
rect 17865 10007 17923 10013
rect 18138 9976 18144 9988
rect 17512 9948 18144 9976
rect 17000 9936 17006 9948
rect 17512 9908 17540 9948
rect 18138 9936 18144 9948
rect 18196 9936 18202 9988
rect 16408 9880 17540 9908
rect 17954 9868 17960 9920
rect 18012 9868 18018 9920
rect 18325 9911 18383 9917
rect 18325 9877 18337 9911
rect 18371 9908 18383 9911
rect 18506 9908 18512 9920
rect 18371 9880 18512 9908
rect 18371 9877 18383 9880
rect 18325 9871 18383 9877
rect 18506 9868 18512 9880
rect 18564 9868 18570 9920
rect 1104 9818 18860 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 18860 9818
rect 1104 9744 18860 9766
rect 2225 9707 2283 9713
rect 2225 9673 2237 9707
rect 2271 9704 2283 9707
rect 4617 9707 4675 9713
rect 2271 9676 3464 9704
rect 2271 9673 2283 9676
rect 2225 9667 2283 9673
rect 2682 9636 2688 9648
rect 2148 9608 2688 9636
rect 2148 9580 2176 9608
rect 2682 9596 2688 9608
rect 2740 9596 2746 9648
rect 3329 9639 3387 9645
rect 3329 9636 3341 9639
rect 2792 9608 3341 9636
rect 1578 9528 1584 9580
rect 1636 9528 1642 9580
rect 1670 9528 1676 9580
rect 1728 9528 1734 9580
rect 2130 9577 2136 9580
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9568 1915 9571
rect 1949 9571 2007 9577
rect 1949 9568 1961 9571
rect 1903 9540 1961 9568
rect 1903 9537 1915 9540
rect 1857 9531 1915 9537
rect 1949 9537 1961 9540
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 2093 9571 2136 9577
rect 2093 9537 2105 9571
rect 2093 9531 2136 9537
rect 2130 9528 2136 9531
rect 2188 9528 2194 9580
rect 2314 9528 2320 9580
rect 2372 9528 2378 9580
rect 2792 9577 2820 9608
rect 3329 9605 3341 9608
rect 3375 9605 3387 9639
rect 3329 9599 3387 9605
rect 3436 9580 3464 9676
rect 4617 9673 4629 9707
rect 4663 9704 4675 9707
rect 5534 9704 5540 9716
rect 4663 9676 5540 9704
rect 4663 9673 4675 9676
rect 4617 9667 4675 9673
rect 5534 9664 5540 9676
rect 5592 9664 5598 9716
rect 5626 9664 5632 9716
rect 5684 9704 5690 9716
rect 9214 9704 9220 9716
rect 5684 9676 9220 9704
rect 5684 9664 5690 9676
rect 9214 9664 9220 9676
rect 9272 9664 9278 9716
rect 16669 9707 16727 9713
rect 16669 9673 16681 9707
rect 16715 9704 16727 9707
rect 16850 9704 16856 9716
rect 16715 9676 16856 9704
rect 16715 9673 16727 9676
rect 16669 9667 16727 9673
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 4525 9639 4583 9645
rect 4525 9605 4537 9639
rect 4571 9636 4583 9639
rect 6089 9639 6147 9645
rect 6089 9636 6101 9639
rect 4571 9608 6101 9636
rect 4571 9605 4583 9608
rect 4525 9599 4583 9605
rect 6089 9605 6101 9608
rect 6135 9605 6147 9639
rect 6089 9599 6147 9605
rect 8113 9639 8171 9645
rect 8113 9605 8125 9639
rect 8159 9636 8171 9639
rect 8386 9636 8392 9648
rect 8159 9608 8392 9636
rect 8159 9605 8171 9608
rect 8113 9599 8171 9605
rect 8386 9596 8392 9608
rect 8444 9596 8450 9648
rect 16758 9596 16764 9648
rect 16816 9636 16822 9648
rect 17037 9639 17095 9645
rect 17037 9636 17049 9639
rect 16816 9608 17049 9636
rect 16816 9596 16822 9608
rect 17037 9605 17049 9608
rect 17083 9636 17095 9639
rect 17405 9639 17463 9645
rect 17083 9608 17356 9636
rect 17083 9605 17095 9608
rect 17037 9599 17095 9605
rect 2777 9571 2835 9577
rect 2777 9537 2789 9571
rect 2823 9537 2835 9571
rect 2777 9531 2835 9537
rect 2866 9528 2872 9580
rect 2924 9568 2930 9580
rect 3237 9571 3295 9577
rect 3237 9568 3249 9571
rect 2924 9540 3249 9568
rect 2924 9528 2930 9540
rect 3237 9537 3249 9540
rect 3283 9537 3295 9571
rect 3237 9531 3295 9537
rect 3418 9528 3424 9580
rect 3476 9528 3482 9580
rect 5994 9568 6000 9580
rect 5644 9540 6000 9568
rect 2332 9500 2360 9528
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 2332 9472 2697 9500
rect 2685 9469 2697 9472
rect 2731 9469 2743 9503
rect 2685 9463 2743 9469
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9500 4491 9503
rect 5442 9500 5448 9512
rect 4479 9472 5448 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 5442 9460 5448 9472
rect 5500 9500 5506 9512
rect 5644 9509 5672 9540
rect 5994 9528 6000 9540
rect 6052 9528 6058 9580
rect 6178 9528 6184 9580
rect 6236 9528 6242 9580
rect 6270 9528 6276 9580
rect 6328 9568 6334 9580
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 6328 9540 6561 9568
rect 6328 9528 6334 9540
rect 6549 9537 6561 9540
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 6638 9528 6644 9580
rect 6696 9528 6702 9580
rect 6914 9528 6920 9580
rect 6972 9528 6978 9580
rect 8018 9528 8024 9580
rect 8076 9528 8082 9580
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 9582 9568 9588 9580
rect 8343 9540 9588 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 9582 9528 9588 9540
rect 9640 9528 9646 9580
rect 11882 9528 11888 9580
rect 11940 9568 11946 9580
rect 12253 9571 12311 9577
rect 12253 9568 12265 9571
rect 11940 9540 12265 9568
rect 11940 9528 11946 9540
rect 12253 9537 12265 9540
rect 12299 9537 12311 9571
rect 12253 9531 12311 9537
rect 16850 9528 16856 9580
rect 16908 9528 16914 9580
rect 16945 9571 17003 9577
rect 16945 9537 16957 9571
rect 16991 9537 17003 9571
rect 16945 9531 17003 9537
rect 5629 9503 5687 9509
rect 5629 9500 5641 9503
rect 5500 9472 5641 9500
rect 5500 9460 5506 9472
rect 5629 9469 5641 9472
rect 5675 9469 5687 9503
rect 5629 9463 5687 9469
rect 5905 9503 5963 9509
rect 5905 9469 5917 9503
rect 5951 9500 5963 9503
rect 6365 9503 6423 9509
rect 6365 9500 6377 9503
rect 5951 9472 6377 9500
rect 5951 9469 5963 9472
rect 5905 9463 5963 9469
rect 6365 9469 6377 9472
rect 6411 9469 6423 9503
rect 6365 9463 6423 9469
rect 6822 9460 6828 9512
rect 6880 9460 6886 9512
rect 2501 9435 2559 9441
rect 2501 9401 2513 9435
rect 2547 9432 2559 9435
rect 2547 9404 8248 9432
rect 2547 9401 2559 9404
rect 2501 9395 2559 9401
rect 3053 9367 3111 9373
rect 3053 9333 3065 9367
rect 3099 9364 3111 9367
rect 4890 9364 4896 9376
rect 3099 9336 4896 9364
rect 3099 9333 3111 9336
rect 3053 9327 3111 9333
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 4985 9367 5043 9373
rect 4985 9333 4997 9367
rect 5031 9364 5043 9367
rect 5258 9364 5264 9376
rect 5031 9336 5264 9364
rect 5031 9333 5043 9336
rect 4985 9327 5043 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 8220 9364 8248 9404
rect 8294 9392 8300 9444
rect 8352 9392 8358 9444
rect 16960 9432 16988 9531
rect 17126 9528 17132 9580
rect 17184 9568 17190 9580
rect 17328 9577 17356 9608
rect 17405 9605 17417 9639
rect 17451 9636 17463 9639
rect 17451 9608 17816 9636
rect 17451 9605 17463 9608
rect 17405 9599 17463 9605
rect 17788 9577 17816 9608
rect 17221 9571 17279 9577
rect 17221 9568 17233 9571
rect 17184 9540 17233 9568
rect 17184 9528 17190 9540
rect 17221 9537 17233 9540
rect 17267 9537 17279 9571
rect 17221 9531 17279 9537
rect 17313 9571 17371 9577
rect 17313 9537 17325 9571
rect 17359 9537 17371 9571
rect 17313 9531 17371 9537
rect 17589 9571 17647 9577
rect 17589 9537 17601 9571
rect 17635 9537 17647 9571
rect 17589 9531 17647 9537
rect 17773 9571 17831 9577
rect 17773 9537 17785 9571
rect 17819 9537 17831 9571
rect 17773 9531 17831 9537
rect 17236 9500 17264 9531
rect 17604 9500 17632 9531
rect 17236 9472 17632 9500
rect 17954 9432 17960 9444
rect 16960 9404 17960 9432
rect 17954 9392 17960 9404
rect 18012 9392 18018 9444
rect 10778 9364 10784 9376
rect 8220 9336 10784 9364
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 12342 9324 12348 9376
rect 12400 9324 12406 9376
rect 17494 9324 17500 9376
rect 17552 9364 17558 9376
rect 17589 9367 17647 9373
rect 17589 9364 17601 9367
rect 17552 9336 17601 9364
rect 17552 9324 17558 9336
rect 17589 9333 17601 9336
rect 17635 9333 17647 9367
rect 17589 9327 17647 9333
rect 1104 9274 18860 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 18860 9274
rect 1104 9200 18860 9222
rect 1949 9163 2007 9169
rect 1949 9129 1961 9163
rect 1995 9160 2007 9163
rect 2314 9160 2320 9172
rect 1995 9132 2320 9160
rect 1995 9129 2007 9132
rect 1949 9123 2007 9129
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 4341 9163 4399 9169
rect 4341 9129 4353 9163
rect 4387 9160 4399 9163
rect 4614 9160 4620 9172
rect 4387 9132 4620 9160
rect 4387 9129 4399 9132
rect 4341 9123 4399 9129
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 4890 9120 4896 9172
rect 4948 9160 4954 9172
rect 4948 9132 9352 9160
rect 4948 9120 4954 9132
rect 3510 9052 3516 9104
rect 3568 9092 3574 9104
rect 3568 9064 4660 9092
rect 3568 9052 3574 9064
rect 1670 8984 1676 9036
rect 1728 8984 1734 9036
rect 4433 9027 4491 9033
rect 4433 8993 4445 9027
rect 4479 8993 4491 9027
rect 4632 9024 4660 9064
rect 4706 9052 4712 9104
rect 4764 9092 4770 9104
rect 9122 9092 9128 9104
rect 4764 9064 9128 9092
rect 4764 9052 4770 9064
rect 9122 9052 9128 9064
rect 9180 9052 9186 9104
rect 9324 9092 9352 9132
rect 9398 9120 9404 9172
rect 9456 9120 9462 9172
rect 9950 9160 9956 9172
rect 9508 9132 9956 9160
rect 9508 9092 9536 9132
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 10229 9163 10287 9169
rect 10229 9129 10241 9163
rect 10275 9160 10287 9163
rect 10275 9132 12296 9160
rect 10275 9129 10287 9132
rect 10229 9123 10287 9129
rect 9324 9064 9536 9092
rect 9585 9095 9643 9101
rect 9585 9061 9597 9095
rect 9631 9092 9643 9095
rect 12161 9095 12219 9101
rect 9631 9064 9812 9092
rect 9631 9061 9643 9064
rect 9585 9055 9643 9061
rect 4632 8996 6040 9024
rect 4433 8987 4491 8993
rect 1578 8916 1584 8968
rect 1636 8916 1642 8968
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8956 3479 8959
rect 3510 8956 3516 8968
rect 3467 8928 3516 8956
rect 3467 8925 3479 8928
rect 3421 8919 3479 8925
rect 3510 8916 3516 8928
rect 3568 8916 3574 8968
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8956 4031 8959
rect 4448 8956 4476 8987
rect 5350 8956 5356 8968
rect 4019 8928 5356 8956
rect 4019 8925 4031 8928
rect 3973 8919 4031 8925
rect 5350 8916 5356 8928
rect 5408 8916 5414 8968
rect 5813 8959 5871 8965
rect 5813 8925 5825 8959
rect 5859 8956 5871 8959
rect 5905 8959 5963 8965
rect 5905 8956 5917 8959
rect 5859 8928 5917 8956
rect 5859 8925 5871 8928
rect 5813 8919 5871 8925
rect 5905 8925 5917 8928
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 3605 8891 3663 8897
rect 3605 8857 3617 8891
rect 3651 8888 3663 8891
rect 3786 8888 3792 8900
rect 3651 8860 3792 8888
rect 3651 8857 3663 8860
rect 3605 8851 3663 8857
rect 3786 8848 3792 8860
rect 3844 8848 3850 8900
rect 4614 8848 4620 8900
rect 4672 8848 4678 8900
rect 4706 8848 4712 8900
rect 4764 8888 4770 8900
rect 5445 8891 5503 8897
rect 5445 8888 5457 8891
rect 4764 8860 5457 8888
rect 4764 8848 4770 8860
rect 5445 8857 5457 8860
rect 5491 8857 5503 8891
rect 5445 8851 5503 8857
rect 5626 8848 5632 8900
rect 5684 8848 5690 8900
rect 6012 8888 6040 8996
rect 6178 8984 6184 9036
rect 6236 8984 6242 9036
rect 6638 8984 6644 9036
rect 6696 8984 6702 9036
rect 8018 8984 8024 9036
rect 8076 8984 8082 9036
rect 9784 9033 9812 9064
rect 12161 9061 12173 9095
rect 12207 9061 12219 9095
rect 12268 9092 12296 9132
rect 12434 9120 12440 9172
rect 12492 9120 12498 9172
rect 13814 9160 13820 9172
rect 12544 9132 13820 9160
rect 12544 9092 12572 9132
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 12268 9064 12572 9092
rect 12621 9095 12679 9101
rect 12161 9055 12219 9061
rect 12621 9061 12633 9095
rect 12667 9061 12679 9095
rect 12621 9055 12679 9061
rect 9769 9027 9827 9033
rect 9769 8993 9781 9027
rect 9815 9024 9827 9027
rect 10042 9024 10048 9036
rect 9815 8996 10048 9024
rect 9815 8993 9827 8996
rect 9769 8987 9827 8993
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 6086 8916 6092 8968
rect 6144 8916 6150 8968
rect 6270 8916 6276 8968
rect 6328 8916 6334 8968
rect 6454 8916 6460 8968
rect 6512 8916 6518 8968
rect 8113 8959 8171 8965
rect 8113 8925 8125 8959
rect 8159 8956 8171 8959
rect 8294 8956 8300 8968
rect 8159 8928 8300 8956
rect 8159 8925 8171 8928
rect 8113 8919 8171 8925
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 9447 8925 9505 8931
rect 9447 8922 9459 8925
rect 8938 8888 8944 8900
rect 6012 8860 8944 8888
rect 8938 8848 8944 8860
rect 8996 8848 9002 8900
rect 9214 8848 9220 8900
rect 9272 8848 9278 8900
rect 9432 8891 9459 8922
rect 9493 8900 9505 8925
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 9861 8959 9919 8965
rect 9861 8956 9873 8959
rect 9732 8928 9873 8956
rect 9732 8916 9738 8928
rect 9861 8925 9873 8928
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 10134 8916 10140 8968
rect 10192 8956 10198 8968
rect 10781 8959 10839 8965
rect 10781 8956 10793 8959
rect 10192 8928 10793 8956
rect 10192 8916 10198 8928
rect 10781 8925 10793 8928
rect 10827 8956 10839 8959
rect 10870 8956 10876 8968
rect 10827 8928 10876 8956
rect 10827 8925 10839 8928
rect 10781 8919 10839 8925
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 11057 8959 11115 8965
rect 11057 8925 11069 8959
rect 11103 8956 11115 8959
rect 11882 8956 11888 8968
rect 11103 8928 11888 8956
rect 11103 8925 11115 8928
rect 11057 8919 11115 8925
rect 11882 8916 11888 8928
rect 11940 8916 11946 8968
rect 12176 8956 12204 9055
rect 12636 9024 12664 9055
rect 13449 9027 13507 9033
rect 13449 9024 13461 9027
rect 12636 8996 13461 9024
rect 13096 8965 13124 8996
rect 13449 8993 13461 8996
rect 13495 8993 13507 9027
rect 13449 8987 13507 8993
rect 12897 8959 12955 8965
rect 12897 8956 12909 8959
rect 12176 8928 12909 8956
rect 12897 8925 12909 8928
rect 12943 8925 12955 8959
rect 12897 8919 12955 8925
rect 13081 8959 13139 8965
rect 13081 8925 13093 8959
rect 13127 8925 13139 8959
rect 13081 8919 13139 8925
rect 13538 8916 13544 8968
rect 13596 8916 13602 8968
rect 9493 8891 9496 8900
rect 9432 8860 9496 8891
rect 9490 8848 9496 8860
rect 9548 8848 9554 8900
rect 10502 8848 10508 8900
rect 10560 8848 10566 8900
rect 10612 8860 11100 8888
rect 3878 8780 3884 8832
rect 3936 8820 3942 8832
rect 4065 8823 4123 8829
rect 4065 8820 4077 8823
rect 3936 8792 4077 8820
rect 3936 8780 3942 8792
rect 4065 8789 4077 8792
rect 4111 8789 4123 8823
rect 4065 8783 4123 8789
rect 4154 8780 4160 8832
rect 4212 8780 4218 8832
rect 5166 8780 5172 8832
rect 5224 8780 5230 8832
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 6362 8820 6368 8832
rect 5592 8792 6368 8820
rect 5592 8780 5598 8792
rect 6362 8780 6368 8792
rect 6420 8780 6426 8832
rect 7742 8780 7748 8832
rect 7800 8780 7806 8832
rect 9582 8780 9588 8832
rect 9640 8820 9646 8832
rect 10612 8820 10640 8860
rect 9640 8792 10640 8820
rect 9640 8780 9646 8792
rect 10686 8780 10692 8832
rect 10744 8780 10750 8832
rect 10778 8780 10784 8832
rect 10836 8820 10842 8832
rect 10873 8823 10931 8829
rect 10873 8820 10885 8823
rect 10836 8792 10885 8820
rect 10836 8780 10842 8792
rect 10873 8789 10885 8792
rect 10919 8789 10931 8823
rect 11072 8820 11100 8860
rect 11146 8848 11152 8900
rect 11204 8888 11210 8900
rect 11977 8891 12035 8897
rect 11977 8888 11989 8891
rect 11204 8860 11989 8888
rect 11204 8848 11210 8860
rect 11977 8857 11989 8860
rect 12023 8857 12035 8891
rect 11977 8851 12035 8857
rect 12161 8891 12219 8897
rect 12161 8857 12173 8891
rect 12207 8888 12219 8891
rect 12253 8891 12311 8897
rect 12253 8888 12265 8891
rect 12207 8860 12265 8888
rect 12207 8857 12219 8860
rect 12161 8851 12219 8857
rect 12253 8857 12265 8860
rect 12299 8857 12311 8891
rect 12253 8851 12311 8857
rect 13265 8891 13323 8897
rect 13265 8857 13277 8891
rect 13311 8888 13323 8891
rect 14182 8888 14188 8900
rect 13311 8860 14188 8888
rect 13311 8857 13323 8860
rect 13265 8851 13323 8857
rect 12176 8820 12204 8851
rect 14182 8848 14188 8860
rect 14240 8848 14246 8900
rect 11072 8792 12204 8820
rect 10873 8783 10931 8789
rect 12342 8780 12348 8832
rect 12400 8820 12406 8832
rect 12453 8823 12511 8829
rect 12453 8820 12465 8823
rect 12400 8792 12465 8820
rect 12400 8780 12406 8792
rect 12453 8789 12465 8792
rect 12499 8789 12511 8823
rect 12453 8783 12511 8789
rect 13906 8780 13912 8832
rect 13964 8780 13970 8832
rect 1104 8730 18860 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 18860 8730
rect 1104 8656 18860 8678
rect 1670 8576 1676 8628
rect 1728 8616 1734 8628
rect 2222 8616 2228 8628
rect 1728 8588 2228 8616
rect 1728 8576 1734 8588
rect 1872 8489 1900 8588
rect 2222 8576 2228 8588
rect 2280 8616 2286 8628
rect 5534 8616 5540 8628
rect 2280 8588 5540 8616
rect 2280 8576 2286 8588
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 6270 8576 6276 8628
rect 6328 8616 6334 8628
rect 6825 8619 6883 8625
rect 6825 8616 6837 8619
rect 6328 8588 6837 8616
rect 6328 8576 6334 8588
rect 6825 8585 6837 8588
rect 6871 8585 6883 8619
rect 6825 8579 6883 8585
rect 8294 8576 8300 8628
rect 8352 8616 8358 8628
rect 12434 8616 12440 8628
rect 8352 8588 12440 8616
rect 8352 8576 8358 8588
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 4985 8551 5043 8557
rect 4985 8517 4997 8551
rect 5031 8548 5043 8551
rect 5813 8551 5871 8557
rect 5813 8548 5825 8551
rect 5031 8520 5825 8548
rect 5031 8517 5043 8520
rect 4985 8511 5043 8517
rect 5813 8517 5825 8520
rect 5859 8517 5871 8551
rect 6178 8548 6184 8560
rect 5813 8511 5871 8517
rect 6012 8520 6184 8548
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8449 1915 8483
rect 1857 8443 1915 8449
rect 4706 8440 4712 8492
rect 4764 8480 4770 8492
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 4764 8452 4905 8480
rect 4764 8440 4770 8452
rect 4893 8449 4905 8452
rect 4939 8480 4951 8483
rect 5537 8483 5595 8489
rect 4939 8452 5488 8480
rect 4939 8449 4951 8452
rect 4893 8443 4951 8449
rect 1578 8372 1584 8424
rect 1636 8372 1642 8424
rect 2501 8415 2559 8421
rect 2501 8381 2513 8415
rect 2547 8412 2559 8415
rect 2774 8412 2780 8424
rect 2547 8384 2780 8412
rect 2547 8381 2559 8384
rect 2501 8375 2559 8381
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 5169 8415 5227 8421
rect 5169 8381 5181 8415
rect 5215 8381 5227 8415
rect 5460 8412 5488 8452
rect 5537 8449 5549 8483
rect 5583 8480 5595 8483
rect 5626 8480 5632 8492
rect 5583 8452 5632 8480
rect 5583 8449 5595 8452
rect 5537 8443 5595 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5905 8484 5963 8489
rect 6012 8484 6040 8520
rect 6178 8508 6184 8520
rect 6236 8548 6242 8560
rect 6457 8551 6515 8557
rect 6457 8548 6469 8551
rect 6236 8520 6469 8548
rect 6236 8508 6242 8520
rect 6457 8517 6469 8520
rect 6503 8548 6515 8551
rect 7742 8548 7748 8560
rect 6503 8520 7748 8548
rect 6503 8517 6515 8520
rect 6457 8511 6515 8517
rect 7742 8508 7748 8520
rect 7800 8508 7806 8560
rect 9214 8508 9220 8560
rect 9272 8548 9278 8560
rect 9769 8551 9827 8557
rect 9769 8548 9781 8551
rect 9272 8520 9781 8548
rect 9272 8508 9278 8520
rect 9769 8517 9781 8520
rect 9815 8517 9827 8551
rect 9769 8511 9827 8517
rect 10137 8551 10195 8557
rect 10137 8517 10149 8551
rect 10183 8548 10195 8551
rect 14090 8548 14096 8560
rect 10183 8520 14096 8548
rect 10183 8517 10195 8520
rect 10137 8511 10195 8517
rect 14090 8508 14096 8520
rect 14148 8508 14154 8560
rect 5905 8483 6040 8484
rect 5905 8449 5917 8483
rect 5951 8456 6040 8483
rect 6365 8483 6423 8489
rect 5951 8449 5963 8456
rect 5905 8443 5963 8449
rect 6365 8449 6377 8483
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8480 6699 8483
rect 6914 8480 6920 8492
rect 6687 8452 6920 8480
rect 6687 8449 6699 8452
rect 6641 8443 6699 8449
rect 6380 8412 6408 8443
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 7558 8440 7564 8492
rect 7616 8440 7622 8492
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8480 9643 8483
rect 9631 8452 9720 8480
rect 9631 8449 9643 8452
rect 9585 8443 9643 8449
rect 5460 8384 6408 8412
rect 5169 8375 5227 8381
rect 4525 8347 4583 8353
rect 4525 8313 4537 8347
rect 4571 8344 4583 8347
rect 4798 8344 4804 8356
rect 4571 8316 4804 8344
rect 4571 8313 4583 8316
rect 4525 8307 4583 8313
rect 4798 8304 4804 8316
rect 4856 8304 4862 8356
rect 5184 8344 5212 8375
rect 9398 8372 9404 8424
rect 9456 8412 9462 8424
rect 9692 8412 9720 8452
rect 10042 8440 10048 8492
rect 10100 8440 10106 8492
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8449 10287 8483
rect 10229 8443 10287 8449
rect 11977 8483 12035 8489
rect 11977 8449 11989 8483
rect 12023 8480 12035 8483
rect 12434 8480 12440 8492
rect 12023 8452 12440 8480
rect 12023 8449 12035 8452
rect 11977 8443 12035 8449
rect 10244 8412 10272 8443
rect 12434 8440 12440 8452
rect 12492 8480 12498 8492
rect 12621 8483 12679 8489
rect 12621 8480 12633 8483
rect 12492 8452 12633 8480
rect 12492 8440 12498 8452
rect 12621 8449 12633 8452
rect 12667 8449 12679 8483
rect 12621 8443 12679 8449
rect 9456 8384 9720 8412
rect 9456 8372 9462 8384
rect 5353 8347 5411 8353
rect 5353 8344 5365 8347
rect 5184 8316 5365 8344
rect 5353 8313 5365 8316
rect 5399 8344 5411 8347
rect 5442 8344 5448 8356
rect 5399 8316 5448 8344
rect 5399 8313 5411 8316
rect 5353 8307 5411 8313
rect 5442 8304 5448 8316
rect 5500 8304 5506 8356
rect 9416 8344 9444 8372
rect 5552 8316 9444 8344
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 5552 8276 5580 8316
rect 4948 8248 5580 8276
rect 4948 8236 4954 8248
rect 5626 8236 5632 8288
rect 5684 8276 5690 8288
rect 6089 8279 6147 8285
rect 6089 8276 6101 8279
rect 5684 8248 6101 8276
rect 5684 8236 5690 8248
rect 6089 8245 6101 8248
rect 6135 8276 6147 8279
rect 7190 8276 7196 8288
rect 6135 8248 7196 8276
rect 6135 8245 6147 8248
rect 6089 8239 6147 8245
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 7742 8236 7748 8288
rect 7800 8236 7806 8288
rect 9692 8276 9720 8384
rect 9784 8384 10272 8412
rect 12069 8415 12127 8421
rect 9784 8353 9812 8384
rect 12069 8381 12081 8415
rect 12115 8412 12127 8415
rect 12158 8412 12164 8424
rect 12115 8384 12164 8412
rect 12115 8381 12127 8384
rect 12069 8375 12127 8381
rect 12158 8372 12164 8384
rect 12216 8412 12222 8424
rect 12342 8412 12348 8424
rect 12216 8384 12348 8412
rect 12216 8372 12222 8384
rect 12342 8372 12348 8384
rect 12400 8412 12406 8424
rect 12529 8415 12587 8421
rect 12529 8412 12541 8415
rect 12400 8384 12541 8412
rect 12400 8372 12406 8384
rect 12529 8381 12541 8384
rect 12575 8381 12587 8415
rect 12529 8375 12587 8381
rect 9769 8347 9827 8353
rect 9769 8313 9781 8347
rect 9815 8313 9827 8347
rect 11698 8344 11704 8356
rect 9769 8307 9827 8313
rect 9876 8316 11704 8344
rect 9876 8276 9904 8316
rect 11698 8304 11704 8316
rect 11756 8304 11762 8356
rect 12986 8304 12992 8356
rect 13044 8304 13050 8356
rect 9692 8248 9904 8276
rect 12250 8236 12256 8288
rect 12308 8236 12314 8288
rect 1104 8186 18860 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 18860 8186
rect 1104 8112 18860 8134
rect 3528 8044 6868 8072
rect 1118 7896 1124 7948
rect 1176 7936 1182 7948
rect 3528 7945 3556 8044
rect 4706 7964 4712 8016
rect 4764 7964 4770 8016
rect 6840 8004 6868 8044
rect 6914 8032 6920 8084
rect 6972 8032 6978 8084
rect 8018 8032 8024 8084
rect 8076 8032 8082 8084
rect 7742 8004 7748 8016
rect 6840 7976 7420 8004
rect 1397 7939 1455 7945
rect 1397 7936 1409 7939
rect 1176 7908 1409 7936
rect 1176 7896 1182 7908
rect 1397 7905 1409 7908
rect 1443 7905 1455 7939
rect 1397 7899 1455 7905
rect 3513 7939 3571 7945
rect 3513 7905 3525 7939
rect 3559 7905 3571 7939
rect 3513 7899 3571 7905
rect 4433 7939 4491 7945
rect 4433 7905 4445 7939
rect 4479 7936 4491 7939
rect 7098 7936 7104 7948
rect 4479 7908 6500 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 2130 7868 2136 7880
rect 1719 7840 2136 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 2130 7828 2136 7840
rect 2188 7868 2194 7880
rect 2501 7871 2559 7877
rect 2501 7868 2513 7871
rect 2188 7840 2513 7868
rect 2188 7828 2194 7840
rect 2501 7837 2513 7840
rect 2547 7837 2559 7871
rect 3418 7868 3424 7880
rect 3174 7840 3424 7868
rect 2501 7831 2559 7837
rect 3418 7828 3424 7840
rect 3476 7828 3482 7880
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7868 4399 7871
rect 4890 7868 4896 7880
rect 4387 7840 4896 7868
rect 4387 7837 4399 7840
rect 4341 7831 4399 7837
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 6270 7828 6276 7880
rect 6328 7828 6334 7880
rect 6472 7877 6500 7908
rect 6656 7908 7104 7936
rect 6656 7877 6684 7908
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 6641 7871 6699 7877
rect 6641 7837 6653 7871
rect 6687 7837 6699 7871
rect 6641 7831 6699 7837
rect 6472 7732 6500 7831
rect 6564 7800 6592 7831
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 6788 7840 7021 7868
rect 6788 7828 6794 7840
rect 7009 7837 7021 7840
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 7282 7828 7288 7880
rect 7340 7828 7346 7880
rect 7392 7868 7420 7976
rect 7484 7976 7748 8004
rect 7484 7945 7512 7976
rect 7742 7964 7748 7976
rect 7800 8004 7806 8016
rect 8573 8007 8631 8013
rect 8573 8004 8585 8007
rect 7800 7976 8585 8004
rect 7800 7964 7806 7976
rect 8573 7973 8585 7976
rect 8619 8004 8631 8007
rect 10502 8004 10508 8016
rect 8619 7976 10508 8004
rect 8619 7973 8631 7976
rect 8573 7967 8631 7973
rect 10502 7964 10508 7976
rect 10560 7964 10566 8016
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7905 7527 7939
rect 9030 7936 9036 7948
rect 7469 7899 7527 7905
rect 7760 7908 9036 7936
rect 7760 7868 7788 7908
rect 9030 7896 9036 7908
rect 9088 7896 9094 7948
rect 7392 7840 7788 7868
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7868 7895 7871
rect 8297 7871 8355 7877
rect 8297 7868 8309 7871
rect 7883 7840 8309 7868
rect 7883 7837 7895 7840
rect 7837 7831 7895 7837
rect 8297 7837 8309 7840
rect 8343 7868 8355 7871
rect 10870 7868 10876 7880
rect 8343 7840 10876 7868
rect 8343 7837 8355 7840
rect 8297 7831 8355 7837
rect 10870 7828 10876 7840
rect 10928 7828 10934 7880
rect 11238 7828 11244 7880
rect 11296 7868 11302 7880
rect 18049 7871 18107 7877
rect 18049 7868 18061 7871
rect 11296 7840 18061 7868
rect 11296 7828 11302 7840
rect 18049 7837 18061 7840
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 6914 7800 6920 7812
rect 6564 7772 6920 7800
rect 6914 7760 6920 7772
rect 6972 7800 6978 7812
rect 7653 7803 7711 7809
rect 7653 7800 7665 7803
rect 6972 7772 7665 7800
rect 6972 7760 6978 7772
rect 7653 7769 7665 7772
rect 7699 7769 7711 7803
rect 7653 7763 7711 7769
rect 8110 7760 8116 7812
rect 8168 7800 8174 7812
rect 8389 7803 8447 7809
rect 8389 7800 8401 7803
rect 8168 7772 8401 7800
rect 8168 7760 8174 7772
rect 8389 7769 8401 7772
rect 8435 7769 8447 7803
rect 8389 7763 8447 7769
rect 18322 7760 18328 7812
rect 18380 7760 18386 7812
rect 6638 7732 6644 7744
rect 6472 7704 6644 7732
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 6730 7692 6736 7744
rect 6788 7732 6794 7744
rect 8205 7735 8263 7741
rect 8205 7732 8217 7735
rect 6788 7704 8217 7732
rect 6788 7692 6794 7704
rect 8205 7701 8217 7704
rect 8251 7701 8263 7735
rect 8205 7695 8263 7701
rect 1104 7642 18860 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 18860 7642
rect 1104 7568 18860 7590
rect 1578 7488 1584 7540
rect 1636 7488 1642 7540
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 4890 7528 4896 7540
rect 4212 7500 4896 7528
rect 4212 7488 4218 7500
rect 4890 7488 4896 7500
rect 4948 7488 4954 7540
rect 9122 7488 9128 7540
rect 9180 7488 9186 7540
rect 9490 7488 9496 7540
rect 9548 7488 9554 7540
rect 12069 7531 12127 7537
rect 12069 7497 12081 7531
rect 12115 7528 12127 7531
rect 12342 7528 12348 7540
rect 12115 7500 12348 7528
rect 12115 7497 12127 7500
rect 12069 7491 12127 7497
rect 12342 7488 12348 7500
rect 12400 7528 12406 7540
rect 12400 7500 12848 7528
rect 12400 7488 12406 7500
rect 1596 7460 1624 7488
rect 2133 7463 2191 7469
rect 1596 7432 2084 7460
rect 1302 7352 1308 7404
rect 1360 7392 1366 7404
rect 2056 7401 2084 7432
rect 2133 7429 2145 7463
rect 2179 7460 2191 7463
rect 3421 7463 3479 7469
rect 2179 7432 3188 7460
rect 2179 7429 2191 7432
rect 2133 7423 2191 7429
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 1360 7364 1409 7392
rect 1360 7352 1366 7364
rect 1397 7361 1409 7364
rect 1443 7392 1455 7395
rect 1857 7395 1915 7401
rect 1857 7392 1869 7395
rect 1443 7364 1869 7392
rect 1443 7361 1455 7364
rect 1397 7355 1455 7361
rect 1857 7361 1869 7364
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7361 2099 7395
rect 2041 7355 2099 7361
rect 2222 7352 2228 7404
rect 2280 7352 2286 7404
rect 2774 7352 2780 7404
rect 2832 7352 2838 7404
rect 3160 7401 3188 7432
rect 3421 7429 3433 7463
rect 3467 7460 3479 7463
rect 6178 7460 6184 7472
rect 3467 7432 6184 7460
rect 3467 7429 3479 7432
rect 3421 7423 3479 7429
rect 6178 7420 6184 7432
rect 6236 7460 6242 7472
rect 6730 7460 6736 7472
rect 6236 7432 6736 7460
rect 6236 7420 6242 7432
rect 6730 7420 6736 7432
rect 6788 7420 6794 7472
rect 7098 7460 7104 7472
rect 6840 7432 7104 7460
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7361 3203 7395
rect 3145 7355 3203 7361
rect 3878 7352 3884 7404
rect 3936 7392 3942 7404
rect 4617 7395 4675 7401
rect 4617 7392 4629 7395
rect 3936 7364 4629 7392
rect 3936 7352 3942 7364
rect 4617 7361 4629 7364
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 4890 7352 4896 7404
rect 4948 7352 4954 7404
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7392 5411 7395
rect 6270 7392 6276 7404
rect 5399 7364 6276 7392
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 1118 7284 1124 7336
rect 1176 7324 1182 7336
rect 1673 7327 1731 7333
rect 1673 7324 1685 7327
rect 1176 7296 1685 7324
rect 1176 7284 1182 7296
rect 1673 7293 1685 7296
rect 1719 7293 1731 7327
rect 1673 7287 1731 7293
rect 2501 7327 2559 7333
rect 2501 7293 2513 7327
rect 2547 7324 2559 7327
rect 2547 7296 2728 7324
rect 2547 7293 2559 7296
rect 2501 7287 2559 7293
rect 2700 7268 2728 7296
rect 3786 7284 3792 7336
rect 3844 7324 3850 7336
rect 4706 7324 4712 7336
rect 3844 7296 4712 7324
rect 3844 7284 3850 7296
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7293 4859 7327
rect 4801 7287 4859 7293
rect 5077 7327 5135 7333
rect 5077 7293 5089 7327
rect 5123 7324 5135 7327
rect 5368 7324 5396 7355
rect 6270 7352 6276 7364
rect 6328 7392 6334 7404
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 6328 7364 6561 7392
rect 6328 7352 6334 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6638 7352 6644 7404
rect 6696 7352 6702 7404
rect 6840 7401 6868 7432
rect 7098 7420 7104 7432
rect 7156 7460 7162 7472
rect 8018 7460 8024 7472
rect 7156 7432 8024 7460
rect 7156 7420 7162 7432
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7361 6883 7395
rect 6825 7355 6883 7361
rect 6914 7352 6920 7404
rect 6972 7392 6978 7404
rect 7208 7401 7236 7432
rect 8018 7420 8024 7432
rect 8076 7420 8082 7472
rect 8938 7420 8944 7472
rect 8996 7420 9002 7472
rect 10686 7460 10692 7472
rect 9048 7432 10692 7460
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 6972 7364 7021 7392
rect 6972 7352 6978 7364
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 7193 7395 7251 7401
rect 7193 7361 7205 7395
rect 7239 7361 7251 7395
rect 7193 7355 7251 7361
rect 7834 7352 7840 7404
rect 7892 7392 7898 7404
rect 9048 7392 9076 7432
rect 7892 7364 9076 7392
rect 7892 7352 7898 7364
rect 9214 7352 9220 7404
rect 9272 7352 9278 7404
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7392 9367 7395
rect 9582 7392 9588 7404
rect 9355 7364 9588 7392
rect 9355 7361 9367 7364
rect 9309 7355 9367 7361
rect 9582 7352 9588 7364
rect 9640 7352 9646 7404
rect 10336 7401 10364 7432
rect 10686 7420 10692 7432
rect 10744 7420 10750 7472
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 10502 7352 10508 7404
rect 10560 7352 10566 7404
rect 10870 7352 10876 7404
rect 10928 7352 10934 7404
rect 11698 7352 11704 7404
rect 11756 7352 11762 7404
rect 12820 7401 12848 7500
rect 12894 7488 12900 7540
rect 12952 7528 12958 7540
rect 13265 7531 13323 7537
rect 13265 7528 13277 7531
rect 12952 7500 13277 7528
rect 12952 7488 12958 7500
rect 13265 7497 13277 7500
rect 13311 7528 13323 7531
rect 15102 7528 15108 7540
rect 13311 7500 15108 7528
rect 13311 7497 13323 7500
rect 13265 7491 13323 7497
rect 15102 7488 15108 7500
rect 15160 7528 15166 7540
rect 18230 7528 18236 7540
rect 15160 7500 18236 7528
rect 15160 7488 15166 7500
rect 18230 7488 18236 7500
rect 18288 7488 18294 7540
rect 13906 7420 13912 7472
rect 13964 7460 13970 7472
rect 14001 7463 14059 7469
rect 14001 7460 14013 7463
rect 13964 7432 14013 7460
rect 13964 7420 13970 7432
rect 14001 7429 14013 7432
rect 14047 7460 14059 7463
rect 14642 7460 14648 7472
rect 14047 7432 14648 7460
rect 14047 7429 14059 7432
rect 14001 7423 14059 7429
rect 14642 7420 14648 7432
rect 14700 7420 14706 7472
rect 12805 7395 12863 7401
rect 12805 7361 12817 7395
rect 12851 7361 12863 7395
rect 12805 7355 12863 7361
rect 12989 7395 13047 7401
rect 12989 7361 13001 7395
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 13449 7395 13507 7401
rect 13449 7361 13461 7395
rect 13495 7361 13507 7395
rect 13449 7355 13507 7361
rect 5123 7296 5396 7324
rect 5537 7327 5595 7333
rect 5123 7293 5135 7296
rect 5077 7287 5135 7293
rect 5537 7293 5549 7327
rect 5583 7324 5595 7327
rect 6656 7324 6684 7352
rect 5583 7296 6684 7324
rect 5583 7293 5595 7296
rect 5537 7287 5595 7293
rect 2682 7216 2688 7268
rect 2740 7216 2746 7268
rect 4816 7256 4844 7287
rect 8938 7284 8944 7336
rect 8996 7324 9002 7336
rect 9766 7324 9772 7336
rect 8996 7296 9772 7324
rect 8996 7284 9002 7296
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 10229 7327 10287 7333
rect 10229 7293 10241 7327
rect 10275 7324 10287 7327
rect 10778 7324 10784 7336
rect 10275 7296 10784 7324
rect 10275 7293 10287 7296
rect 10229 7287 10287 7293
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 11790 7284 11796 7336
rect 11848 7284 11854 7336
rect 12250 7284 12256 7336
rect 12308 7324 12314 7336
rect 13004 7324 13032 7355
rect 12308 7296 13032 7324
rect 13464 7324 13492 7355
rect 13814 7352 13820 7404
rect 13872 7352 13878 7404
rect 14090 7352 14096 7404
rect 14148 7352 14154 7404
rect 14182 7352 14188 7404
rect 14240 7352 14246 7404
rect 13906 7324 13912 7336
rect 13464 7296 13912 7324
rect 12308 7284 12314 7296
rect 13906 7284 13912 7296
rect 13964 7284 13970 7336
rect 5350 7256 5356 7268
rect 4816 7228 5356 7256
rect 5350 7216 5356 7228
rect 5408 7216 5414 7268
rect 5626 7216 5632 7268
rect 5684 7256 5690 7268
rect 7009 7259 7067 7265
rect 7009 7256 7021 7259
rect 5684 7228 7021 7256
rect 5684 7216 5690 7228
rect 7009 7225 7021 7228
rect 7055 7225 7067 7259
rect 7009 7219 7067 7225
rect 7282 7216 7288 7268
rect 7340 7256 7346 7268
rect 7653 7259 7711 7265
rect 7653 7256 7665 7259
rect 7340 7228 7665 7256
rect 7340 7216 7346 7228
rect 7653 7225 7665 7228
rect 7699 7256 7711 7259
rect 8110 7256 8116 7268
rect 7699 7228 8116 7256
rect 7699 7225 7711 7228
rect 7653 7219 7711 7225
rect 8110 7216 8116 7228
rect 8168 7216 8174 7268
rect 10873 7259 10931 7265
rect 10873 7225 10885 7259
rect 10919 7256 10931 7259
rect 11330 7256 11336 7268
rect 10919 7228 11336 7256
rect 10919 7225 10931 7228
rect 10873 7219 10931 7225
rect 11330 7216 11336 7228
rect 11388 7216 11394 7268
rect 5166 7148 5172 7200
rect 5224 7148 5230 7200
rect 6365 7191 6423 7197
rect 6365 7157 6377 7191
rect 6411 7188 6423 7191
rect 6914 7188 6920 7200
rect 6411 7160 6920 7188
rect 6411 7157 6423 7160
rect 6365 7151 6423 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 9122 7148 9128 7200
rect 9180 7188 9186 7200
rect 9950 7188 9956 7200
rect 9180 7160 9956 7188
rect 9180 7148 9186 7160
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 13078 7148 13084 7200
rect 13136 7188 13142 7200
rect 13173 7191 13231 7197
rect 13173 7188 13185 7191
rect 13136 7160 13185 7188
rect 13136 7148 13142 7160
rect 13173 7157 13185 7160
rect 13219 7157 13231 7191
rect 13173 7151 13231 7157
rect 14274 7148 14280 7200
rect 14332 7188 14338 7200
rect 14369 7191 14427 7197
rect 14369 7188 14381 7191
rect 14332 7160 14381 7188
rect 14332 7148 14338 7160
rect 14369 7157 14381 7160
rect 14415 7157 14427 7191
rect 14369 7151 14427 7157
rect 1104 7098 18860 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 18860 7098
rect 1104 7024 18860 7046
rect 3878 6944 3884 6996
rect 3936 6984 3942 6996
rect 8205 6987 8263 6993
rect 3936 6956 8156 6984
rect 3936 6944 3942 6956
rect 4890 6876 4896 6928
rect 4948 6916 4954 6928
rect 8128 6916 8156 6956
rect 8205 6953 8217 6987
rect 8251 6984 8263 6987
rect 9122 6984 9128 6996
rect 8251 6956 9128 6984
rect 8251 6953 8263 6956
rect 8205 6947 8263 6953
rect 9122 6944 9128 6956
rect 9180 6944 9186 6996
rect 9582 6944 9588 6996
rect 9640 6984 9646 6996
rect 9640 6956 9996 6984
rect 9640 6944 9646 6956
rect 8754 6916 8760 6928
rect 4948 6888 5580 6916
rect 8128 6888 8760 6916
rect 4948 6876 4954 6888
rect 4801 6851 4859 6857
rect 4801 6817 4813 6851
rect 4847 6848 4859 6851
rect 5442 6848 5448 6860
rect 4847 6820 5448 6848
rect 4847 6817 4859 6820
rect 4801 6811 4859 6817
rect 5442 6808 5448 6820
rect 5500 6808 5506 6860
rect 2133 6783 2191 6789
rect 2133 6749 2145 6783
rect 2179 6780 2191 6783
rect 2866 6780 2872 6792
rect 2179 6752 2872 6780
rect 2179 6749 2191 6752
rect 2133 6743 2191 6749
rect 2866 6740 2872 6752
rect 2924 6780 2930 6792
rect 3418 6780 3424 6792
rect 2924 6752 3424 6780
rect 2924 6740 2930 6752
rect 3418 6740 3424 6752
rect 3476 6740 3482 6792
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6780 4583 6783
rect 5166 6780 5172 6792
rect 4571 6752 5172 6780
rect 4571 6749 4583 6752
rect 4525 6743 4583 6749
rect 5166 6740 5172 6752
rect 5224 6740 5230 6792
rect 5552 6780 5580 6888
rect 8754 6876 8760 6888
rect 8812 6916 8818 6928
rect 9214 6916 9220 6928
rect 8812 6888 9220 6916
rect 8812 6876 8818 6888
rect 9214 6876 9220 6888
rect 9272 6916 9278 6928
rect 9272 6888 9720 6916
rect 9272 6876 9278 6888
rect 8128 6820 9260 6848
rect 7742 6780 7748 6792
rect 5552 6752 7748 6780
rect 7742 6740 7748 6752
rect 7800 6780 7806 6792
rect 8018 6780 8024 6792
rect 7800 6752 8024 6780
rect 7800 6740 7806 6752
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 8128 6789 8156 6820
rect 9232 6792 9260 6820
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 1578 6672 1584 6724
rect 1636 6712 1642 6724
rect 1949 6715 2007 6721
rect 1949 6712 1961 6715
rect 1636 6684 1961 6712
rect 1636 6672 1642 6684
rect 1949 6681 1961 6684
rect 1995 6681 2007 6715
rect 1949 6675 2007 6681
rect 4617 6715 4675 6721
rect 4617 6681 4629 6715
rect 4663 6712 4675 6715
rect 5626 6712 5632 6724
rect 4663 6684 5632 6712
rect 4663 6681 4675 6684
rect 4617 6675 4675 6681
rect 5626 6672 5632 6684
rect 5684 6672 5690 6724
rect 8404 6712 8432 6743
rect 8754 6740 8760 6792
rect 8812 6740 8818 6792
rect 8941 6783 8999 6789
rect 8941 6749 8953 6783
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 8665 6715 8723 6721
rect 8665 6712 8677 6715
rect 8404 6684 8677 6712
rect 8665 6681 8677 6684
rect 8711 6712 8723 6715
rect 8956 6712 8984 6743
rect 9214 6740 9220 6792
rect 9272 6740 9278 6792
rect 9582 6740 9588 6792
rect 9640 6740 9646 6792
rect 9692 6780 9720 6888
rect 9766 6876 9772 6928
rect 9824 6916 9830 6928
rect 9824 6888 9904 6916
rect 9824 6876 9830 6888
rect 9876 6789 9904 6888
rect 9968 6848 9996 6956
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 14553 6987 14611 6993
rect 14553 6984 14565 6987
rect 13872 6956 14565 6984
rect 13872 6944 13878 6956
rect 14553 6953 14565 6956
rect 14599 6984 14611 6987
rect 14599 6956 14872 6984
rect 14599 6953 14611 6956
rect 14553 6947 14611 6953
rect 14844 6925 14872 6956
rect 14829 6919 14887 6925
rect 14829 6885 14841 6919
rect 14875 6885 14887 6919
rect 14829 6879 14887 6885
rect 10045 6851 10103 6857
rect 10045 6848 10057 6851
rect 9968 6820 10057 6848
rect 10045 6817 10057 6820
rect 10091 6817 10103 6851
rect 10045 6811 10103 6817
rect 10229 6851 10287 6857
rect 10229 6817 10241 6851
rect 10275 6848 10287 6851
rect 12342 6848 12348 6860
rect 10275 6820 11100 6848
rect 10275 6817 10287 6820
rect 10229 6811 10287 6817
rect 9769 6783 9827 6789
rect 9769 6780 9781 6783
rect 9692 6752 9781 6780
rect 9769 6749 9781 6752
rect 9815 6749 9827 6783
rect 9769 6743 9827 6749
rect 9861 6783 9919 6789
rect 9861 6749 9873 6783
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 9950 6740 9956 6792
rect 10008 6740 10014 6792
rect 11072 6789 11100 6820
rect 12268 6820 12348 6848
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6780 11115 6783
rect 11146 6780 11152 6792
rect 11103 6752 11152 6780
rect 11103 6749 11115 6752
rect 11057 6743 11115 6749
rect 11146 6740 11152 6752
rect 11204 6740 11210 6792
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6749 11299 6783
rect 11241 6743 11299 6749
rect 11256 6712 11284 6743
rect 11330 6740 11336 6792
rect 11388 6740 11394 6792
rect 11425 6783 11483 6789
rect 11425 6749 11437 6783
rect 11471 6780 11483 6783
rect 11606 6780 11612 6792
rect 11471 6752 11612 6780
rect 11471 6749 11483 6752
rect 11425 6743 11483 6749
rect 11606 6740 11612 6752
rect 11664 6780 11670 6792
rect 12158 6780 12164 6792
rect 11664 6752 12164 6780
rect 11664 6740 11670 6752
rect 12158 6740 12164 6752
rect 12216 6740 12222 6792
rect 12268 6789 12296 6820
rect 12342 6808 12348 6820
rect 12400 6848 12406 6860
rect 12400 6820 12848 6848
rect 12400 6808 12406 6820
rect 12253 6783 12311 6789
rect 12253 6749 12265 6783
rect 12299 6749 12311 6783
rect 12253 6743 12311 6749
rect 12529 6783 12587 6789
rect 12529 6749 12541 6783
rect 12575 6749 12587 6783
rect 12820 6780 12848 6820
rect 12894 6808 12900 6860
rect 12952 6808 12958 6860
rect 12986 6808 12992 6860
rect 13044 6848 13050 6860
rect 13081 6851 13139 6857
rect 13081 6848 13093 6851
rect 13044 6820 13093 6848
rect 13044 6808 13050 6820
rect 13081 6817 13093 6820
rect 13127 6817 13139 6851
rect 13081 6811 13139 6817
rect 13906 6808 13912 6860
rect 13964 6848 13970 6860
rect 14093 6851 14151 6857
rect 14093 6848 14105 6851
rect 13964 6820 14105 6848
rect 13964 6808 13970 6820
rect 14093 6817 14105 6820
rect 14139 6817 14151 6851
rect 14093 6811 14151 6817
rect 13173 6783 13231 6789
rect 13173 6780 13185 6783
rect 12820 6752 13185 6780
rect 12529 6743 12587 6749
rect 13173 6749 13185 6752
rect 13219 6749 13231 6783
rect 13173 6743 13231 6749
rect 8711 6684 8984 6712
rect 9416 6684 11284 6712
rect 11701 6715 11759 6721
rect 8711 6681 8723 6684
rect 8665 6675 8723 6681
rect 2317 6647 2375 6653
rect 2317 6613 2329 6647
rect 2363 6644 2375 6647
rect 2498 6644 2504 6656
rect 2363 6616 2504 6644
rect 2363 6613 2375 6616
rect 2317 6607 2375 6613
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 4157 6647 4215 6653
rect 4157 6613 4169 6647
rect 4203 6644 4215 6647
rect 4522 6644 4528 6656
rect 4203 6616 4528 6644
rect 4203 6613 4215 6616
rect 4157 6607 4215 6613
rect 4522 6604 4528 6616
rect 4580 6604 4586 6656
rect 6638 6604 6644 6656
rect 6696 6644 6702 6656
rect 9416 6653 9444 6684
rect 11072 6656 11100 6684
rect 11701 6681 11713 6715
rect 11747 6712 11759 6715
rect 12544 6712 12572 6743
rect 14274 6740 14280 6792
rect 14332 6740 14338 6792
rect 14366 6740 14372 6792
rect 14424 6740 14430 6792
rect 14642 6740 14648 6792
rect 14700 6780 14706 6792
rect 15197 6783 15255 6789
rect 15197 6780 15209 6783
rect 14700 6752 15209 6780
rect 14700 6740 14706 6752
rect 15197 6749 15209 6752
rect 15243 6749 15255 6783
rect 15197 6743 15255 6749
rect 11747 6684 12572 6712
rect 11747 6681 11759 6684
rect 11701 6675 11759 6681
rect 7929 6647 7987 6653
rect 7929 6644 7941 6647
rect 6696 6616 7941 6644
rect 6696 6604 6702 6616
rect 7929 6613 7941 6616
rect 7975 6613 7987 6647
rect 7929 6607 7987 6613
rect 9401 6647 9459 6653
rect 9401 6613 9413 6647
rect 9447 6613 9459 6647
rect 9401 6607 9459 6613
rect 11054 6604 11060 6656
rect 11112 6644 11118 6656
rect 11790 6644 11796 6656
rect 11112 6616 11796 6644
rect 11112 6604 11118 6616
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 12250 6604 12256 6656
rect 12308 6644 12314 6656
rect 12345 6647 12403 6653
rect 12345 6644 12357 6647
rect 12308 6616 12357 6644
rect 12308 6604 12314 6616
rect 12345 6613 12357 6616
rect 12391 6613 12403 6647
rect 12345 6607 12403 6613
rect 12713 6647 12771 6653
rect 12713 6613 12725 6647
rect 12759 6644 12771 6647
rect 13354 6644 13360 6656
rect 12759 6616 13360 6644
rect 12759 6613 12771 6616
rect 12713 6607 12771 6613
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 13541 6647 13599 6653
rect 13541 6613 13553 6647
rect 13587 6644 13599 6647
rect 13630 6644 13636 6656
rect 13587 6616 13636 6644
rect 13587 6613 13599 6616
rect 13541 6607 13599 6613
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 14642 6604 14648 6656
rect 14700 6644 14706 6656
rect 14737 6647 14795 6653
rect 14737 6644 14749 6647
rect 14700 6616 14749 6644
rect 14700 6604 14706 6616
rect 14737 6613 14749 6616
rect 14783 6613 14795 6647
rect 14737 6607 14795 6613
rect 1104 6554 18860 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 18860 6554
rect 1104 6480 18860 6502
rect 1578 6400 1584 6452
rect 1636 6400 1642 6452
rect 6365 6443 6423 6449
rect 6365 6409 6377 6443
rect 6411 6440 6423 6443
rect 6454 6440 6460 6452
rect 6411 6412 6460 6440
rect 6411 6409 6423 6412
rect 6365 6403 6423 6409
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 8849 6443 8907 6449
rect 8849 6409 8861 6443
rect 8895 6440 8907 6443
rect 9214 6440 9220 6452
rect 8895 6412 9220 6440
rect 8895 6409 8907 6412
rect 8849 6403 8907 6409
rect 8864 6372 8892 6403
rect 9214 6400 9220 6412
rect 9272 6400 9278 6452
rect 13725 6443 13783 6449
rect 13725 6409 13737 6443
rect 13771 6440 13783 6443
rect 14366 6440 14372 6452
rect 13771 6412 14372 6440
rect 13771 6409 13783 6412
rect 13725 6403 13783 6409
rect 14366 6400 14372 6412
rect 14424 6400 14430 6452
rect 14090 6372 14096 6384
rect 7944 6344 8892 6372
rect 11164 6344 11928 6372
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 1360 6276 1409 6304
rect 1360 6264 1366 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6304 2007 6307
rect 2682 6304 2688 6316
rect 1995 6276 2688 6304
rect 1995 6273 2007 6276
rect 1949 6267 2007 6273
rect 2682 6264 2688 6276
rect 2740 6304 2746 6316
rect 2777 6307 2835 6313
rect 2777 6304 2789 6307
rect 2740 6276 2789 6304
rect 2740 6264 2746 6276
rect 2777 6273 2789 6276
rect 2823 6273 2835 6307
rect 2777 6267 2835 6273
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 5592 6276 6561 6304
rect 5592 6264 5598 6276
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6822 6264 6828 6316
rect 6880 6264 6886 6316
rect 6914 6264 6920 6316
rect 6972 6304 6978 6316
rect 7944 6313 7972 6344
rect 11164 6316 11192 6344
rect 7009 6307 7067 6313
rect 7009 6304 7021 6307
rect 6972 6276 7021 6304
rect 6972 6264 6978 6276
rect 7009 6273 7021 6276
rect 7055 6273 7067 6307
rect 7009 6267 7067 6273
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 8018 6264 8024 6316
rect 8076 6304 8082 6316
rect 8205 6307 8263 6313
rect 8765 6308 8823 6313
rect 8205 6304 8217 6307
rect 8076 6276 8217 6304
rect 8076 6264 8082 6276
rect 8205 6273 8217 6276
rect 8251 6273 8263 6307
rect 8680 6307 8823 6308
rect 8680 6304 8777 6307
rect 8205 6267 8263 6273
rect 8312 6280 8777 6304
rect 8312 6276 8708 6280
rect 2041 6239 2099 6245
rect 2041 6205 2053 6239
rect 2087 6236 2099 6239
rect 2869 6239 2927 6245
rect 2869 6236 2881 6239
rect 2087 6208 2881 6236
rect 2087 6205 2099 6208
rect 2041 6199 2099 6205
rect 2746 6180 2774 6208
rect 2869 6205 2881 6208
rect 2915 6205 2927 6239
rect 2869 6199 2927 6205
rect 4706 6196 4712 6248
rect 4764 6236 4770 6248
rect 8312 6236 8340 6276
rect 8765 6273 8777 6280
rect 8811 6304 8823 6307
rect 8938 6304 8944 6316
rect 8811 6276 8944 6304
rect 8811 6273 8823 6276
rect 8765 6267 8823 6273
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 9033 6307 9091 6313
rect 9033 6273 9045 6307
rect 9079 6273 9091 6307
rect 9033 6267 9091 6273
rect 4764 6208 8340 6236
rect 4764 6196 4770 6208
rect 2746 6140 2780 6180
rect 2774 6128 2780 6140
rect 2832 6128 2838 6180
rect 3145 6171 3203 6177
rect 3145 6137 3157 6171
rect 3191 6168 3203 6171
rect 3694 6168 3700 6180
rect 3191 6140 3700 6168
rect 3191 6137 3203 6140
rect 3145 6131 3203 6137
rect 3694 6128 3700 6140
rect 3752 6128 3758 6180
rect 6638 6128 6644 6180
rect 6696 6128 6702 6180
rect 6730 6128 6736 6180
rect 6788 6128 6794 6180
rect 9048 6168 9076 6267
rect 11054 6264 11060 6316
rect 11112 6264 11118 6316
rect 11146 6264 11152 6316
rect 11204 6264 11210 6316
rect 11330 6264 11336 6316
rect 11388 6304 11394 6316
rect 11517 6307 11575 6313
rect 11517 6304 11529 6307
rect 11388 6276 11529 6304
rect 11388 6264 11394 6276
rect 11517 6273 11529 6276
rect 11563 6273 11575 6307
rect 11517 6267 11575 6273
rect 11532 6236 11560 6267
rect 11606 6264 11612 6316
rect 11664 6264 11670 6316
rect 11790 6264 11796 6316
rect 11848 6264 11854 6316
rect 11900 6313 11928 6344
rect 13188 6344 14096 6372
rect 11885 6307 11943 6313
rect 11885 6273 11897 6307
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 12161 6307 12219 6313
rect 12161 6273 12173 6307
rect 12207 6273 12219 6307
rect 12161 6267 12219 6273
rect 12176 6236 12204 6267
rect 12250 6264 12256 6316
rect 12308 6304 12314 6316
rect 12345 6307 12403 6313
rect 12345 6304 12357 6307
rect 12308 6276 12357 6304
rect 12308 6264 12314 6276
rect 12345 6273 12357 6276
rect 12391 6273 12403 6307
rect 12345 6267 12403 6273
rect 12989 6307 13047 6313
rect 12989 6273 13001 6307
rect 13035 6304 13047 6307
rect 13078 6304 13084 6316
rect 13035 6276 13084 6304
rect 13035 6273 13047 6276
rect 12989 6267 13047 6273
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 13188 6313 13216 6344
rect 14090 6332 14096 6344
rect 14148 6332 14154 6384
rect 13173 6307 13231 6313
rect 13173 6273 13185 6307
rect 13219 6273 13231 6307
rect 13173 6267 13231 6273
rect 13354 6264 13360 6316
rect 13412 6264 13418 6316
rect 13538 6264 13544 6316
rect 13596 6264 13602 6316
rect 11532 6208 12204 6236
rect 13265 6239 13323 6245
rect 13265 6205 13277 6239
rect 13311 6236 13323 6239
rect 14182 6236 14188 6248
rect 13311 6208 14188 6236
rect 13311 6205 13323 6208
rect 13265 6199 13323 6205
rect 14182 6196 14188 6208
rect 14240 6196 14246 6248
rect 9398 6168 9404 6180
rect 6840 6140 9404 6168
rect 2317 6103 2375 6109
rect 2317 6069 2329 6103
rect 2363 6100 2375 6103
rect 2590 6100 2596 6112
rect 2363 6072 2596 6100
rect 2363 6069 2375 6072
rect 2317 6063 2375 6069
rect 2590 6060 2596 6072
rect 2648 6060 2654 6112
rect 5350 6060 5356 6112
rect 5408 6100 5414 6112
rect 6840 6100 6868 6140
rect 9398 6128 9404 6140
rect 9456 6128 9462 6180
rect 11333 6171 11391 6177
rect 11333 6137 11345 6171
rect 11379 6168 11391 6171
rect 12434 6168 12440 6180
rect 11379 6140 12440 6168
rect 11379 6137 11391 6140
rect 11333 6131 11391 6137
rect 12434 6128 12440 6140
rect 12492 6128 12498 6180
rect 5408 6072 6868 6100
rect 5408 6060 5414 6072
rect 6914 6060 6920 6112
rect 6972 6100 6978 6112
rect 7653 6103 7711 6109
rect 7653 6100 7665 6103
rect 6972 6072 7665 6100
rect 6972 6060 6978 6072
rect 7653 6069 7665 6072
rect 7699 6069 7711 6103
rect 7653 6063 7711 6069
rect 8113 6103 8171 6109
rect 8113 6069 8125 6103
rect 8159 6100 8171 6103
rect 9125 6103 9183 6109
rect 9125 6100 9137 6103
rect 8159 6072 9137 6100
rect 8159 6069 8171 6072
rect 8113 6063 8171 6069
rect 9125 6069 9137 6072
rect 9171 6100 9183 6103
rect 9214 6100 9220 6112
rect 9171 6072 9220 6100
rect 9171 6069 9183 6072
rect 9125 6063 9183 6069
rect 9214 6060 9220 6072
rect 9272 6060 9278 6112
rect 12066 6060 12072 6112
rect 12124 6060 12130 6112
rect 12161 6103 12219 6109
rect 12161 6069 12173 6103
rect 12207 6100 12219 6103
rect 12526 6100 12532 6112
rect 12207 6072 12532 6100
rect 12207 6069 12219 6072
rect 12161 6063 12219 6069
rect 12526 6060 12532 6072
rect 12584 6060 12590 6112
rect 1104 6010 18860 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 18860 6010
rect 1104 5936 18860 5958
rect 1302 5856 1308 5908
rect 1360 5896 1366 5908
rect 1397 5899 1455 5905
rect 1397 5896 1409 5899
rect 1360 5868 1409 5896
rect 1360 5856 1366 5868
rect 1397 5865 1409 5868
rect 1443 5865 1455 5899
rect 1397 5859 1455 5865
rect 6365 5899 6423 5905
rect 6365 5865 6377 5899
rect 6411 5896 6423 5899
rect 6638 5896 6644 5908
rect 6411 5868 6644 5896
rect 6411 5865 6423 5868
rect 6365 5859 6423 5865
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 6822 5856 6828 5908
rect 6880 5896 6886 5908
rect 7009 5899 7067 5905
rect 7009 5896 7021 5899
rect 6880 5868 7021 5896
rect 6880 5856 6886 5868
rect 7009 5865 7021 5868
rect 7055 5865 7067 5899
rect 7009 5859 7067 5865
rect 7282 5856 7288 5908
rect 7340 5856 7346 5908
rect 9398 5856 9404 5908
rect 9456 5856 9462 5908
rect 13081 5899 13139 5905
rect 13081 5865 13093 5899
rect 13127 5896 13139 5899
rect 13538 5896 13544 5908
rect 13127 5868 13544 5896
rect 13127 5865 13139 5868
rect 13081 5859 13139 5865
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 5920 5800 6776 5828
rect 2866 5760 2872 5772
rect 2148 5732 2872 5760
rect 1578 5652 1584 5704
rect 1636 5692 1642 5704
rect 2148 5701 2176 5732
rect 2866 5720 2872 5732
rect 2924 5720 2930 5772
rect 5350 5760 5356 5772
rect 4632 5732 5356 5760
rect 1857 5695 1915 5701
rect 1857 5692 1869 5695
rect 1636 5664 1869 5692
rect 1636 5652 1642 5664
rect 1857 5661 1869 5664
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5661 2191 5695
rect 2133 5655 2191 5661
rect 2498 5652 2504 5704
rect 2556 5652 2562 5704
rect 2682 5652 2688 5704
rect 2740 5652 2746 5704
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5661 2835 5695
rect 2961 5695 3019 5701
rect 2961 5692 2973 5695
rect 2777 5655 2835 5661
rect 2884 5664 2973 5692
rect 2225 5627 2283 5633
rect 2225 5593 2237 5627
rect 2271 5624 2283 5627
rect 2516 5624 2544 5652
rect 2792 5624 2820 5655
rect 2271 5596 2452 5624
rect 2516 5596 2820 5624
rect 2271 5593 2283 5596
rect 2225 5587 2283 5593
rect 2314 5516 2320 5568
rect 2372 5516 2378 5568
rect 2424 5556 2452 5596
rect 2682 5556 2688 5568
rect 2424 5528 2688 5556
rect 2682 5516 2688 5528
rect 2740 5556 2746 5568
rect 2884 5556 2912 5664
rect 2961 5661 2973 5664
rect 3007 5661 3019 5695
rect 2961 5655 3019 5661
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 4632 5701 4660 5732
rect 5350 5720 5356 5732
rect 5408 5720 5414 5772
rect 5445 5763 5503 5769
rect 5445 5729 5457 5763
rect 5491 5760 5503 5763
rect 5920 5760 5948 5800
rect 6270 5760 6276 5772
rect 5491 5732 5948 5760
rect 5491 5729 5503 5732
rect 5445 5723 5503 5729
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 4212 5664 4537 5692
rect 4212 5652 4218 5664
rect 4525 5661 4537 5664
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 4706 5652 4712 5704
rect 4764 5692 4770 5704
rect 5920 5701 5948 5732
rect 6012 5732 6276 5760
rect 6012 5701 6040 5732
rect 6270 5720 6276 5732
rect 6328 5760 6334 5772
rect 6748 5760 6776 5800
rect 6914 5760 6920 5772
rect 6328 5732 6500 5760
rect 6328 5720 6334 5732
rect 4801 5695 4859 5701
rect 4801 5692 4813 5695
rect 4764 5664 4813 5692
rect 4764 5652 4770 5664
rect 4801 5661 4813 5664
rect 4847 5661 4859 5695
rect 4801 5655 4859 5661
rect 4985 5695 5043 5701
rect 4985 5661 4997 5695
rect 5031 5692 5043 5695
rect 5261 5695 5319 5701
rect 5261 5692 5273 5695
rect 5031 5664 5273 5692
rect 5031 5661 5043 5664
rect 4985 5655 5043 5661
rect 5261 5661 5273 5664
rect 5307 5692 5319 5695
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 5307 5664 5733 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 5721 5661 5733 5664
rect 5767 5661 5779 5695
rect 5721 5655 5779 5661
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5661 5963 5695
rect 5905 5655 5963 5661
rect 5997 5695 6055 5701
rect 5997 5661 6009 5695
rect 6043 5661 6055 5695
rect 5997 5655 6055 5661
rect 6089 5695 6147 5701
rect 6089 5661 6101 5695
rect 6135 5692 6147 5695
rect 6362 5692 6368 5704
rect 6135 5664 6368 5692
rect 6135 5661 6147 5664
rect 6089 5655 6147 5661
rect 5736 5624 5764 5655
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 6472 5701 6500 5732
rect 6748 5732 6920 5760
rect 6457 5695 6515 5701
rect 6457 5661 6469 5695
rect 6503 5661 6515 5695
rect 6457 5655 6515 5661
rect 6546 5652 6552 5704
rect 6604 5652 6610 5704
rect 6748 5701 6776 5732
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 9416 5760 9444 5856
rect 9677 5831 9735 5837
rect 9677 5797 9689 5831
rect 9723 5828 9735 5831
rect 11514 5828 11520 5840
rect 9723 5800 11520 5828
rect 9723 5797 9735 5800
rect 9677 5791 9735 5797
rect 11514 5788 11520 5800
rect 11572 5788 11578 5840
rect 9416 5732 10088 5760
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5661 6791 5695
rect 6733 5655 6791 5661
rect 6825 5695 6883 5701
rect 6825 5661 6837 5695
rect 6871 5661 6883 5695
rect 6825 5655 6883 5661
rect 6840 5624 6868 5655
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 7064 5664 7328 5692
rect 7064 5652 7070 5664
rect 7300 5633 7328 5664
rect 7558 5652 7564 5704
rect 7616 5692 7622 5704
rect 7653 5695 7711 5701
rect 7653 5692 7665 5695
rect 7616 5664 7665 5692
rect 7616 5652 7622 5664
rect 7653 5661 7665 5664
rect 7699 5661 7711 5695
rect 7653 5655 7711 5661
rect 9122 5652 9128 5704
rect 9180 5692 9186 5704
rect 9582 5692 9588 5704
rect 9180 5664 9588 5692
rect 9180 5652 9186 5664
rect 9582 5652 9588 5664
rect 9640 5692 9646 5704
rect 9953 5695 10011 5701
rect 9953 5692 9965 5695
rect 9640 5664 9965 5692
rect 9640 5652 9646 5664
rect 9953 5661 9965 5664
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 5736 5596 6868 5624
rect 7269 5627 7328 5633
rect 7269 5593 7281 5627
rect 7315 5596 7328 5627
rect 7469 5627 7527 5633
rect 7315 5593 7327 5596
rect 7269 5587 7327 5593
rect 7469 5593 7481 5627
rect 7515 5624 7527 5627
rect 7834 5624 7840 5636
rect 7515 5596 7840 5624
rect 7515 5593 7527 5596
rect 7469 5587 7527 5593
rect 7834 5584 7840 5596
rect 7892 5584 7898 5636
rect 8938 5584 8944 5636
rect 8996 5624 9002 5636
rect 9217 5627 9275 5633
rect 9217 5624 9229 5627
rect 8996 5596 9229 5624
rect 8996 5584 9002 5596
rect 9217 5593 9229 5596
rect 9263 5624 9275 5627
rect 9677 5627 9735 5633
rect 9677 5624 9689 5627
rect 9263 5596 9689 5624
rect 9263 5593 9275 5596
rect 9217 5587 9275 5593
rect 9677 5593 9689 5596
rect 9723 5593 9735 5627
rect 9677 5587 9735 5593
rect 9861 5627 9919 5633
rect 9861 5593 9873 5627
rect 9907 5624 9919 5627
rect 10060 5624 10088 5732
rect 12066 5652 12072 5704
rect 12124 5692 12130 5704
rect 12437 5695 12495 5701
rect 12437 5692 12449 5695
rect 12124 5664 12449 5692
rect 12124 5652 12130 5664
rect 12437 5661 12449 5664
rect 12483 5661 12495 5695
rect 12437 5655 12495 5661
rect 12618 5652 12624 5704
rect 12676 5652 12682 5704
rect 12710 5652 12716 5704
rect 12768 5652 12774 5704
rect 12802 5652 12808 5704
rect 12860 5652 12866 5704
rect 12897 5695 12955 5701
rect 12897 5661 12909 5695
rect 12943 5661 12955 5695
rect 12897 5655 12955 5661
rect 9907 5596 10088 5624
rect 9907 5593 9919 5596
rect 9861 5587 9919 5593
rect 12158 5584 12164 5636
rect 12216 5624 12222 5636
rect 12912 5624 12940 5655
rect 12216 5596 12940 5624
rect 12216 5584 12222 5596
rect 2740 5528 2912 5556
rect 2740 5516 2746 5528
rect 2958 5516 2964 5568
rect 3016 5516 3022 5568
rect 5077 5559 5135 5565
rect 5077 5525 5089 5559
rect 5123 5556 5135 5559
rect 5350 5556 5356 5568
rect 5123 5528 5356 5556
rect 5123 5525 5135 5528
rect 5077 5519 5135 5525
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 5442 5516 5448 5568
rect 5500 5556 5506 5568
rect 5626 5556 5632 5568
rect 5500 5528 5632 5556
rect 5500 5516 5506 5528
rect 5626 5516 5632 5528
rect 5684 5516 5690 5568
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 7101 5559 7159 5565
rect 7101 5556 7113 5559
rect 6604 5528 7113 5556
rect 6604 5516 6610 5528
rect 7101 5525 7113 5528
rect 7147 5525 7159 5559
rect 7101 5519 7159 5525
rect 9122 5516 9128 5568
rect 9180 5556 9186 5568
rect 9417 5559 9475 5565
rect 9417 5556 9429 5559
rect 9180 5528 9429 5556
rect 9180 5516 9186 5528
rect 9417 5525 9429 5528
rect 9463 5525 9475 5559
rect 9417 5519 9475 5525
rect 9585 5559 9643 5565
rect 9585 5525 9597 5559
rect 9631 5556 9643 5559
rect 9766 5556 9772 5568
rect 9631 5528 9772 5556
rect 9631 5525 9643 5528
rect 9585 5519 9643 5525
rect 9766 5516 9772 5528
rect 9824 5516 9830 5568
rect 1104 5466 18860 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 18860 5466
rect 1104 5392 18860 5414
rect 4985 5355 5043 5361
rect 4985 5321 4997 5355
rect 5031 5352 5043 5355
rect 5534 5352 5540 5364
rect 5031 5324 5540 5352
rect 5031 5321 5043 5324
rect 4985 5315 5043 5321
rect 5534 5312 5540 5324
rect 5592 5312 5598 5364
rect 6089 5355 6147 5361
rect 6089 5321 6101 5355
rect 6135 5352 6147 5355
rect 6730 5352 6736 5364
rect 6135 5324 6736 5352
rect 6135 5321 6147 5324
rect 6089 5315 6147 5321
rect 6730 5312 6736 5324
rect 6788 5312 6794 5364
rect 10965 5355 11023 5361
rect 10965 5321 10977 5355
rect 11011 5352 11023 5355
rect 11011 5324 11468 5352
rect 11011 5321 11023 5324
rect 10965 5315 11023 5321
rect 2958 5244 2964 5296
rect 3016 5284 3022 5296
rect 3605 5287 3663 5293
rect 3605 5284 3617 5287
rect 3016 5256 3617 5284
rect 3016 5244 3022 5256
rect 3605 5253 3617 5256
rect 3651 5253 3663 5287
rect 3605 5247 3663 5253
rect 3694 5244 3700 5296
rect 3752 5284 3758 5296
rect 3752 5256 4476 5284
rect 3752 5244 3758 5256
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 1360 5188 1409 5216
rect 1360 5176 1366 5188
rect 1397 5185 1409 5188
rect 1443 5216 1455 5219
rect 1673 5219 1731 5225
rect 1673 5216 1685 5219
rect 1443 5188 1685 5216
rect 1443 5185 1455 5188
rect 1397 5179 1455 5185
rect 1673 5185 1685 5188
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 3418 5176 3424 5228
rect 3476 5176 3482 5228
rect 4448 5225 4476 5256
rect 5442 5244 5448 5296
rect 5500 5284 5506 5296
rect 6457 5287 6515 5293
rect 6457 5284 6469 5287
rect 5500 5256 6469 5284
rect 5500 5244 5506 5256
rect 6457 5253 6469 5256
rect 6503 5253 6515 5287
rect 6457 5247 6515 5253
rect 6914 5244 6920 5296
rect 6972 5284 6978 5296
rect 7834 5284 7840 5296
rect 6972 5256 7840 5284
rect 6972 5244 6978 5256
rect 7834 5244 7840 5256
rect 7892 5284 7898 5296
rect 10594 5284 10600 5296
rect 7892 5256 10600 5284
rect 7892 5244 7898 5256
rect 10594 5244 10600 5256
rect 10652 5244 10658 5296
rect 3789 5219 3847 5225
rect 3789 5185 3801 5219
rect 3835 5216 3847 5219
rect 4249 5219 4307 5225
rect 4249 5216 4261 5219
rect 3835 5188 3924 5216
rect 3835 5185 3847 5188
rect 3789 5179 3847 5185
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 2130 5012 2136 5024
rect 1627 4984 2136 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 3896 5012 3924 5188
rect 3988 5188 4261 5216
rect 3988 5089 4016 5188
rect 4249 5185 4261 5188
rect 4295 5185 4307 5219
rect 4249 5179 4307 5185
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5185 4491 5219
rect 4433 5179 4491 5185
rect 4525 5219 4583 5225
rect 4525 5185 4537 5219
rect 4571 5216 4583 5219
rect 4706 5216 4712 5228
rect 4571 5188 4712 5216
rect 4571 5185 4583 5188
rect 4525 5179 4583 5185
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 4801 5219 4859 5225
rect 4801 5185 4813 5219
rect 4847 5216 4859 5219
rect 4890 5216 4896 5228
rect 4847 5188 4896 5216
rect 4847 5185 4859 5188
rect 4801 5179 4859 5185
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 5902 5216 5908 5228
rect 5644 5188 5908 5216
rect 4617 5151 4675 5157
rect 4617 5117 4629 5151
rect 4663 5148 4675 5151
rect 5644 5148 5672 5188
rect 5902 5176 5908 5188
rect 5960 5176 5966 5228
rect 6270 5176 6276 5228
rect 6328 5216 6334 5228
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 6328 5188 6377 5216
rect 6328 5176 6334 5188
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 4663 5120 5672 5148
rect 5721 5151 5779 5157
rect 4663 5117 4675 5120
rect 4617 5111 4675 5117
rect 5721 5117 5733 5151
rect 5767 5117 5779 5151
rect 6380 5148 6408 5179
rect 6546 5176 6552 5228
rect 6604 5176 6610 5228
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 6788 5188 6837 5216
rect 6788 5176 6794 5188
rect 6825 5185 6837 5188
rect 6871 5216 6883 5219
rect 7006 5216 7012 5228
rect 6871 5188 7012 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 7101 5219 7159 5225
rect 7101 5185 7113 5219
rect 7147 5216 7159 5219
rect 7282 5216 7288 5228
rect 7147 5188 7288 5216
rect 7147 5185 7159 5188
rect 7101 5179 7159 5185
rect 7282 5176 7288 5188
rect 7340 5216 7346 5228
rect 7929 5219 7987 5225
rect 7340 5188 7788 5216
rect 7340 5176 7346 5188
rect 6380 5120 7144 5148
rect 5721 5111 5779 5117
rect 3973 5083 4031 5089
rect 3973 5049 3985 5083
rect 4019 5049 4031 5083
rect 3973 5043 4031 5049
rect 4706 5012 4712 5024
rect 3896 4984 4712 5012
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 4890 4972 4896 5024
rect 4948 5012 4954 5024
rect 5534 5012 5540 5024
rect 4948 4984 5540 5012
rect 4948 4972 4954 4984
rect 5534 4972 5540 4984
rect 5592 5012 5598 5024
rect 5736 5012 5764 5111
rect 7116 5089 7144 5120
rect 7101 5083 7159 5089
rect 7101 5049 7113 5083
rect 7147 5049 7159 5083
rect 7760 5080 7788 5188
rect 7929 5185 7941 5219
rect 7975 5216 7987 5219
rect 9214 5216 9220 5228
rect 7975 5188 9220 5216
rect 7975 5185 7987 5188
rect 7929 5179 7987 5185
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 10505 5219 10563 5225
rect 10505 5185 10517 5219
rect 10551 5216 10563 5219
rect 10686 5216 10692 5228
rect 10551 5188 10692 5216
rect 10551 5185 10563 5188
rect 10505 5179 10563 5185
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 10781 5219 10839 5225
rect 11060 5222 11118 5225
rect 10781 5185 10793 5219
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 10888 5219 11118 5222
rect 10888 5194 11072 5219
rect 7834 5108 7840 5160
rect 7892 5108 7898 5160
rect 9122 5108 9128 5160
rect 9180 5108 9186 5160
rect 10796 5148 10824 5179
rect 10888 5160 10916 5194
rect 11060 5185 11072 5194
rect 11106 5185 11118 5219
rect 11060 5179 11118 5185
rect 11241 5219 11299 5225
rect 11241 5185 11253 5219
rect 11287 5185 11299 5219
rect 11241 5179 11299 5185
rect 9232 5120 10824 5148
rect 9232 5080 9260 5120
rect 7760 5052 9260 5080
rect 9585 5083 9643 5089
rect 7101 5043 7159 5049
rect 9585 5049 9597 5083
rect 9631 5080 9643 5083
rect 10686 5080 10692 5092
rect 9631 5052 10692 5080
rect 9631 5049 9643 5052
rect 9585 5043 9643 5049
rect 10686 5040 10692 5052
rect 10744 5040 10750 5092
rect 10796 5080 10824 5120
rect 10870 5108 10876 5160
rect 10928 5108 10934 5160
rect 11256 5080 11284 5179
rect 11330 5176 11336 5228
rect 11388 5176 11394 5228
rect 11440 5148 11468 5324
rect 12618 5312 12624 5364
rect 12676 5352 12682 5364
rect 13449 5355 13507 5361
rect 13449 5352 13461 5355
rect 12676 5324 13461 5352
rect 12676 5312 12682 5324
rect 13449 5321 13461 5324
rect 13495 5321 13507 5355
rect 13449 5315 13507 5321
rect 12529 5287 12587 5293
rect 12529 5253 12541 5287
rect 12575 5284 12587 5287
rect 12802 5284 12808 5296
rect 12575 5256 12808 5284
rect 12575 5253 12587 5256
rect 12529 5247 12587 5253
rect 12802 5244 12808 5256
rect 12860 5244 12866 5296
rect 12894 5244 12900 5296
rect 12952 5284 12958 5296
rect 12952 5256 13400 5284
rect 12952 5244 12958 5256
rect 11514 5176 11520 5228
rect 11572 5216 11578 5228
rect 12342 5216 12348 5228
rect 11572 5188 12348 5216
rect 11572 5176 11578 5188
rect 12342 5176 12348 5188
rect 12400 5216 12406 5228
rect 12621 5219 12679 5225
rect 12400 5214 12480 5216
rect 12621 5214 12633 5219
rect 12400 5188 12633 5214
rect 12400 5176 12406 5188
rect 12452 5186 12633 5188
rect 12621 5185 12633 5186
rect 12667 5185 12679 5219
rect 12621 5179 12679 5185
rect 12989 5219 13047 5225
rect 12989 5185 13001 5219
rect 13035 5185 13047 5219
rect 12989 5179 13047 5185
rect 12802 5148 12808 5160
rect 11440 5120 12808 5148
rect 12802 5108 12808 5120
rect 12860 5148 12866 5160
rect 13004 5148 13032 5179
rect 13078 5176 13084 5228
rect 13136 5176 13142 5228
rect 13372 5225 13400 5256
rect 13357 5219 13415 5225
rect 13357 5185 13369 5219
rect 13403 5185 13415 5219
rect 13357 5179 13415 5185
rect 14001 5219 14059 5225
rect 14001 5185 14013 5219
rect 14047 5216 14059 5219
rect 14182 5216 14188 5228
rect 14047 5188 14188 5216
rect 14047 5185 14059 5188
rect 14001 5179 14059 5185
rect 14182 5176 14188 5188
rect 14240 5176 14246 5228
rect 13449 5151 13507 5157
rect 13449 5148 13461 5151
rect 12860 5120 13461 5148
rect 12860 5108 12866 5120
rect 13449 5117 13461 5120
rect 13495 5117 13507 5151
rect 13449 5111 13507 5117
rect 10796 5052 11284 5080
rect 11333 5083 11391 5089
rect 11333 5049 11345 5083
rect 11379 5080 11391 5083
rect 12526 5080 12532 5092
rect 11379 5052 12532 5080
rect 11379 5049 11391 5052
rect 11333 5043 11391 5049
rect 12526 5040 12532 5052
rect 12584 5080 12590 5092
rect 12894 5080 12900 5092
rect 12584 5052 12900 5080
rect 12584 5040 12590 5052
rect 12894 5040 12900 5052
rect 12952 5040 12958 5092
rect 7653 5015 7711 5021
rect 7653 5012 7665 5015
rect 5592 4984 7665 5012
rect 5592 4972 5598 4984
rect 7653 4981 7665 4984
rect 7699 4981 7711 5015
rect 7653 4975 7711 4981
rect 9766 4972 9772 5024
rect 9824 5012 9830 5024
rect 12713 5015 12771 5021
rect 12713 5012 12725 5015
rect 9824 4984 12725 5012
rect 9824 4972 9830 4984
rect 12713 4981 12725 4984
rect 12759 5012 12771 5015
rect 13078 5012 13084 5024
rect 12759 4984 13084 5012
rect 12759 4981 12771 4984
rect 12713 4975 12771 4981
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 13170 4972 13176 5024
rect 13228 4972 13234 5024
rect 14093 5015 14151 5021
rect 14093 4981 14105 5015
rect 14139 5012 14151 5015
rect 14550 5012 14556 5024
rect 14139 4984 14556 5012
rect 14139 4981 14151 4984
rect 14093 4975 14151 4981
rect 14550 4972 14556 4984
rect 14608 4972 14614 5024
rect 1104 4922 18860 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 18860 4922
rect 1104 4848 18860 4870
rect 5902 4768 5908 4820
rect 5960 4808 5966 4820
rect 6549 4811 6607 4817
rect 6549 4808 6561 4811
rect 5960 4780 6561 4808
rect 5960 4768 5966 4780
rect 6549 4777 6561 4780
rect 6595 4777 6607 4811
rect 6549 4771 6607 4777
rect 8665 4811 8723 4817
rect 8665 4777 8677 4811
rect 8711 4808 8723 4811
rect 9122 4808 9128 4820
rect 8711 4780 9128 4808
rect 8711 4777 8723 4780
rect 8665 4771 8723 4777
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 3068 4712 8524 4740
rect 3068 4681 3096 4712
rect 8496 4684 8524 4712
rect 10778 4700 10784 4752
rect 10836 4740 10842 4752
rect 10836 4712 10916 4740
rect 10836 4700 10842 4712
rect 3053 4675 3111 4681
rect 3053 4641 3065 4675
rect 3099 4641 3111 4675
rect 3053 4635 3111 4641
rect 6178 4632 6184 4684
rect 6236 4672 6242 4684
rect 6730 4672 6736 4684
rect 6236 4644 6736 4672
rect 6236 4632 6242 4644
rect 6730 4632 6736 4644
rect 6788 4632 6794 4684
rect 8478 4632 8484 4684
rect 8536 4632 8542 4684
rect 10888 4681 10916 4712
rect 10873 4675 10931 4681
rect 10873 4641 10885 4675
rect 10919 4641 10931 4675
rect 10873 4635 10931 4641
rect 11330 4632 11336 4684
rect 11388 4632 11394 4684
rect 12526 4632 12532 4684
rect 12584 4632 12590 4684
rect 14550 4632 14556 4684
rect 14608 4632 14614 4684
rect 14734 4632 14740 4684
rect 14792 4672 14798 4684
rect 14921 4675 14979 4681
rect 14921 4672 14933 4675
rect 14792 4644 14933 4672
rect 14792 4632 14798 4644
rect 14921 4641 14933 4644
rect 14967 4641 14979 4675
rect 14921 4635 14979 4641
rect 2136 4616 2188 4622
rect 2038 4564 2044 4616
rect 2096 4564 2102 4616
rect 6825 4607 6883 4613
rect 6825 4573 6837 4607
rect 6871 4604 6883 4607
rect 6914 4604 6920 4616
rect 6871 4576 6920 4604
rect 6871 4573 6883 4576
rect 6825 4567 6883 4573
rect 6914 4564 6920 4576
rect 6972 4564 6978 4616
rect 8205 4607 8263 4613
rect 8205 4604 8217 4607
rect 7024 4576 8217 4604
rect 2136 4558 2188 4564
rect 2498 4496 2504 4548
rect 2556 4536 2562 4548
rect 7024 4536 7052 4576
rect 8205 4573 8217 4576
rect 8251 4573 8263 4607
rect 8205 4567 8263 4573
rect 8297 4607 8355 4613
rect 8297 4573 8309 4607
rect 8343 4573 8355 4607
rect 8297 4567 8355 4573
rect 8312 4536 8340 4567
rect 8386 4564 8392 4616
rect 8444 4564 8450 4616
rect 10778 4564 10784 4616
rect 10836 4564 10842 4616
rect 11241 4607 11299 4613
rect 11241 4573 11253 4607
rect 11287 4604 11299 4607
rect 11348 4604 11376 4632
rect 11287 4576 11376 4604
rect 12713 4607 12771 4613
rect 11287 4573 11299 4576
rect 11241 4567 11299 4573
rect 12713 4573 12725 4607
rect 12759 4604 12771 4607
rect 12802 4604 12808 4616
rect 12759 4576 12808 4604
rect 12759 4573 12771 4576
rect 12713 4567 12771 4573
rect 12802 4564 12808 4576
rect 12860 4564 12866 4616
rect 12989 4607 13047 4613
rect 12989 4573 13001 4607
rect 13035 4604 13047 4607
rect 13078 4604 13084 4616
rect 13035 4576 13084 4604
rect 13035 4573 13047 4576
rect 12989 4567 13047 4573
rect 13078 4564 13084 4576
rect 13136 4564 13142 4616
rect 13170 4564 13176 4616
rect 13228 4564 13234 4616
rect 14090 4564 14096 4616
rect 14148 4604 14154 4616
rect 14461 4607 14519 4613
rect 14461 4604 14473 4607
rect 14148 4576 14473 4604
rect 14148 4564 14154 4576
rect 14461 4573 14473 4576
rect 14507 4573 14519 4607
rect 14461 4567 14519 4573
rect 15102 4564 15108 4616
rect 15160 4564 15166 4616
rect 2556 4508 7052 4536
rect 7944 4508 8340 4536
rect 10796 4536 10824 4564
rect 11333 4539 11391 4545
rect 11333 4536 11345 4539
rect 10796 4508 11345 4536
rect 2556 4496 2562 4508
rect 6454 4428 6460 4480
rect 6512 4468 6518 4480
rect 7944 4477 7972 4508
rect 11333 4505 11345 4508
rect 11379 4505 11391 4539
rect 11333 4499 11391 4505
rect 12342 4496 12348 4548
rect 12400 4536 12406 4548
rect 13188 4536 13216 4564
rect 12400 4508 13216 4536
rect 12400 4496 12406 4508
rect 7929 4471 7987 4477
rect 7929 4468 7941 4471
rect 6512 4440 7941 4468
rect 6512 4428 6518 4440
rect 7929 4437 7941 4440
rect 7975 4437 7987 4471
rect 7929 4431 7987 4437
rect 11146 4428 11152 4480
rect 11204 4428 11210 4480
rect 12894 4428 12900 4480
rect 12952 4428 12958 4480
rect 13078 4428 13084 4480
rect 13136 4428 13142 4480
rect 14090 4428 14096 4480
rect 14148 4428 14154 4480
rect 1104 4378 18860 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 18860 4378
rect 1104 4304 18860 4326
rect 1762 4224 1768 4276
rect 1820 4264 1826 4276
rect 1820 4236 2452 4264
rect 1820 4224 1826 4236
rect 2130 4156 2136 4208
rect 2188 4156 2194 4208
rect 2424 4196 2452 4236
rect 2498 4224 2504 4276
rect 2556 4224 2562 4276
rect 5350 4224 5356 4276
rect 5408 4224 5414 4276
rect 3881 4199 3939 4205
rect 3881 4196 3893 4199
rect 2424 4168 3893 4196
rect 3881 4165 3893 4168
rect 3927 4165 3939 4199
rect 3881 4159 3939 4165
rect 1946 4088 1952 4140
rect 2004 4088 2010 4140
rect 2148 4128 2176 4156
rect 2317 4131 2375 4137
rect 2317 4128 2329 4131
rect 2148 4100 2329 4128
rect 2317 4097 2329 4100
rect 2363 4097 2375 4131
rect 2317 4091 2375 4097
rect 1394 4020 1400 4072
rect 1452 4060 1458 4072
rect 1673 4063 1731 4069
rect 1673 4060 1685 4063
rect 1452 4032 1685 4060
rect 1452 4020 1458 4032
rect 1673 4029 1685 4032
rect 1719 4029 1731 4063
rect 1673 4023 1731 4029
rect 2038 4020 2044 4072
rect 2096 4060 2102 4072
rect 2133 4063 2191 4069
rect 2133 4060 2145 4063
rect 2096 4032 2145 4060
rect 2096 4020 2102 4032
rect 2133 4029 2145 4032
rect 2179 4029 2191 4063
rect 3896 4060 3924 4159
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 4617 4131 4675 4137
rect 4617 4128 4629 4131
rect 4028 4100 4629 4128
rect 4028 4088 4034 4100
rect 4617 4097 4629 4100
rect 4663 4128 4675 4131
rect 5074 4128 5080 4140
rect 4663 4100 5080 4128
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 5442 4088 5448 4140
rect 5500 4088 5506 4140
rect 6454 4128 6460 4140
rect 5552 4100 6460 4128
rect 4893 4063 4951 4069
rect 4893 4060 4905 4063
rect 3896 4032 4905 4060
rect 2133 4023 2191 4029
rect 4893 4029 4905 4032
rect 4939 4060 4951 4063
rect 5552 4060 5580 4100
rect 6454 4088 6460 4100
rect 6512 4088 6518 4140
rect 6733 4131 6791 4137
rect 6733 4097 6745 4131
rect 6779 4128 6791 4131
rect 10778 4128 10784 4140
rect 6779 4100 10784 4128
rect 6779 4097 6791 4100
rect 6733 4091 6791 4097
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 11146 4088 11152 4140
rect 11204 4128 11210 4140
rect 12342 4128 12348 4140
rect 11204 4100 12348 4128
rect 11204 4088 11210 4100
rect 12342 4088 12348 4100
rect 12400 4128 12406 4140
rect 12437 4131 12495 4137
rect 12437 4128 12449 4131
rect 12400 4100 12449 4128
rect 12400 4088 12406 4100
rect 12437 4097 12449 4100
rect 12483 4097 12495 4131
rect 12437 4091 12495 4097
rect 12618 4088 12624 4140
rect 12676 4088 12682 4140
rect 4939 4032 5580 4060
rect 4939 4029 4951 4032
rect 4893 4023 4951 4029
rect 5626 4020 5632 4072
rect 5684 4020 5690 4072
rect 6822 4020 6828 4072
rect 6880 4020 6886 4072
rect 12621 3995 12679 4001
rect 12621 3961 12633 3995
rect 12667 3992 12679 3995
rect 12710 3992 12716 4004
rect 12667 3964 12716 3992
rect 12667 3961 12679 3964
rect 12621 3955 12679 3961
rect 12710 3952 12716 3964
rect 12768 3952 12774 4004
rect 4982 3884 4988 3936
rect 5040 3884 5046 3936
rect 5350 3884 5356 3936
rect 5408 3924 5414 3936
rect 6457 3927 6515 3933
rect 6457 3924 6469 3927
rect 5408 3896 6469 3924
rect 5408 3884 5414 3896
rect 6457 3893 6469 3896
rect 6503 3893 6515 3927
rect 6457 3887 6515 3893
rect 7190 3884 7196 3936
rect 7248 3924 7254 3936
rect 17957 3927 18015 3933
rect 17957 3924 17969 3927
rect 7248 3896 17969 3924
rect 7248 3884 7254 3896
rect 17957 3893 17969 3896
rect 18003 3924 18015 3927
rect 18046 3924 18052 3936
rect 18003 3896 18052 3924
rect 18003 3893 18015 3896
rect 17957 3887 18015 3893
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 1104 3834 18860 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 18860 3834
rect 1104 3760 18860 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 1627 3692 4108 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 3326 3612 3332 3664
rect 3384 3652 3390 3664
rect 3970 3652 3976 3664
rect 3384 3624 3976 3652
rect 3384 3612 3390 3624
rect 3970 3612 3976 3624
rect 4028 3612 4034 3664
rect 4080 3652 4108 3692
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 4341 3723 4399 3729
rect 4341 3720 4353 3723
rect 4304 3692 4353 3720
rect 4304 3680 4310 3692
rect 4341 3689 4353 3692
rect 4387 3689 4399 3723
rect 4341 3683 4399 3689
rect 4430 3680 4436 3732
rect 4488 3720 4494 3732
rect 4706 3720 4712 3732
rect 4488 3692 4712 3720
rect 4488 3680 4494 3692
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 9030 3680 9036 3732
rect 9088 3720 9094 3732
rect 9766 3720 9772 3732
rect 9088 3692 9772 3720
rect 9088 3680 9094 3692
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 12158 3680 12164 3732
rect 12216 3680 12222 3732
rect 8757 3655 8815 3661
rect 4080 3624 5028 3652
rect 1578 3544 1584 3596
rect 1636 3584 1642 3596
rect 1949 3587 2007 3593
rect 1949 3584 1961 3587
rect 1636 3556 1961 3584
rect 1636 3544 1642 3556
rect 1949 3553 1961 3556
rect 1995 3553 2007 3587
rect 1949 3547 2007 3553
rect 2409 3587 2467 3593
rect 2409 3553 2421 3587
rect 2455 3584 2467 3587
rect 4157 3587 4215 3593
rect 4157 3584 4169 3587
rect 2455 3556 4169 3584
rect 2455 3553 2467 3556
rect 2409 3547 2467 3553
rect 4157 3553 4169 3556
rect 4203 3584 4215 3587
rect 4709 3587 4767 3593
rect 4709 3584 4721 3587
rect 4203 3556 4721 3584
rect 4203 3553 4215 3556
rect 4157 3547 4215 3553
rect 4709 3553 4721 3556
rect 4755 3553 4767 3587
rect 4709 3547 4767 3553
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 1360 3488 1409 3516
rect 1360 3476 1366 3488
rect 1397 3485 1409 3488
rect 1443 3516 1455 3519
rect 1673 3519 1731 3525
rect 1673 3516 1685 3519
rect 1443 3488 1685 3516
rect 1443 3485 1455 3488
rect 1397 3479 1455 3485
rect 1673 3485 1685 3488
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 1964 3448 1992 3547
rect 2038 3476 2044 3528
rect 2096 3516 2102 3528
rect 2501 3519 2559 3525
rect 2501 3516 2513 3519
rect 2096 3488 2513 3516
rect 2096 3476 2102 3488
rect 2501 3485 2513 3488
rect 2547 3485 2559 3519
rect 2501 3479 2559 3485
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3485 2743 3519
rect 2685 3479 2743 3485
rect 2869 3519 2927 3525
rect 2869 3485 2881 3519
rect 2915 3516 2927 3519
rect 3881 3519 3939 3525
rect 3881 3516 3893 3519
rect 2915 3488 3893 3516
rect 2915 3485 2927 3488
rect 2869 3479 2927 3485
rect 3881 3485 3893 3488
rect 3927 3485 3939 3519
rect 3881 3479 3939 3485
rect 2700 3448 2728 3479
rect 3970 3476 3976 3528
rect 4028 3476 4034 3528
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 4801 3519 4859 3525
rect 4801 3485 4813 3519
rect 4847 3485 4859 3519
rect 5000 3516 5028 3624
rect 8757 3621 8769 3655
rect 8803 3652 8815 3655
rect 10505 3655 10563 3661
rect 8803 3624 10456 3652
rect 8803 3621 8815 3624
rect 8757 3615 8815 3621
rect 5074 3544 5080 3596
rect 5132 3584 5138 3596
rect 5132 3556 8156 3584
rect 5132 3544 5138 3556
rect 8128 3528 8156 3556
rect 8478 3544 8484 3596
rect 8536 3584 8542 3596
rect 9677 3587 9735 3593
rect 8536 3556 8984 3584
rect 8536 3544 8542 3556
rect 7929 3519 7987 3525
rect 7929 3516 7941 3519
rect 5000 3488 7941 3516
rect 4801 3479 4859 3485
rect 7929 3485 7941 3488
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 1964 3420 2728 3448
rect 3237 3451 3295 3457
rect 3237 3417 3249 3451
rect 3283 3417 3295 3451
rect 3237 3411 3295 3417
rect 3252 3380 3280 3411
rect 3326 3408 3332 3460
rect 3384 3448 3390 3460
rect 3421 3451 3479 3457
rect 3421 3448 3433 3451
rect 3384 3420 3433 3448
rect 3384 3408 3390 3420
rect 3421 3417 3433 3420
rect 3467 3417 3479 3451
rect 3786 3448 3792 3460
rect 3421 3411 3479 3417
rect 3528 3420 3792 3448
rect 3528 3380 3556 3420
rect 3786 3408 3792 3420
rect 3844 3448 3850 3460
rect 4080 3448 4108 3479
rect 3844 3420 4108 3448
rect 3844 3408 3850 3420
rect 4154 3408 4160 3460
rect 4212 3448 4218 3460
rect 4212 3420 4568 3448
rect 4212 3408 4218 3420
rect 3252 3352 3556 3380
rect 3605 3383 3663 3389
rect 3605 3349 3617 3383
rect 3651 3380 3663 3383
rect 4246 3380 4252 3392
rect 3651 3352 4252 3380
rect 3651 3349 3663 3352
rect 3605 3343 3663 3349
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 4430 3340 4436 3392
rect 4488 3340 4494 3392
rect 4540 3380 4568 3420
rect 4706 3408 4712 3460
rect 4764 3448 4770 3460
rect 4816 3448 4844 3479
rect 4764 3420 4844 3448
rect 4764 3408 4770 3420
rect 4982 3380 4988 3392
rect 4540 3352 4988 3380
rect 4982 3340 4988 3352
rect 5040 3340 5046 3392
rect 7944 3380 7972 3479
rect 8110 3476 8116 3528
rect 8168 3476 8174 3528
rect 8956 3525 8984 3556
rect 9677 3553 9689 3587
rect 9723 3584 9735 3587
rect 10321 3587 10379 3593
rect 10321 3584 10333 3587
rect 9723 3556 10333 3584
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 10321 3553 10333 3556
rect 10367 3553 10379 3587
rect 10321 3547 10379 3553
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 8941 3519 8999 3525
rect 8941 3485 8953 3519
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 8021 3451 8079 3457
rect 8021 3417 8033 3451
rect 8067 3448 8079 3451
rect 8404 3448 8432 3479
rect 9214 3476 9220 3528
rect 9272 3516 9278 3528
rect 9585 3519 9643 3525
rect 9585 3516 9597 3519
rect 9272 3488 9597 3516
rect 9272 3476 9278 3488
rect 9585 3485 9597 3488
rect 9631 3485 9643 3519
rect 9585 3479 9643 3485
rect 9766 3476 9772 3528
rect 9824 3476 9830 3528
rect 9953 3519 10011 3525
rect 9953 3485 9965 3519
rect 9999 3516 10011 3519
rect 10042 3516 10048 3528
rect 9999 3488 10048 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 10229 3519 10287 3525
rect 10229 3485 10241 3519
rect 10275 3516 10287 3519
rect 10428 3516 10456 3624
rect 10505 3621 10517 3655
rect 10551 3652 10563 3655
rect 10551 3624 12434 3652
rect 10551 3621 10563 3624
rect 10505 3615 10563 3621
rect 10686 3544 10692 3596
rect 10744 3584 10750 3596
rect 11882 3584 11888 3596
rect 10744 3556 11888 3584
rect 10744 3544 10750 3556
rect 11882 3544 11888 3556
rect 11940 3584 11946 3596
rect 11977 3587 12035 3593
rect 11977 3584 11989 3587
rect 11940 3556 11989 3584
rect 11940 3544 11946 3556
rect 11977 3553 11989 3556
rect 12023 3553 12035 3587
rect 12406 3584 12434 3624
rect 12618 3584 12624 3596
rect 12406 3556 12624 3584
rect 11977 3547 12035 3553
rect 10870 3516 10876 3528
rect 10275 3488 10876 3516
rect 10275 3485 10287 3488
rect 10229 3479 10287 3485
rect 10870 3476 10876 3488
rect 10928 3476 10934 3528
rect 12342 3476 12348 3528
rect 12400 3476 12406 3528
rect 12452 3525 12480 3556
rect 12618 3544 12624 3556
rect 12676 3544 12682 3596
rect 17773 3587 17831 3593
rect 17773 3553 17785 3587
rect 17819 3584 17831 3587
rect 18414 3584 18420 3596
rect 17819 3556 18420 3584
rect 17819 3553 17831 3556
rect 17773 3547 17831 3553
rect 18414 3544 18420 3556
rect 18472 3544 18478 3596
rect 12437 3519 12495 3525
rect 12437 3485 12449 3519
rect 12483 3516 12495 3519
rect 12483 3488 12517 3516
rect 12483 3485 12495 3488
rect 12437 3479 12495 3485
rect 17494 3476 17500 3528
rect 17552 3476 17558 3528
rect 18046 3476 18052 3528
rect 18104 3476 18110 3528
rect 8478 3448 8484 3460
rect 8067 3420 8484 3448
rect 8067 3417 8079 3420
rect 8021 3411 8079 3417
rect 8478 3408 8484 3420
rect 8536 3408 8542 3460
rect 9861 3451 9919 3457
rect 9861 3448 9873 3451
rect 9508 3420 9873 3448
rect 8294 3380 8300 3392
rect 7944 3352 8300 3380
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 9508 3389 9536 3420
rect 9861 3417 9873 3420
rect 9907 3417 9919 3451
rect 9861 3411 9919 3417
rect 18322 3408 18328 3460
rect 18380 3408 18386 3460
rect 9493 3383 9551 3389
rect 9493 3349 9505 3383
rect 9539 3349 9551 3383
rect 9493 3343 9551 3349
rect 1104 3290 18860 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 18860 3290
rect 1104 3216 18860 3238
rect 2133 3179 2191 3185
rect 2133 3145 2145 3179
rect 2179 3145 2191 3179
rect 2133 3139 2191 3145
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3040 2099 3043
rect 2148 3040 2176 3139
rect 2590 3136 2596 3188
rect 2648 3136 2654 3188
rect 4430 3176 4436 3188
rect 2746 3148 4436 3176
rect 2501 3111 2559 3117
rect 2501 3077 2513 3111
rect 2547 3108 2559 3111
rect 2746 3108 2774 3148
rect 4430 3136 4436 3148
rect 4488 3136 4494 3188
rect 5350 3136 5356 3188
rect 5408 3136 5414 3188
rect 7745 3179 7803 3185
rect 7745 3145 7757 3179
rect 7791 3176 7803 3179
rect 9214 3176 9220 3188
rect 7791 3148 9220 3176
rect 7791 3145 7803 3148
rect 7745 3139 7803 3145
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 9953 3179 10011 3185
rect 9953 3176 9965 3179
rect 9824 3148 9965 3176
rect 9824 3136 9830 3148
rect 9953 3145 9965 3148
rect 9999 3145 10011 3179
rect 9953 3139 10011 3145
rect 10042 3136 10048 3188
rect 10100 3176 10106 3188
rect 10781 3179 10839 3185
rect 10781 3176 10793 3179
rect 10100 3148 10793 3176
rect 10100 3136 10106 3148
rect 10781 3145 10793 3148
rect 10827 3145 10839 3179
rect 10781 3139 10839 3145
rect 10870 3136 10876 3188
rect 10928 3136 10934 3188
rect 11882 3136 11888 3188
rect 11940 3136 11946 3188
rect 11977 3179 12035 3185
rect 11977 3145 11989 3179
rect 12023 3176 12035 3179
rect 12342 3176 12348 3188
rect 12023 3148 12348 3176
rect 12023 3145 12035 3148
rect 11977 3139 12035 3145
rect 12342 3136 12348 3148
rect 12400 3136 12406 3188
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 12713 3179 12771 3185
rect 12713 3176 12725 3179
rect 12492 3148 12725 3176
rect 12492 3136 12498 3148
rect 12713 3145 12725 3148
rect 12759 3145 12771 3179
rect 12713 3139 12771 3145
rect 13078 3136 13084 3188
rect 13136 3176 13142 3188
rect 13541 3179 13599 3185
rect 13541 3176 13553 3179
rect 13136 3148 13553 3176
rect 13136 3136 13142 3148
rect 13541 3145 13553 3148
rect 13587 3145 13599 3179
rect 13541 3139 13599 3145
rect 4614 3108 4620 3120
rect 2547 3080 2774 3108
rect 3344 3080 4108 3108
rect 2547 3077 2559 3080
rect 2501 3071 2559 3077
rect 3344 3040 3372 3080
rect 2087 3012 2176 3040
rect 2700 3012 3372 3040
rect 3421 3043 3479 3049
rect 2087 3009 2099 3012
rect 2041 3003 2099 3009
rect 1854 2932 1860 2984
rect 1912 2932 1918 2984
rect 2590 2932 2596 2984
rect 2648 2972 2654 2984
rect 2700 2981 2728 3012
rect 3421 3009 3433 3043
rect 3467 3009 3479 3043
rect 3421 3003 3479 3009
rect 2685 2975 2743 2981
rect 2685 2972 2697 2975
rect 2648 2944 2697 2972
rect 2648 2932 2654 2944
rect 2685 2941 2697 2944
rect 2731 2941 2743 2975
rect 2685 2935 2743 2941
rect 3145 2975 3203 2981
rect 3145 2941 3157 2975
rect 3191 2941 3203 2975
rect 3145 2935 3203 2941
rect 2498 2864 2504 2916
rect 2556 2904 2562 2916
rect 3160 2904 3188 2935
rect 2556 2876 3188 2904
rect 3436 2904 3464 3003
rect 3602 2932 3608 2984
rect 3660 2972 3666 2984
rect 3881 2975 3939 2981
rect 3881 2972 3893 2975
rect 3660 2944 3893 2972
rect 3660 2932 3666 2944
rect 3881 2941 3893 2944
rect 3927 2941 3939 2975
rect 4080 2972 4108 3080
rect 4172 3080 4620 3108
rect 4172 3049 4200 3080
rect 4614 3068 4620 3080
rect 4672 3068 4678 3120
rect 5261 3111 5319 3117
rect 5261 3077 5273 3111
rect 5307 3108 5319 3111
rect 5442 3108 5448 3120
rect 5307 3080 5448 3108
rect 5307 3077 5319 3080
rect 5261 3071 5319 3077
rect 5442 3068 5448 3080
rect 5500 3068 5506 3120
rect 6638 3068 6644 3120
rect 6696 3068 6702 3120
rect 8110 3108 8116 3120
rect 7392 3080 8116 3108
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 4246 3000 4252 3052
rect 4304 3040 4310 3052
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 4304 3012 4445 3040
rect 4304 3000 4310 3012
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 5626 3040 5632 3052
rect 4433 3003 4491 3009
rect 4540 3012 5632 3040
rect 4540 2972 4568 3012
rect 4080 2944 4568 2972
rect 3881 2935 3939 2941
rect 4614 2932 4620 2984
rect 4672 2932 4678 2984
rect 5460 2981 5488 3012
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 6457 3043 6515 3049
rect 6457 3009 6469 3043
rect 6503 3040 6515 3043
rect 6656 3040 6684 3068
rect 7392 3049 7420 3080
rect 8110 3068 8116 3080
rect 8168 3108 8174 3120
rect 8205 3111 8263 3117
rect 8205 3108 8217 3111
rect 8168 3080 8217 3108
rect 8168 3068 8174 3080
rect 8205 3077 8217 3080
rect 8251 3077 8263 3111
rect 8205 3071 8263 3077
rect 12526 3068 12532 3120
rect 12584 3108 12590 3120
rect 12805 3111 12863 3117
rect 12805 3108 12817 3111
rect 12584 3080 12817 3108
rect 12584 3068 12590 3080
rect 12805 3077 12817 3080
rect 12851 3077 12863 3111
rect 12805 3071 12863 3077
rect 12894 3068 12900 3120
rect 12952 3108 12958 3120
rect 13633 3111 13691 3117
rect 13633 3108 13645 3111
rect 12952 3080 13645 3108
rect 12952 3068 12958 3080
rect 13633 3077 13645 3080
rect 13679 3077 13691 3111
rect 13633 3071 13691 3077
rect 6503 3012 6684 3040
rect 7377 3043 7435 3049
rect 6503 3009 6515 3012
rect 6457 3003 6515 3009
rect 7377 3009 7389 3043
rect 7423 3009 7435 3043
rect 8021 3043 8079 3049
rect 8021 3040 8033 3043
rect 7377 3003 7435 3009
rect 7484 3012 8033 3040
rect 5445 2975 5503 2981
rect 5445 2941 5457 2975
rect 5491 2941 5503 2975
rect 5445 2935 5503 2941
rect 6362 2932 6368 2984
rect 6420 2972 6426 2984
rect 7484 2981 7512 3012
rect 8021 3009 8033 3012
rect 8067 3040 8079 3043
rect 8294 3040 8300 3052
rect 8067 3012 8300 3040
rect 8067 3009 8079 3012
rect 8021 3003 8079 3009
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 8389 3043 8447 3049
rect 8389 3009 8401 3043
rect 8435 3040 8447 3043
rect 8665 3043 8723 3049
rect 8665 3040 8677 3043
rect 8435 3012 8677 3040
rect 8435 3009 8447 3012
rect 8389 3003 8447 3009
rect 8665 3009 8677 3012
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 8849 3043 8907 3049
rect 8849 3009 8861 3043
rect 8895 3040 8907 3043
rect 10045 3043 10103 3049
rect 10045 3040 10057 3043
rect 8895 3012 10057 3040
rect 8895 3009 8907 3012
rect 8849 3003 8907 3009
rect 10045 3009 10057 3012
rect 10091 3009 10103 3043
rect 17497 3043 17555 3049
rect 10045 3003 10103 3009
rect 12406 3012 13032 3040
rect 6641 2975 6699 2981
rect 6641 2972 6653 2975
rect 6420 2944 6653 2972
rect 6420 2932 6426 2944
rect 6641 2941 6653 2944
rect 6687 2941 6699 2975
rect 6641 2935 6699 2941
rect 7469 2975 7527 2981
rect 7469 2941 7481 2975
rect 7515 2941 7527 2975
rect 7469 2935 7527 2941
rect 8478 2932 8484 2984
rect 8536 2932 8542 2984
rect 9861 2975 9919 2981
rect 9861 2941 9873 2975
rect 9907 2941 9919 2975
rect 9861 2935 9919 2941
rect 10597 2975 10655 2981
rect 10597 2941 10609 2975
rect 10643 2941 10655 2975
rect 10597 2935 10655 2941
rect 12069 2975 12127 2981
rect 12069 2941 12081 2975
rect 12115 2972 12127 2975
rect 12406 2972 12434 3012
rect 13004 2981 13032 3012
rect 17497 3009 17509 3043
rect 17543 3040 17555 3043
rect 17586 3040 17592 3052
rect 17543 3012 17592 3040
rect 17543 3009 17555 3012
rect 17497 3003 17555 3009
rect 17586 3000 17592 3012
rect 17644 3000 17650 3052
rect 18506 3000 18512 3052
rect 18564 3000 18570 3052
rect 12115 2944 12434 2972
rect 12989 2975 13047 2981
rect 12115 2941 12127 2944
rect 12069 2935 12127 2941
rect 12989 2941 13001 2975
rect 13035 2972 13047 2975
rect 13725 2975 13783 2981
rect 13725 2972 13737 2975
rect 13035 2944 13737 2972
rect 13035 2941 13047 2944
rect 12989 2935 13047 2941
rect 13725 2941 13737 2944
rect 13771 2972 13783 2975
rect 14734 2972 14740 2984
rect 13771 2944 14740 2972
rect 13771 2941 13783 2944
rect 13725 2935 13783 2941
rect 4893 2907 4951 2913
rect 4893 2904 4905 2907
rect 3436 2876 4905 2904
rect 2556 2864 2562 2876
rect 4893 2873 4905 2876
rect 4939 2873 4951 2907
rect 9876 2904 9904 2935
rect 10612 2904 10640 2935
rect 12084 2904 12112 2935
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 17402 2932 17408 2984
rect 17460 2972 17466 2984
rect 17681 2975 17739 2981
rect 17681 2972 17693 2975
rect 17460 2944 17693 2972
rect 17460 2932 17466 2944
rect 17681 2941 17693 2944
rect 17727 2941 17739 2975
rect 17681 2935 17739 2941
rect 17954 2932 17960 2984
rect 18012 2972 18018 2984
rect 18233 2975 18291 2981
rect 18233 2972 18245 2975
rect 18012 2944 18245 2972
rect 18012 2932 18018 2944
rect 18233 2941 18245 2944
rect 18279 2941 18291 2975
rect 18233 2935 18291 2941
rect 9876 2876 12112 2904
rect 4893 2867 4951 2873
rect 12526 2864 12532 2916
rect 12584 2904 12590 2916
rect 13173 2907 13231 2913
rect 13173 2904 13185 2907
rect 12584 2876 13185 2904
rect 12584 2864 12590 2876
rect 13173 2873 13185 2876
rect 13219 2873 13231 2907
rect 13173 2867 13231 2873
rect 3970 2796 3976 2848
rect 4028 2836 4034 2848
rect 4249 2839 4307 2845
rect 4249 2836 4261 2839
rect 4028 2808 4261 2836
rect 4028 2796 4034 2808
rect 4249 2805 4261 2808
rect 4295 2805 4307 2839
rect 4249 2799 4307 2805
rect 10318 2796 10324 2848
rect 10376 2836 10382 2848
rect 10413 2839 10471 2845
rect 10413 2836 10425 2839
rect 10376 2808 10425 2836
rect 10376 2796 10382 2808
rect 10413 2805 10425 2808
rect 10459 2805 10471 2839
rect 10413 2799 10471 2805
rect 11241 2839 11299 2845
rect 11241 2805 11253 2839
rect 11287 2836 11299 2839
rect 11330 2836 11336 2848
rect 11287 2808 11336 2836
rect 11287 2805 11299 2808
rect 11241 2799 11299 2805
rect 11330 2796 11336 2808
rect 11388 2796 11394 2848
rect 11514 2796 11520 2848
rect 11572 2796 11578 2848
rect 12345 2839 12403 2845
rect 12345 2805 12357 2839
rect 12391 2836 12403 2839
rect 12618 2836 12624 2848
rect 12391 2808 12624 2836
rect 12391 2805 12403 2808
rect 12345 2799 12403 2805
rect 12618 2796 12624 2808
rect 12676 2796 12682 2848
rect 1104 2746 18860 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 18860 2746
rect 1104 2672 18860 2694
rect 1578 2592 1584 2644
rect 1636 2592 1642 2644
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 1946 2632 1952 2644
rect 1903 2604 1952 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 3786 2632 3792 2644
rect 2915 2604 3792 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 3786 2592 3792 2604
rect 3844 2592 3850 2644
rect 3881 2635 3939 2641
rect 3881 2601 3893 2635
rect 3927 2632 3939 2635
rect 4614 2632 4620 2644
rect 3927 2604 4620 2632
rect 3927 2601 3939 2604
rect 3881 2595 3939 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 8110 2564 8116 2576
rect 5644 2536 8116 2564
rect 2314 2456 2320 2508
rect 2372 2456 2378 2508
rect 2501 2499 2559 2505
rect 2501 2465 2513 2499
rect 2547 2496 2559 2499
rect 2590 2496 2596 2508
rect 2547 2468 2596 2496
rect 2547 2465 2559 2468
rect 2501 2459 2559 2465
rect 2590 2456 2596 2468
rect 2648 2456 2654 2508
rect 4062 2496 4068 2508
rect 3620 2468 4068 2496
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 3620 2437 3648 2468
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 4706 2456 4712 2508
rect 4764 2456 4770 2508
rect 5258 2456 5264 2508
rect 5316 2456 5322 2508
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 1360 2400 1409 2428
rect 1360 2388 1366 2400
rect 1397 2397 1409 2400
rect 1443 2428 1455 2431
rect 1673 2431 1731 2437
rect 1673 2428 1685 2431
rect 1443 2400 1685 2428
rect 1443 2397 1455 2400
rect 1397 2391 1455 2397
rect 1673 2397 1685 2400
rect 1719 2397 1731 2431
rect 1673 2391 1731 2397
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2397 3663 2431
rect 3605 2391 3663 2397
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 2700 2360 2728 2391
rect 3786 2388 3792 2440
rect 3844 2388 3850 2440
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3936 2400 3985 2428
rect 3936 2388 3942 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4525 2431 4583 2437
rect 4525 2397 4537 2431
rect 4571 2428 4583 2431
rect 4724 2428 4752 2456
rect 4571 2400 4752 2428
rect 5077 2431 5135 2437
rect 4571 2397 4583 2400
rect 4525 2391 4583 2397
rect 5077 2397 5089 2431
rect 5123 2428 5135 2431
rect 5276 2428 5304 2456
rect 5644 2437 5672 2536
rect 8110 2524 8116 2536
rect 8168 2524 8174 2576
rect 5810 2456 5816 2508
rect 5868 2456 5874 2508
rect 11422 2496 11428 2508
rect 10244 2468 11428 2496
rect 5123 2400 5304 2428
rect 5629 2431 5687 2437
rect 5123 2397 5135 2400
rect 5077 2391 5135 2397
rect 5629 2397 5641 2431
rect 5675 2397 5687 2431
rect 5629 2391 5687 2397
rect 5718 2388 5724 2440
rect 5776 2388 5782 2440
rect 5828 2428 5856 2456
rect 6641 2431 6699 2437
rect 6641 2428 6653 2431
rect 5828 2400 6653 2428
rect 6641 2397 6653 2400
rect 6687 2397 6699 2431
rect 6641 2391 6699 2397
rect 7650 2388 7656 2440
rect 7708 2388 7714 2440
rect 8202 2388 8208 2440
rect 8260 2388 8266 2440
rect 8754 2388 8760 2440
rect 8812 2388 8818 2440
rect 9677 2431 9735 2437
rect 9677 2397 9689 2431
rect 9723 2428 9735 2431
rect 9766 2428 9772 2440
rect 9723 2400 9772 2428
rect 9723 2397 9735 2400
rect 9677 2391 9735 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 10244 2437 10272 2468
rect 11422 2456 11428 2468
rect 11480 2456 11486 2508
rect 14734 2456 14740 2508
rect 14792 2496 14798 2508
rect 15381 2499 15439 2505
rect 15381 2496 15393 2499
rect 14792 2468 15393 2496
rect 14792 2456 14798 2468
rect 15381 2465 15393 2468
rect 15427 2465 15439 2499
rect 15381 2459 15439 2465
rect 15746 2456 15752 2508
rect 15804 2496 15810 2508
rect 15804 2468 16804 2496
rect 15804 2456 15810 2468
rect 10229 2431 10287 2437
rect 10229 2397 10241 2431
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 10318 2388 10324 2440
rect 10376 2388 10382 2440
rect 11330 2388 11336 2440
rect 11388 2388 11394 2440
rect 11514 2388 11520 2440
rect 11572 2388 11578 2440
rect 12526 2388 12532 2440
rect 12584 2388 12590 2440
rect 12618 2388 12624 2440
rect 12676 2388 12682 2440
rect 13630 2388 13636 2440
rect 13688 2388 13694 2440
rect 14090 2388 14096 2440
rect 14148 2388 14154 2440
rect 14642 2388 14648 2440
rect 14700 2388 14706 2440
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2428 15255 2431
rect 15562 2428 15568 2440
rect 15243 2400 15568 2428
rect 15243 2397 15255 2400
rect 15197 2391 15255 2397
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 16206 2388 16212 2440
rect 16264 2388 16270 2440
rect 16666 2388 16672 2440
rect 16724 2388 16730 2440
rect 16776 2428 16804 2468
rect 16945 2431 17003 2437
rect 16945 2428 16957 2431
rect 16776 2400 16957 2428
rect 16945 2397 16957 2400
rect 16991 2397 17003 2431
rect 16945 2391 17003 2397
rect 17218 2388 17224 2440
rect 17276 2388 17282 2440
rect 17770 2388 17776 2440
rect 17828 2388 17834 2440
rect 2961 2363 3019 2369
rect 2961 2360 2973 2363
rect 1268 2332 2973 2360
rect 1268 2320 1274 2332
rect 2961 2329 2973 2332
rect 3007 2329 3019 2363
rect 2961 2323 3019 2329
rect 3050 2320 3056 2372
rect 3108 2360 3114 2372
rect 3329 2363 3387 2369
rect 3329 2360 3341 2363
rect 3108 2332 3341 2360
rect 3108 2320 3114 2332
rect 3329 2329 3341 2332
rect 3375 2329 3387 2363
rect 3329 2323 3387 2329
rect 4154 2320 4160 2372
rect 4212 2360 4218 2372
rect 4249 2363 4307 2369
rect 4249 2360 4261 2363
rect 4212 2332 4261 2360
rect 4212 2320 4218 2332
rect 4249 2329 4261 2332
rect 4295 2329 4307 2363
rect 4249 2323 4307 2329
rect 4706 2320 4712 2372
rect 4764 2360 4770 2372
rect 4801 2363 4859 2369
rect 4801 2360 4813 2363
rect 4764 2332 4813 2360
rect 4764 2320 4770 2332
rect 4801 2329 4813 2332
rect 4847 2329 4859 2363
rect 4801 2323 4859 2329
rect 5258 2320 5264 2372
rect 5316 2360 5322 2372
rect 5353 2363 5411 2369
rect 5353 2360 5365 2363
rect 5316 2332 5365 2360
rect 5316 2320 5322 2332
rect 5353 2329 5365 2332
rect 5399 2329 5411 2363
rect 5353 2323 5411 2329
rect 5810 2320 5816 2372
rect 5868 2360 5874 2372
rect 5997 2363 6055 2369
rect 5997 2360 6009 2363
rect 5868 2332 6009 2360
rect 5868 2320 5874 2332
rect 5997 2329 6009 2332
rect 6043 2329 6055 2363
rect 5997 2323 6055 2329
rect 6914 2320 6920 2372
rect 6972 2320 6978 2372
rect 7377 2363 7435 2369
rect 7377 2329 7389 2363
rect 7423 2360 7435 2363
rect 7466 2360 7472 2372
rect 7423 2332 7472 2360
rect 7423 2329 7435 2332
rect 7377 2323 7435 2329
rect 7466 2320 7472 2332
rect 7524 2320 7530 2372
rect 7929 2363 7987 2369
rect 7929 2329 7941 2363
rect 7975 2360 7987 2363
rect 8018 2360 8024 2372
rect 7975 2332 8024 2360
rect 7975 2329 7987 2332
rect 7929 2323 7987 2329
rect 8018 2320 8024 2332
rect 8076 2320 8082 2372
rect 8481 2363 8539 2369
rect 8481 2329 8493 2363
rect 8527 2360 8539 2363
rect 8570 2360 8576 2372
rect 8527 2332 8576 2360
rect 8527 2329 8539 2332
rect 8481 2323 8539 2329
rect 8570 2320 8576 2332
rect 8628 2320 8634 2372
rect 9122 2320 9128 2372
rect 9180 2360 9186 2372
rect 9401 2363 9459 2369
rect 9401 2360 9413 2363
rect 9180 2332 9413 2360
rect 9180 2320 9186 2332
rect 9401 2329 9413 2332
rect 9447 2329 9459 2363
rect 9953 2363 10011 2369
rect 9953 2360 9965 2363
rect 9401 2323 9459 2329
rect 9692 2332 9965 2360
rect 9692 2304 9720 2332
rect 9953 2329 9965 2332
rect 9999 2329 10011 2363
rect 10597 2363 10655 2369
rect 10597 2360 10609 2363
rect 9953 2323 10011 2329
rect 10244 2332 10609 2360
rect 10244 2304 10272 2332
rect 10597 2329 10609 2332
rect 10643 2329 10655 2363
rect 10597 2323 10655 2329
rect 10778 2320 10784 2372
rect 10836 2360 10842 2372
rect 11057 2363 11115 2369
rect 11057 2360 11069 2363
rect 10836 2332 11069 2360
rect 10836 2320 10842 2332
rect 11057 2329 11069 2332
rect 11103 2329 11115 2363
rect 11793 2363 11851 2369
rect 11793 2360 11805 2363
rect 11057 2323 11115 2329
rect 11348 2332 11805 2360
rect 11348 2304 11376 2332
rect 11793 2329 11805 2332
rect 11839 2329 11851 2363
rect 11793 2323 11851 2329
rect 11882 2320 11888 2372
rect 11940 2360 11946 2372
rect 12253 2363 12311 2369
rect 12253 2360 12265 2363
rect 11940 2332 12265 2360
rect 11940 2320 11946 2332
rect 12253 2329 12265 2332
rect 12299 2329 12311 2363
rect 12253 2323 12311 2329
rect 12434 2320 12440 2372
rect 12492 2360 12498 2372
rect 12897 2363 12955 2369
rect 12897 2360 12909 2363
rect 12492 2332 12909 2360
rect 12492 2320 12498 2332
rect 12897 2329 12909 2332
rect 12943 2329 12955 2363
rect 12897 2323 12955 2329
rect 12986 2320 12992 2372
rect 13044 2360 13050 2372
rect 13357 2363 13415 2369
rect 13357 2360 13369 2363
rect 13044 2332 13369 2360
rect 13044 2320 13050 2332
rect 13357 2329 13369 2332
rect 13403 2329 13415 2363
rect 13357 2323 13415 2329
rect 13538 2320 13544 2372
rect 13596 2360 13602 2372
rect 14369 2363 14427 2369
rect 14369 2360 14381 2363
rect 13596 2332 14381 2360
rect 13596 2320 13602 2332
rect 14369 2329 14381 2332
rect 14415 2329 14427 2363
rect 14369 2323 14427 2329
rect 14921 2363 14979 2369
rect 14921 2329 14933 2363
rect 14967 2329 14979 2363
rect 14921 2323 14979 2329
rect 15933 2363 15991 2369
rect 15933 2329 15945 2363
rect 15979 2329 15991 2363
rect 15933 2323 15991 2329
rect 2225 2295 2283 2301
rect 2225 2261 2237 2295
rect 2271 2292 2283 2295
rect 3418 2292 3424 2304
rect 2271 2264 3424 2292
rect 2271 2261 2283 2264
rect 2225 2255 2283 2261
rect 3418 2252 3424 2264
rect 3476 2292 3482 2304
rect 3970 2292 3976 2304
rect 3476 2264 3976 2292
rect 3476 2252 3482 2264
rect 3970 2252 3976 2264
rect 4028 2252 4034 2304
rect 9674 2252 9680 2304
rect 9732 2252 9738 2304
rect 10226 2252 10232 2304
rect 10284 2252 10290 2304
rect 11330 2252 11336 2304
rect 11388 2252 11394 2304
rect 14090 2252 14096 2304
rect 14148 2292 14154 2304
rect 14936 2292 14964 2323
rect 14148 2264 14964 2292
rect 14148 2252 14154 2264
rect 15194 2252 15200 2304
rect 15252 2292 15258 2304
rect 15948 2292 15976 2323
rect 16298 2320 16304 2372
rect 16356 2360 16362 2372
rect 17497 2363 17555 2369
rect 17497 2360 17509 2363
rect 16356 2332 17509 2360
rect 16356 2320 16362 2332
rect 17497 2329 17509 2332
rect 17543 2329 17555 2363
rect 17497 2323 17555 2329
rect 18049 2363 18107 2369
rect 18049 2329 18061 2363
rect 18095 2329 18107 2363
rect 18049 2323 18107 2329
rect 15252 2264 15976 2292
rect 15252 2252 15258 2264
rect 16850 2252 16856 2304
rect 16908 2292 16914 2304
rect 18064 2292 18092 2323
rect 16908 2264 18092 2292
rect 16908 2252 16914 2264
rect 1104 2202 18860 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 18860 2202
rect 1104 2128 18860 2150
<< via1 >>
rect 7012 17688 7064 17740
rect 15016 17688 15068 17740
rect 12256 17552 12308 17604
rect 16764 17552 16816 17604
rect 7748 17484 7800 17536
rect 15384 17484 15436 17536
rect 15752 17484 15804 17536
rect 16488 17484 16540 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 2504 17323 2556 17332
rect 2504 17289 2513 17323
rect 2513 17289 2547 17323
rect 2547 17289 2556 17323
rect 2504 17280 2556 17289
rect 3056 17323 3108 17332
rect 3056 17289 3065 17323
rect 3065 17289 3099 17323
rect 3099 17289 3108 17323
rect 3056 17280 3108 17289
rect 3608 17323 3660 17332
rect 3608 17289 3617 17323
rect 3617 17289 3651 17323
rect 3651 17289 3660 17323
rect 3608 17280 3660 17289
rect 1952 17212 2004 17264
rect 1492 17187 1544 17196
rect 1492 17153 1501 17187
rect 1501 17153 1535 17187
rect 1535 17153 1544 17187
rect 1492 17144 1544 17153
rect 1308 17076 1360 17128
rect 3424 17144 3476 17196
rect 6736 17280 6788 17332
rect 7012 17280 7064 17332
rect 7472 17323 7524 17332
rect 7472 17289 7481 17323
rect 7481 17289 7515 17323
rect 7515 17289 7524 17323
rect 7472 17280 7524 17289
rect 8024 17323 8076 17332
rect 8024 17289 8033 17323
rect 8033 17289 8067 17323
rect 8067 17289 8076 17323
rect 8024 17280 8076 17289
rect 4160 17212 4212 17264
rect 6368 17212 6420 17264
rect 6920 17212 6972 17264
rect 4712 17144 4764 17196
rect 5264 17144 5316 17196
rect 5908 17144 5960 17196
rect 1676 16983 1728 16992
rect 1676 16949 1685 16983
rect 1685 16949 1719 16983
rect 1719 16949 1728 16983
rect 1676 16940 1728 16949
rect 2044 16940 2096 16992
rect 3516 16940 3568 16992
rect 3884 16940 3936 16992
rect 4620 17008 4672 17060
rect 6552 17144 6604 17196
rect 7012 17187 7064 17196
rect 7012 17153 7021 17187
rect 7021 17153 7055 17187
rect 7055 17153 7064 17187
rect 7012 17144 7064 17153
rect 8576 17323 8628 17332
rect 8576 17289 8585 17323
rect 8585 17289 8619 17323
rect 8619 17289 8628 17323
rect 8576 17280 8628 17289
rect 9680 17323 9732 17332
rect 9680 17289 9689 17323
rect 9689 17289 9723 17323
rect 9723 17289 9732 17323
rect 9680 17280 9732 17289
rect 10232 17323 10284 17332
rect 10232 17289 10241 17323
rect 10241 17289 10275 17323
rect 10275 17289 10284 17323
rect 10232 17280 10284 17289
rect 9128 17144 9180 17196
rect 10784 17280 10836 17332
rect 12992 17280 13044 17332
rect 14004 17280 14056 17332
rect 15200 17280 15252 17332
rect 16028 17280 16080 17332
rect 16856 17280 16908 17332
rect 11336 17144 11388 17196
rect 12440 17144 12492 17196
rect 6644 17076 6696 17128
rect 11704 17076 11756 17128
rect 11796 17119 11848 17128
rect 11796 17085 11805 17119
rect 11805 17085 11839 17119
rect 11839 17085 11848 17119
rect 11796 17076 11848 17085
rect 12808 17119 12860 17128
rect 12808 17085 12817 17119
rect 12817 17085 12851 17119
rect 12851 17085 12860 17119
rect 12808 17076 12860 17085
rect 6276 17008 6328 17060
rect 10048 17008 10100 17060
rect 10692 17008 10744 17060
rect 11888 17008 11940 17060
rect 13268 17144 13320 17196
rect 13912 17144 13964 17196
rect 14096 17144 14148 17196
rect 14648 17144 14700 17196
rect 15108 17144 15160 17196
rect 15660 17187 15712 17196
rect 15660 17153 15669 17187
rect 15669 17153 15703 17187
rect 15703 17153 15712 17187
rect 15660 17144 15712 17153
rect 15752 17187 15804 17196
rect 15752 17153 15761 17187
rect 15761 17153 15795 17187
rect 15795 17153 15804 17187
rect 15752 17144 15804 17153
rect 15936 17187 15988 17196
rect 15936 17153 15945 17187
rect 15945 17153 15979 17187
rect 15979 17153 15988 17187
rect 15936 17144 15988 17153
rect 16028 17144 16080 17196
rect 16488 17212 16540 17264
rect 16764 17144 16816 17196
rect 18512 17187 18564 17196
rect 18512 17153 18521 17187
rect 18521 17153 18555 17187
rect 18555 17153 18564 17187
rect 18512 17144 18564 17153
rect 14464 17119 14516 17128
rect 14464 17085 14473 17119
rect 14473 17085 14507 17119
rect 14507 17085 14516 17119
rect 14464 17076 14516 17085
rect 16212 17076 16264 17128
rect 15016 17008 15068 17060
rect 15292 17008 15344 17060
rect 4804 16940 4856 16992
rect 5356 16940 5408 16992
rect 5908 16940 5960 16992
rect 6920 16983 6972 16992
rect 6920 16949 6929 16983
rect 6929 16949 6963 16983
rect 6963 16949 6972 16983
rect 6920 16940 6972 16949
rect 7564 16940 7616 16992
rect 7932 16940 7984 16992
rect 9036 16940 9088 16992
rect 9588 16940 9640 16992
rect 10232 16940 10284 16992
rect 11336 16983 11388 16992
rect 11336 16949 11345 16983
rect 11345 16949 11379 16983
rect 11379 16949 11388 16983
rect 11336 16940 11388 16949
rect 12900 16940 12952 16992
rect 13912 16983 13964 16992
rect 13912 16949 13921 16983
rect 13921 16949 13955 16983
rect 13955 16949 13964 16983
rect 13912 16940 13964 16949
rect 14648 16940 14700 16992
rect 15568 16940 15620 16992
rect 16028 16940 16080 16992
rect 16120 16983 16172 16992
rect 16120 16949 16129 16983
rect 16129 16949 16163 16983
rect 16163 16949 16172 16983
rect 16120 16940 16172 16949
rect 16672 16940 16724 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 1952 16779 2004 16788
rect 1952 16745 1961 16779
rect 1961 16745 1995 16779
rect 1995 16745 2004 16779
rect 1952 16736 2004 16745
rect 4160 16779 4212 16788
rect 4160 16745 4169 16779
rect 4169 16745 4203 16779
rect 4203 16745 4212 16779
rect 4160 16736 4212 16745
rect 4712 16779 4764 16788
rect 4712 16745 4721 16779
rect 4721 16745 4755 16779
rect 4755 16745 4764 16779
rect 4712 16736 4764 16745
rect 7012 16736 7064 16788
rect 12256 16779 12308 16788
rect 12256 16745 12265 16779
rect 12265 16745 12299 16779
rect 12299 16745 12308 16779
rect 12256 16736 12308 16745
rect 1676 16668 1728 16720
rect 1308 16600 1360 16652
rect 1400 16575 1452 16584
rect 1400 16541 1409 16575
rect 1409 16541 1443 16575
rect 1443 16541 1452 16575
rect 1400 16532 1452 16541
rect 5816 16532 5868 16584
rect 6644 16532 6696 16584
rect 6920 16600 6972 16652
rect 7748 16643 7800 16652
rect 7748 16609 7757 16643
rect 7757 16609 7791 16643
rect 7791 16609 7800 16643
rect 7748 16600 7800 16609
rect 8760 16643 8812 16652
rect 8760 16609 8769 16643
rect 8769 16609 8803 16643
rect 8803 16609 8812 16643
rect 8760 16600 8812 16609
rect 9220 16668 9272 16720
rect 12716 16736 12768 16788
rect 9956 16600 10008 16652
rect 7012 16575 7064 16584
rect 7012 16541 7021 16575
rect 7021 16541 7055 16575
rect 7055 16541 7064 16575
rect 7012 16532 7064 16541
rect 7472 16575 7524 16584
rect 7472 16541 7481 16575
rect 7481 16541 7515 16575
rect 7515 16541 7524 16575
rect 7472 16532 7524 16541
rect 11060 16600 11112 16652
rect 12532 16643 12584 16652
rect 5632 16464 5684 16516
rect 11704 16575 11756 16584
rect 11704 16541 11713 16575
rect 11713 16541 11747 16575
rect 11747 16541 11756 16575
rect 11704 16532 11756 16541
rect 11888 16532 11940 16584
rect 12532 16609 12541 16643
rect 12541 16609 12575 16643
rect 12575 16609 12584 16643
rect 12532 16600 12584 16609
rect 12164 16532 12216 16584
rect 14648 16779 14700 16788
rect 14648 16745 14657 16779
rect 14657 16745 14691 16779
rect 14691 16745 14700 16779
rect 14648 16736 14700 16745
rect 15292 16736 15344 16788
rect 15660 16736 15712 16788
rect 16764 16736 16816 16788
rect 15108 16668 15160 16720
rect 16212 16668 16264 16720
rect 18052 16668 18104 16720
rect 9772 16439 9824 16448
rect 9772 16405 9781 16439
rect 9781 16405 9815 16439
rect 9815 16405 9824 16439
rect 9772 16396 9824 16405
rect 12348 16464 12400 16516
rect 10876 16396 10928 16448
rect 11244 16396 11296 16448
rect 11980 16396 12032 16448
rect 12716 16507 12768 16516
rect 12716 16473 12725 16507
rect 12725 16473 12759 16507
rect 12759 16473 12768 16507
rect 12716 16464 12768 16473
rect 13176 16464 13228 16516
rect 13544 16464 13596 16516
rect 15384 16532 15436 16584
rect 16028 16600 16080 16652
rect 16580 16532 16632 16584
rect 14740 16507 14792 16516
rect 14740 16473 14749 16507
rect 14749 16473 14783 16507
rect 14783 16473 14792 16507
rect 14740 16464 14792 16473
rect 12992 16396 13044 16448
rect 13084 16439 13136 16448
rect 13084 16405 13093 16439
rect 13093 16405 13127 16439
rect 13127 16405 13136 16439
rect 13084 16396 13136 16405
rect 13360 16439 13412 16448
rect 13360 16405 13369 16439
rect 13369 16405 13403 16439
rect 13403 16405 13412 16439
rect 13360 16396 13412 16405
rect 13452 16396 13504 16448
rect 15108 16507 15160 16516
rect 15108 16473 15117 16507
rect 15117 16473 15151 16507
rect 15151 16473 15160 16507
rect 15108 16464 15160 16473
rect 15568 16464 15620 16516
rect 16672 16464 16724 16516
rect 16764 16464 16816 16516
rect 17500 16532 17552 16584
rect 17776 16575 17828 16584
rect 17776 16541 17785 16575
rect 17785 16541 17819 16575
rect 17819 16541 17828 16575
rect 17776 16532 17828 16541
rect 18328 16575 18380 16584
rect 18328 16541 18337 16575
rect 18337 16541 18371 16575
rect 18371 16541 18380 16575
rect 18328 16532 18380 16541
rect 16304 16396 16356 16448
rect 17224 16439 17276 16448
rect 17224 16405 17233 16439
rect 17233 16405 17267 16439
rect 17267 16405 17276 16439
rect 17224 16396 17276 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 1492 16192 1544 16244
rect 7472 16192 7524 16244
rect 8760 16192 8812 16244
rect 9312 16192 9364 16244
rect 1308 16056 1360 16108
rect 11152 16124 11204 16176
rect 11704 16235 11756 16244
rect 11704 16201 11713 16235
rect 11713 16201 11747 16235
rect 11747 16201 11756 16235
rect 11704 16192 11756 16201
rect 12164 16192 12216 16244
rect 12440 16192 12492 16244
rect 13268 16235 13320 16244
rect 13268 16201 13277 16235
rect 13277 16201 13311 16235
rect 13311 16201 13320 16235
rect 13268 16192 13320 16201
rect 14004 16235 14056 16244
rect 14004 16201 14013 16235
rect 14013 16201 14047 16235
rect 14047 16201 14056 16235
rect 14004 16192 14056 16201
rect 15108 16235 15160 16244
rect 15108 16201 15117 16235
rect 15117 16201 15151 16235
rect 15151 16201 15160 16235
rect 15108 16192 15160 16201
rect 15660 16235 15712 16244
rect 15660 16201 15685 16235
rect 15685 16201 15712 16235
rect 15660 16192 15712 16201
rect 16580 16192 16632 16244
rect 16856 16235 16908 16244
rect 16856 16201 16865 16235
rect 16865 16201 16899 16235
rect 16899 16201 16908 16235
rect 16856 16192 16908 16201
rect 17500 16192 17552 16244
rect 17960 16235 18012 16244
rect 17960 16201 17969 16235
rect 17969 16201 18003 16235
rect 18003 16201 18012 16235
rect 17960 16192 18012 16201
rect 18512 16235 18564 16244
rect 18512 16201 18521 16235
rect 18521 16201 18555 16235
rect 18555 16201 18564 16235
rect 18512 16192 18564 16201
rect 4988 16031 5040 16040
rect 4988 15997 4997 16031
rect 4997 15997 5031 16031
rect 5031 15997 5040 16031
rect 4988 15988 5040 15997
rect 5632 16099 5684 16108
rect 5632 16065 5641 16099
rect 5641 16065 5675 16099
rect 5675 16065 5684 16099
rect 5632 16056 5684 16065
rect 5816 16099 5868 16108
rect 5816 16065 5825 16099
rect 5825 16065 5859 16099
rect 5859 16065 5868 16099
rect 5816 16056 5868 16065
rect 6920 16099 6972 16108
rect 6920 16065 6929 16099
rect 6929 16065 6963 16099
rect 6963 16065 6972 16099
rect 6920 16056 6972 16065
rect 7012 16031 7064 16040
rect 7012 15997 7021 16031
rect 7021 15997 7055 16031
rect 7055 15997 7064 16031
rect 7012 15988 7064 15997
rect 9220 15988 9272 16040
rect 9772 16056 9824 16108
rect 10600 15988 10652 16040
rect 11244 16056 11296 16108
rect 11888 16099 11940 16108
rect 11888 16065 11897 16099
rect 11897 16065 11931 16099
rect 11931 16065 11940 16099
rect 11888 16056 11940 16065
rect 11980 16099 12032 16108
rect 11980 16065 11989 16099
rect 11989 16065 12023 16099
rect 12023 16065 12032 16099
rect 11980 16056 12032 16065
rect 8208 15920 8260 15972
rect 9864 15920 9916 15972
rect 5632 15852 5684 15904
rect 8484 15895 8536 15904
rect 8484 15861 8493 15895
rect 8493 15861 8527 15895
rect 8527 15861 8536 15895
rect 8484 15852 8536 15861
rect 8760 15895 8812 15904
rect 8760 15861 8769 15895
rect 8769 15861 8803 15895
rect 8803 15861 8812 15895
rect 8760 15852 8812 15861
rect 10416 15895 10468 15904
rect 10416 15861 10425 15895
rect 10425 15861 10459 15895
rect 10459 15861 10468 15895
rect 10416 15852 10468 15861
rect 10784 15852 10836 15904
rect 11060 16031 11112 16040
rect 11060 15997 11069 16031
rect 11069 15997 11103 16031
rect 11103 15997 11112 16031
rect 11060 15988 11112 15997
rect 11244 15920 11296 15972
rect 12440 16056 12492 16108
rect 13360 16124 13412 16176
rect 12624 16099 12676 16108
rect 12624 16065 12633 16099
rect 12633 16065 12667 16099
rect 12667 16065 12676 16099
rect 12624 16056 12676 16065
rect 12716 16056 12768 16108
rect 13176 16056 13228 16108
rect 16028 16124 16080 16176
rect 16304 16124 16356 16176
rect 13912 16056 13964 16108
rect 14556 16056 14608 16108
rect 16488 16056 16540 16108
rect 15936 15988 15988 16040
rect 17224 15988 17276 16040
rect 13084 15920 13136 15972
rect 12808 15895 12860 15904
rect 12808 15861 12817 15895
rect 12817 15861 12851 15895
rect 12851 15861 12860 15895
rect 12808 15852 12860 15861
rect 13728 15895 13780 15904
rect 13728 15861 13737 15895
rect 13737 15861 13771 15895
rect 13771 15861 13780 15895
rect 13728 15852 13780 15861
rect 15752 15920 15804 15972
rect 16580 15920 16632 15972
rect 16028 15852 16080 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 9312 15580 9364 15632
rect 4988 15555 5040 15564
rect 4988 15521 4997 15555
rect 4997 15521 5031 15555
rect 5031 15521 5040 15555
rect 4988 15512 5040 15521
rect 6736 15555 6788 15564
rect 6736 15521 6745 15555
rect 6745 15521 6779 15555
rect 6779 15521 6788 15555
rect 6736 15512 6788 15521
rect 9772 15580 9824 15632
rect 11244 15691 11296 15700
rect 11244 15657 11253 15691
rect 11253 15657 11287 15691
rect 11287 15657 11296 15691
rect 11244 15648 11296 15657
rect 12992 15648 13044 15700
rect 13728 15648 13780 15700
rect 11888 15580 11940 15632
rect 5264 15487 5316 15496
rect 5264 15453 5273 15487
rect 5273 15453 5307 15487
rect 5307 15453 5316 15487
rect 5264 15444 5316 15453
rect 5632 15487 5684 15496
rect 5632 15453 5641 15487
rect 5641 15453 5675 15487
rect 5675 15453 5684 15487
rect 5632 15444 5684 15453
rect 6552 15444 6604 15496
rect 6460 15376 6512 15428
rect 8852 15376 8904 15428
rect 9680 15487 9732 15496
rect 9680 15453 9689 15487
rect 9689 15453 9723 15487
rect 9723 15453 9732 15487
rect 9680 15444 9732 15453
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 9772 15444 9824 15453
rect 9956 15444 10008 15496
rect 10416 15444 10468 15496
rect 10784 15487 10836 15496
rect 10784 15453 10791 15487
rect 10791 15453 10836 15487
rect 10784 15444 10836 15453
rect 11980 15512 12032 15564
rect 13452 15580 13504 15632
rect 13820 15623 13872 15632
rect 13820 15589 13829 15623
rect 13829 15589 13863 15623
rect 13863 15589 13872 15623
rect 13820 15580 13872 15589
rect 12624 15512 12676 15564
rect 15200 15512 15252 15564
rect 15660 15512 15712 15564
rect 12440 15444 12492 15496
rect 13084 15487 13136 15496
rect 13084 15453 13093 15487
rect 13093 15453 13127 15487
rect 13127 15453 13136 15487
rect 13084 15444 13136 15453
rect 10508 15376 10560 15428
rect 8484 15351 8536 15360
rect 8484 15317 8493 15351
rect 8493 15317 8527 15351
rect 8527 15317 8536 15351
rect 8484 15308 8536 15317
rect 8576 15351 8628 15360
rect 8576 15317 8585 15351
rect 8585 15317 8619 15351
rect 8619 15317 8628 15351
rect 8576 15308 8628 15317
rect 8668 15308 8720 15360
rect 10784 15308 10836 15360
rect 10968 15419 11020 15428
rect 10968 15385 10977 15419
rect 10977 15385 11011 15419
rect 11011 15385 11020 15419
rect 10968 15376 11020 15385
rect 12532 15376 12584 15428
rect 13360 15419 13412 15428
rect 13360 15385 13369 15419
rect 13369 15385 13403 15419
rect 13403 15385 13412 15419
rect 13360 15376 13412 15385
rect 14464 15487 14516 15496
rect 14464 15453 14473 15487
rect 14473 15453 14507 15487
rect 14507 15453 14516 15487
rect 14464 15444 14516 15453
rect 15384 15487 15436 15496
rect 15384 15453 15393 15487
rect 15393 15453 15427 15487
rect 15427 15453 15436 15487
rect 15384 15444 15436 15453
rect 15568 15487 15620 15496
rect 15568 15453 15577 15487
rect 15577 15453 15611 15487
rect 15611 15453 15620 15487
rect 15568 15444 15620 15453
rect 16028 15512 16080 15564
rect 16120 15487 16172 15496
rect 16120 15453 16129 15487
rect 16129 15453 16163 15487
rect 16163 15453 16172 15487
rect 16120 15444 16172 15453
rect 16580 15444 16632 15496
rect 11428 15308 11480 15360
rect 12992 15308 13044 15360
rect 17132 15351 17184 15360
rect 17132 15317 17141 15351
rect 17141 15317 17175 15351
rect 17175 15317 17184 15351
rect 17132 15308 17184 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 1308 14968 1360 15020
rect 6736 15104 6788 15156
rect 9772 15104 9824 15156
rect 12808 15104 12860 15156
rect 4068 14968 4120 15020
rect 5540 15036 5592 15088
rect 4804 14968 4856 15020
rect 6736 14968 6788 15020
rect 8484 14968 8536 15020
rect 8852 15036 8904 15088
rect 15292 15036 15344 15088
rect 9312 14968 9364 15020
rect 12900 14968 12952 15020
rect 13452 15011 13504 15020
rect 13452 14977 13461 15011
rect 13461 14977 13495 15011
rect 13495 14977 13504 15011
rect 13452 14968 13504 14977
rect 13820 14968 13872 15020
rect 15384 14968 15436 15020
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 15660 14968 15712 14977
rect 16120 15036 16172 15088
rect 5264 14900 5316 14952
rect 6460 14900 6512 14952
rect 5448 14832 5500 14884
rect 8576 14900 8628 14952
rect 9956 14900 10008 14952
rect 15568 14943 15620 14952
rect 15568 14909 15577 14943
rect 15577 14909 15611 14943
rect 15611 14909 15620 14943
rect 15568 14900 15620 14909
rect 8392 14832 8444 14884
rect 8760 14832 8812 14884
rect 12348 14764 12400 14816
rect 15292 14807 15344 14816
rect 15292 14773 15301 14807
rect 15301 14773 15335 14807
rect 15335 14773 15344 14807
rect 15292 14764 15344 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 4068 14424 4120 14476
rect 4528 14467 4580 14476
rect 4528 14433 4537 14467
rect 4537 14433 4571 14467
rect 4571 14433 4580 14467
rect 4528 14424 4580 14433
rect 6460 14467 6512 14476
rect 6460 14433 6469 14467
rect 6469 14433 6503 14467
rect 6503 14433 6512 14467
rect 6460 14424 6512 14433
rect 5540 14356 5592 14408
rect 6736 14356 6788 14408
rect 9956 14560 10008 14612
rect 13084 14560 13136 14612
rect 9772 14492 9824 14544
rect 10600 14535 10652 14544
rect 10600 14501 10609 14535
rect 10609 14501 10643 14535
rect 10643 14501 10652 14535
rect 10600 14492 10652 14501
rect 11520 14492 11572 14544
rect 12624 14492 12676 14544
rect 9220 14424 9272 14476
rect 9680 14356 9732 14408
rect 9956 14356 10008 14408
rect 11612 14424 11664 14476
rect 10416 14399 10468 14408
rect 10416 14365 10425 14399
rect 10425 14365 10459 14399
rect 10459 14365 10468 14399
rect 10416 14356 10468 14365
rect 11336 14356 11388 14408
rect 17500 14424 17552 14476
rect 12624 14356 12676 14408
rect 12992 14356 13044 14408
rect 13636 14356 13688 14408
rect 16396 14399 16448 14408
rect 16396 14365 16405 14399
rect 16405 14365 16439 14399
rect 16439 14365 16448 14399
rect 16396 14356 16448 14365
rect 6920 14263 6972 14272
rect 6920 14229 6929 14263
rect 6929 14229 6963 14263
rect 6963 14229 6972 14263
rect 6920 14220 6972 14229
rect 8944 14263 8996 14272
rect 8944 14229 8953 14263
rect 8953 14229 8987 14263
rect 8987 14229 8996 14263
rect 8944 14220 8996 14229
rect 9496 14220 9548 14272
rect 11060 14220 11112 14272
rect 14188 14331 14240 14340
rect 14188 14297 14197 14331
rect 14197 14297 14231 14331
rect 14231 14297 14240 14331
rect 14188 14288 14240 14297
rect 14372 14331 14424 14340
rect 14372 14297 14381 14331
rect 14381 14297 14415 14331
rect 14415 14297 14424 14331
rect 14372 14288 14424 14297
rect 16212 14288 16264 14340
rect 12348 14263 12400 14272
rect 12348 14229 12357 14263
rect 12357 14229 12391 14263
rect 12391 14229 12400 14263
rect 12348 14220 12400 14229
rect 12532 14263 12584 14272
rect 12532 14229 12541 14263
rect 12541 14229 12575 14263
rect 12575 14229 12584 14263
rect 12532 14220 12584 14229
rect 16948 14220 17000 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 5724 14016 5776 14068
rect 4528 13991 4580 14000
rect 4528 13957 4537 13991
rect 4537 13957 4571 13991
rect 4571 13957 4580 13991
rect 4528 13948 4580 13957
rect 6920 13991 6972 14000
rect 6920 13957 6929 13991
rect 6929 13957 6963 13991
rect 6963 13957 6972 13991
rect 6920 13948 6972 13957
rect 8300 13948 8352 14000
rect 9680 14016 9732 14068
rect 10416 14016 10468 14068
rect 12440 14016 12492 14068
rect 16948 14059 17000 14068
rect 16948 14025 16957 14059
rect 16957 14025 16991 14059
rect 16991 14025 17000 14059
rect 16948 14016 17000 14025
rect 17684 14016 17736 14068
rect 1308 13880 1360 13932
rect 4896 13787 4948 13796
rect 4896 13753 4905 13787
rect 4905 13753 4939 13787
rect 4939 13753 4948 13787
rect 5908 13880 5960 13932
rect 6828 13923 6880 13932
rect 6828 13889 6837 13923
rect 6837 13889 6871 13923
rect 6871 13889 6880 13923
rect 6828 13880 6880 13889
rect 7196 13880 7248 13932
rect 9496 13948 9548 14000
rect 8852 13923 8904 13932
rect 8852 13889 8861 13923
rect 8861 13889 8895 13923
rect 8895 13889 8904 13923
rect 8852 13880 8904 13889
rect 11060 13923 11112 13932
rect 11060 13889 11069 13923
rect 11069 13889 11103 13923
rect 11103 13889 11112 13923
rect 11060 13880 11112 13889
rect 11520 13923 11572 13932
rect 11520 13889 11529 13923
rect 11529 13889 11563 13923
rect 11563 13889 11572 13923
rect 11520 13880 11572 13889
rect 11612 13923 11664 13932
rect 11612 13889 11621 13923
rect 11621 13889 11655 13923
rect 11655 13889 11664 13923
rect 11612 13880 11664 13889
rect 4896 13744 4948 13753
rect 1584 13719 1636 13728
rect 1584 13685 1593 13719
rect 1593 13685 1627 13719
rect 1627 13685 1636 13719
rect 1584 13676 1636 13685
rect 8668 13812 8720 13864
rect 10968 13855 11020 13864
rect 10968 13821 10977 13855
rect 10977 13821 11011 13855
rect 11011 13821 11020 13855
rect 10968 13812 11020 13821
rect 12532 13880 12584 13932
rect 15752 13948 15804 14000
rect 12992 13923 13044 13932
rect 12992 13889 13001 13923
rect 13001 13889 13035 13923
rect 13035 13889 13044 13923
rect 12992 13880 13044 13889
rect 13636 13923 13688 13932
rect 13636 13889 13645 13923
rect 13645 13889 13679 13923
rect 13679 13889 13688 13923
rect 13636 13880 13688 13889
rect 14464 13923 14516 13932
rect 14464 13889 14473 13923
rect 14473 13889 14507 13923
rect 14507 13889 14516 13923
rect 14464 13880 14516 13889
rect 15292 13880 15344 13932
rect 16028 13923 16080 13932
rect 16028 13889 16037 13923
rect 16037 13889 16071 13923
rect 16071 13889 16080 13923
rect 16028 13880 16080 13889
rect 16396 13948 16448 14000
rect 16212 13923 16264 13932
rect 16212 13889 16221 13923
rect 16221 13889 16255 13923
rect 16255 13889 16264 13923
rect 16212 13880 16264 13889
rect 17040 13923 17092 13932
rect 17040 13889 17049 13923
rect 17049 13889 17083 13923
rect 17083 13889 17092 13923
rect 17040 13880 17092 13889
rect 12256 13812 12308 13864
rect 12440 13855 12492 13864
rect 12440 13821 12449 13855
rect 12449 13821 12483 13855
rect 12483 13821 12492 13855
rect 12440 13812 12492 13821
rect 11612 13744 11664 13796
rect 12716 13812 12768 13864
rect 14372 13855 14424 13864
rect 14372 13821 14381 13855
rect 14381 13821 14415 13855
rect 14415 13821 14424 13855
rect 14372 13812 14424 13821
rect 5632 13676 5684 13728
rect 5816 13719 5868 13728
rect 5816 13685 5825 13719
rect 5825 13685 5859 13719
rect 5859 13685 5868 13719
rect 5816 13676 5868 13685
rect 10968 13676 11020 13728
rect 12624 13744 12676 13796
rect 14280 13744 14332 13796
rect 16488 13855 16540 13864
rect 16488 13821 16497 13855
rect 16497 13821 16531 13855
rect 16531 13821 16540 13855
rect 16488 13812 16540 13821
rect 14004 13676 14056 13728
rect 16580 13744 16632 13796
rect 17316 13744 17368 13796
rect 17776 13744 17828 13796
rect 17868 13676 17920 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 4896 13472 4948 13524
rect 5908 13515 5960 13524
rect 5908 13481 5917 13515
rect 5917 13481 5951 13515
rect 5951 13481 5960 13515
rect 5908 13472 5960 13481
rect 6828 13472 6880 13524
rect 14188 13472 14240 13524
rect 14280 13515 14332 13524
rect 14280 13481 14289 13515
rect 14289 13481 14323 13515
rect 14323 13481 14332 13515
rect 14280 13472 14332 13481
rect 14372 13472 14424 13524
rect 8668 13447 8720 13456
rect 8668 13413 8677 13447
rect 8677 13413 8711 13447
rect 8711 13413 8720 13447
rect 8668 13404 8720 13413
rect 8944 13404 8996 13456
rect 9404 13404 9456 13456
rect 15660 13472 15712 13524
rect 17040 13472 17092 13524
rect 4068 13379 4120 13388
rect 4068 13345 4077 13379
rect 4077 13345 4111 13379
rect 4111 13345 4120 13379
rect 4068 13336 4120 13345
rect 12900 13336 12952 13388
rect 12992 13379 13044 13388
rect 12992 13345 13001 13379
rect 13001 13345 13035 13379
rect 13035 13345 13044 13379
rect 12992 13336 13044 13345
rect 4804 13268 4856 13320
rect 5448 13311 5500 13320
rect 5448 13277 5457 13311
rect 5457 13277 5491 13311
rect 5491 13277 5500 13311
rect 5448 13268 5500 13277
rect 5724 13311 5776 13320
rect 5724 13277 5733 13311
rect 5733 13277 5767 13311
rect 5767 13277 5776 13311
rect 5724 13268 5776 13277
rect 8392 13311 8444 13320
rect 8392 13277 8401 13311
rect 8401 13277 8435 13311
rect 8435 13277 8444 13311
rect 8392 13268 8444 13277
rect 8576 13268 8628 13320
rect 13360 13268 13412 13320
rect 15476 13404 15528 13456
rect 16028 13404 16080 13456
rect 16212 13404 16264 13456
rect 14004 13336 14056 13388
rect 18052 13336 18104 13388
rect 5540 13175 5592 13184
rect 5540 13141 5549 13175
rect 5549 13141 5583 13175
rect 5583 13141 5592 13175
rect 5540 13132 5592 13141
rect 8484 13175 8536 13184
rect 8484 13141 8493 13175
rect 8493 13141 8527 13175
rect 8527 13141 8536 13175
rect 8484 13132 8536 13141
rect 14188 13200 14240 13252
rect 15292 13268 15344 13320
rect 14556 13200 14608 13252
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 15660 13311 15712 13320
rect 15660 13277 15669 13311
rect 15669 13277 15703 13311
rect 15703 13277 15712 13311
rect 15660 13268 15712 13277
rect 15752 13311 15804 13320
rect 15752 13277 15761 13311
rect 15761 13277 15795 13311
rect 15795 13277 15804 13311
rect 15752 13268 15804 13277
rect 16028 13268 16080 13320
rect 8760 13132 8812 13184
rect 11336 13132 11388 13184
rect 15200 13175 15252 13184
rect 15200 13141 15209 13175
rect 15209 13141 15243 13175
rect 15243 13141 15252 13175
rect 15200 13132 15252 13141
rect 17868 13311 17920 13320
rect 17868 13277 17877 13311
rect 17877 13277 17911 13311
rect 17911 13277 17920 13311
rect 17868 13268 17920 13277
rect 17592 13175 17644 13184
rect 17592 13141 17601 13175
rect 17601 13141 17635 13175
rect 17635 13141 17644 13175
rect 17592 13132 17644 13141
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 8300 12928 8352 12980
rect 8852 12928 8904 12980
rect 14924 12928 14976 12980
rect 15384 12928 15436 12980
rect 1308 12792 1360 12844
rect 5448 12792 5500 12844
rect 9128 12860 9180 12912
rect 8300 12792 8352 12844
rect 8852 12835 8904 12844
rect 8852 12801 8875 12835
rect 8875 12801 8904 12835
rect 8852 12792 8904 12801
rect 8944 12801 8950 12828
rect 8950 12801 8984 12828
rect 8984 12801 8996 12828
rect 8944 12776 8996 12801
rect 8668 12724 8720 12776
rect 10876 12835 10928 12844
rect 10876 12801 10885 12835
rect 10885 12801 10919 12835
rect 10919 12801 10928 12835
rect 10876 12792 10928 12801
rect 12992 12860 13044 12912
rect 14372 12860 14424 12912
rect 15568 12860 15620 12912
rect 15936 12860 15988 12912
rect 11152 12792 11204 12844
rect 14924 12835 14976 12844
rect 14924 12801 14933 12835
rect 14933 12801 14967 12835
rect 14967 12801 14976 12835
rect 14924 12792 14976 12801
rect 6092 12631 6144 12640
rect 6092 12597 6101 12631
rect 6101 12597 6135 12631
rect 6135 12597 6144 12631
rect 6092 12588 6144 12597
rect 9312 12656 9364 12708
rect 10324 12588 10376 12640
rect 11336 12724 11388 12776
rect 15384 12792 15436 12844
rect 18144 12792 18196 12844
rect 18328 12767 18380 12776
rect 18328 12733 18337 12767
rect 18337 12733 18371 12767
rect 18371 12733 18380 12767
rect 18328 12724 18380 12733
rect 12256 12588 12308 12640
rect 13636 12588 13688 12640
rect 15660 12588 15712 12640
rect 15752 12631 15804 12640
rect 15752 12597 15761 12631
rect 15761 12597 15795 12631
rect 15795 12597 15804 12631
rect 15752 12588 15804 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 6736 12384 6788 12436
rect 8484 12384 8536 12436
rect 8668 12384 8720 12436
rect 10876 12384 10928 12436
rect 13268 12384 13320 12436
rect 13636 12384 13688 12436
rect 4068 12316 4120 12368
rect 5080 12316 5132 12368
rect 4436 12291 4488 12300
rect 4436 12257 4445 12291
rect 4445 12257 4479 12291
rect 4479 12257 4488 12291
rect 4436 12248 4488 12257
rect 5632 12248 5684 12300
rect 6000 12291 6052 12300
rect 6000 12257 6009 12291
rect 6009 12257 6043 12291
rect 6043 12257 6052 12291
rect 6000 12248 6052 12257
rect 6092 12291 6144 12300
rect 6092 12257 6101 12291
rect 6101 12257 6135 12291
rect 6135 12257 6144 12291
rect 6092 12248 6144 12257
rect 8300 12316 8352 12368
rect 8852 12316 8904 12368
rect 8668 12248 8720 12300
rect 9312 12291 9364 12300
rect 9312 12257 9321 12291
rect 9321 12257 9355 12291
rect 9355 12257 9364 12291
rect 9312 12248 9364 12257
rect 3792 12180 3844 12232
rect 4252 12112 4304 12164
rect 5540 12112 5592 12164
rect 8760 12155 8812 12164
rect 8760 12121 8769 12155
rect 8769 12121 8803 12155
rect 8803 12121 8812 12155
rect 8760 12112 8812 12121
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 9404 12223 9456 12232
rect 9404 12189 9413 12223
rect 9413 12189 9447 12223
rect 9447 12189 9456 12223
rect 9404 12180 9456 12189
rect 14004 12316 14056 12368
rect 14924 12248 14976 12300
rect 16488 12248 16540 12300
rect 12532 12180 12584 12232
rect 14372 12180 14424 12232
rect 17132 12223 17184 12232
rect 17132 12189 17141 12223
rect 17141 12189 17175 12223
rect 17175 12189 17184 12223
rect 17132 12180 17184 12189
rect 17592 12180 17644 12232
rect 12256 12155 12308 12164
rect 12256 12121 12265 12155
rect 12265 12121 12299 12155
rect 12299 12121 12308 12155
rect 12256 12112 12308 12121
rect 4988 12087 5040 12096
rect 4988 12053 4997 12087
rect 4997 12053 5031 12087
rect 5031 12053 5040 12087
rect 4988 12044 5040 12053
rect 5080 12087 5132 12096
rect 5080 12053 5089 12087
rect 5089 12053 5123 12087
rect 5123 12053 5132 12087
rect 5080 12044 5132 12053
rect 6552 12087 6604 12096
rect 6552 12053 6561 12087
rect 6561 12053 6595 12087
rect 6595 12053 6604 12087
rect 6552 12044 6604 12053
rect 7196 12087 7248 12096
rect 7196 12053 7205 12087
rect 7205 12053 7239 12087
rect 7239 12053 7248 12087
rect 7196 12044 7248 12053
rect 8576 12087 8628 12096
rect 8576 12053 8603 12087
rect 8603 12053 8628 12087
rect 8576 12044 8628 12053
rect 8944 12087 8996 12096
rect 8944 12053 8953 12087
rect 8953 12053 8987 12087
rect 8987 12053 8996 12087
rect 8944 12044 8996 12053
rect 9496 12087 9548 12096
rect 9496 12053 9505 12087
rect 9505 12053 9539 12087
rect 9539 12053 9548 12087
rect 9496 12044 9548 12053
rect 11612 12087 11664 12096
rect 11612 12053 11621 12087
rect 11621 12053 11655 12087
rect 11655 12053 11664 12087
rect 11612 12044 11664 12053
rect 12992 12044 13044 12096
rect 13268 12112 13320 12164
rect 15384 12112 15436 12164
rect 13360 12087 13412 12096
rect 13360 12053 13385 12087
rect 13385 12053 13412 12087
rect 13360 12044 13412 12053
rect 15292 12044 15344 12096
rect 17776 12044 17828 12096
rect 17868 12044 17920 12096
rect 18236 12044 18288 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 4252 11883 4304 11892
rect 4252 11849 4261 11883
rect 4261 11849 4295 11883
rect 4295 11849 4304 11883
rect 4252 11840 4304 11849
rect 4436 11883 4488 11892
rect 4436 11849 4445 11883
rect 4445 11849 4479 11883
rect 4479 11849 4488 11883
rect 4436 11840 4488 11849
rect 8944 11840 8996 11892
rect 12532 11840 12584 11892
rect 13360 11840 13412 11892
rect 1308 11704 1360 11756
rect 4804 11772 4856 11824
rect 3792 11679 3844 11688
rect 3792 11645 3801 11679
rect 3801 11645 3835 11679
rect 3835 11645 3844 11679
rect 3792 11636 3844 11645
rect 3976 11636 4028 11688
rect 6736 11704 6788 11756
rect 9496 11772 9548 11824
rect 8576 11636 8628 11688
rect 8760 11679 8812 11688
rect 8760 11645 8769 11679
rect 8769 11645 8803 11679
rect 8803 11645 8812 11679
rect 8760 11636 8812 11645
rect 9220 11636 9272 11688
rect 9680 11679 9732 11688
rect 9680 11645 9689 11679
rect 9689 11645 9723 11679
rect 9723 11645 9732 11679
rect 9680 11636 9732 11645
rect 9312 11568 9364 11620
rect 10324 11747 10376 11756
rect 10324 11713 10333 11747
rect 10333 11713 10367 11747
rect 10367 11713 10376 11747
rect 10324 11704 10376 11713
rect 11612 11772 11664 11824
rect 10692 11704 10744 11756
rect 14004 11747 14056 11756
rect 14004 11713 14013 11747
rect 14013 11713 14047 11747
rect 14047 11713 14056 11747
rect 14004 11704 14056 11713
rect 14188 11747 14240 11756
rect 14188 11713 14197 11747
rect 14197 11713 14231 11747
rect 14231 11713 14240 11747
rect 14188 11704 14240 11713
rect 15200 11840 15252 11892
rect 15292 11840 15344 11892
rect 10508 11679 10560 11688
rect 10508 11645 10517 11679
rect 10517 11645 10551 11679
rect 10551 11645 10560 11679
rect 10508 11636 10560 11645
rect 15292 11747 15344 11756
rect 15292 11713 15301 11747
rect 15301 11713 15335 11747
rect 15335 11713 15344 11747
rect 15292 11704 15344 11713
rect 15384 11747 15436 11756
rect 15384 11713 15393 11747
rect 15393 11713 15427 11747
rect 15427 11713 15436 11747
rect 15384 11704 15436 11713
rect 15660 11747 15712 11756
rect 15660 11713 15669 11747
rect 15669 11713 15703 11747
rect 15703 11713 15712 11747
rect 15660 11704 15712 11713
rect 15752 11747 15804 11756
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 17132 11840 17184 11892
rect 17868 11840 17920 11892
rect 17960 11772 18012 11824
rect 16396 11747 16448 11756
rect 16396 11713 16399 11747
rect 16399 11713 16433 11747
rect 16433 11713 16448 11747
rect 14832 11636 14884 11688
rect 16396 11704 16448 11713
rect 11796 11568 11848 11620
rect 14648 11611 14700 11620
rect 14648 11577 14657 11611
rect 14657 11577 14691 11611
rect 14691 11577 14700 11611
rect 14648 11568 14700 11577
rect 17776 11704 17828 11756
rect 18236 11747 18288 11756
rect 18236 11713 18245 11747
rect 18245 11713 18279 11747
rect 18279 11713 18288 11747
rect 18236 11704 18288 11713
rect 16856 11679 16908 11688
rect 16856 11645 16865 11679
rect 16865 11645 16899 11679
rect 16899 11645 16908 11679
rect 16856 11636 16908 11645
rect 17408 11636 17460 11688
rect 16948 11568 17000 11620
rect 7288 11500 7340 11552
rect 7656 11500 7708 11552
rect 15384 11500 15436 11552
rect 16396 11500 16448 11552
rect 17224 11500 17276 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 5816 11296 5868 11348
rect 14648 11296 14700 11348
rect 14832 11339 14884 11348
rect 14832 11305 14841 11339
rect 14841 11305 14875 11339
rect 14875 11305 14884 11339
rect 14832 11296 14884 11305
rect 6000 11228 6052 11280
rect 7288 11203 7340 11212
rect 7288 11169 7297 11203
rect 7297 11169 7331 11203
rect 7331 11169 7340 11203
rect 7288 11160 7340 11169
rect 8760 11160 8812 11212
rect 9312 11160 9364 11212
rect 10508 11160 10560 11212
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 1584 11024 1636 11076
rect 9680 11092 9732 11144
rect 13452 11067 13504 11076
rect 13452 11033 13461 11067
rect 13461 11033 13495 11067
rect 13495 11033 13504 11067
rect 13452 11024 13504 11033
rect 14004 11024 14056 11076
rect 14188 11092 14240 11144
rect 15660 11228 15712 11280
rect 16856 11228 16908 11280
rect 15752 11160 15804 11212
rect 18052 11203 18104 11212
rect 18052 11169 18061 11203
rect 18061 11169 18095 11203
rect 18095 11169 18104 11203
rect 18052 11160 18104 11169
rect 18144 11203 18196 11212
rect 18144 11169 18153 11203
rect 18153 11169 18187 11203
rect 18187 11169 18196 11203
rect 18144 11160 18196 11169
rect 15292 11135 15344 11144
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 15384 11135 15436 11144
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 17868 11092 17920 11144
rect 15200 11024 15252 11076
rect 8208 10956 8260 11008
rect 12808 10956 12860 11008
rect 17592 10999 17644 11008
rect 17592 10965 17601 10999
rect 17601 10965 17635 10999
rect 17635 10965 17644 10999
rect 17592 10956 17644 10965
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 3976 10752 4028 10804
rect 10508 10752 10560 10804
rect 1308 10616 1360 10668
rect 5908 10684 5960 10736
rect 9680 10684 9732 10736
rect 10692 10684 10744 10736
rect 5356 10591 5408 10600
rect 5356 10557 5365 10591
rect 5365 10557 5399 10591
rect 5399 10557 5408 10591
rect 5356 10548 5408 10557
rect 8392 10480 8444 10532
rect 6828 10412 6880 10464
rect 10324 10616 10376 10668
rect 13452 10752 13504 10804
rect 17316 10752 17368 10804
rect 10692 10548 10744 10600
rect 12808 10659 12860 10668
rect 12808 10625 12817 10659
rect 12817 10625 12851 10659
rect 12851 10625 12860 10659
rect 12808 10616 12860 10625
rect 12992 10616 13044 10668
rect 13176 10659 13228 10668
rect 13176 10625 13185 10659
rect 13185 10625 13219 10659
rect 13219 10625 13228 10659
rect 13176 10616 13228 10625
rect 14004 10616 14056 10668
rect 16764 10616 16816 10668
rect 16948 10659 17000 10668
rect 16948 10625 16957 10659
rect 16957 10625 16991 10659
rect 16991 10625 17000 10659
rect 16948 10616 17000 10625
rect 11980 10548 12032 10600
rect 15752 10548 15804 10600
rect 16856 10548 16908 10600
rect 9036 10412 9088 10464
rect 11152 10412 11204 10464
rect 13176 10480 13228 10532
rect 16580 10480 16632 10532
rect 17132 10480 17184 10532
rect 12532 10455 12584 10464
rect 12532 10421 12541 10455
rect 12541 10421 12575 10455
rect 12575 10421 12584 10455
rect 12532 10412 12584 10421
rect 15292 10412 15344 10464
rect 18144 10412 18196 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 4620 10251 4672 10260
rect 4620 10217 4629 10251
rect 4629 10217 4663 10251
rect 4663 10217 4672 10251
rect 4620 10208 4672 10217
rect 5356 10208 5408 10260
rect 4896 10140 4948 10192
rect 1308 10004 1360 10056
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 4620 9911 4672 9920
rect 4620 9877 4645 9911
rect 4645 9877 4672 9911
rect 6184 10004 6236 10056
rect 8392 10208 8444 10260
rect 12992 10251 13044 10260
rect 12992 10217 13001 10251
rect 13001 10217 13035 10251
rect 13035 10217 13044 10251
rect 12992 10208 13044 10217
rect 13176 10208 13228 10260
rect 6828 10140 6880 10192
rect 6920 10072 6972 10124
rect 12532 10140 12584 10192
rect 15568 10140 15620 10192
rect 16672 10140 16724 10192
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 10232 10004 10284 10056
rect 15200 10115 15252 10124
rect 15200 10081 15209 10115
rect 15209 10081 15243 10115
rect 15243 10081 15252 10115
rect 15200 10072 15252 10081
rect 16948 10072 17000 10124
rect 4620 9868 4672 9877
rect 4988 9911 5040 9920
rect 4988 9877 4997 9911
rect 4997 9877 5031 9911
rect 5031 9877 5040 9911
rect 4988 9868 5040 9877
rect 5540 9936 5592 9988
rect 6092 9936 6144 9988
rect 8300 9936 8352 9988
rect 9588 9936 9640 9988
rect 5264 9868 5316 9920
rect 5632 9868 5684 9920
rect 6000 9911 6052 9920
rect 6000 9877 6009 9911
rect 6009 9877 6043 9911
rect 6043 9877 6052 9911
rect 6000 9868 6052 9877
rect 6276 9911 6328 9920
rect 6276 9877 6285 9911
rect 6285 9877 6319 9911
rect 6319 9877 6328 9911
rect 6276 9868 6328 9877
rect 7932 9868 7984 9920
rect 8024 9868 8076 9920
rect 11980 9936 12032 9988
rect 15292 10047 15344 10056
rect 15292 10013 15301 10047
rect 15301 10013 15335 10047
rect 15335 10013 15344 10047
rect 15292 10004 15344 10013
rect 15752 10047 15804 10056
rect 15752 10013 15761 10047
rect 15761 10013 15795 10047
rect 15795 10013 15804 10047
rect 15752 10004 15804 10013
rect 16580 10004 16632 10056
rect 16856 10047 16908 10056
rect 16856 10013 16865 10047
rect 16865 10013 16899 10047
rect 16899 10013 16908 10047
rect 16856 10004 16908 10013
rect 13544 9868 13596 9920
rect 16212 9868 16264 9920
rect 16764 9936 16816 9988
rect 16948 9936 17000 9988
rect 17408 10004 17460 10056
rect 18144 9936 18196 9988
rect 17960 9911 18012 9920
rect 17960 9877 17969 9911
rect 17969 9877 18003 9911
rect 18003 9877 18012 9911
rect 17960 9868 18012 9877
rect 18512 9868 18564 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 2688 9596 2740 9648
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 1584 9528 1636 9537
rect 1676 9571 1728 9580
rect 1676 9537 1685 9571
rect 1685 9537 1719 9571
rect 1719 9537 1728 9571
rect 1676 9528 1728 9537
rect 2136 9571 2188 9580
rect 2136 9537 2139 9571
rect 2139 9537 2188 9571
rect 2136 9528 2188 9537
rect 2320 9571 2372 9580
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 5540 9664 5592 9716
rect 5632 9664 5684 9716
rect 9220 9664 9272 9716
rect 16856 9664 16908 9716
rect 8392 9596 8444 9648
rect 16764 9596 16816 9648
rect 2872 9528 2924 9580
rect 3424 9571 3476 9580
rect 3424 9537 3433 9571
rect 3433 9537 3467 9571
rect 3467 9537 3476 9571
rect 3424 9528 3476 9537
rect 5448 9460 5500 9512
rect 6000 9528 6052 9580
rect 6184 9571 6236 9580
rect 6184 9537 6193 9571
rect 6193 9537 6227 9571
rect 6227 9537 6236 9571
rect 6184 9528 6236 9537
rect 6276 9528 6328 9580
rect 6644 9571 6696 9580
rect 6644 9537 6653 9571
rect 6653 9537 6687 9571
rect 6687 9537 6696 9571
rect 6644 9528 6696 9537
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 8024 9571 8076 9580
rect 8024 9537 8033 9571
rect 8033 9537 8067 9571
rect 8067 9537 8076 9571
rect 8024 9528 8076 9537
rect 9588 9528 9640 9580
rect 11888 9528 11940 9580
rect 16856 9571 16908 9580
rect 16856 9537 16865 9571
rect 16865 9537 16899 9571
rect 16899 9537 16908 9571
rect 16856 9528 16908 9537
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 4896 9324 4948 9376
rect 5264 9324 5316 9376
rect 8300 9435 8352 9444
rect 8300 9401 8309 9435
rect 8309 9401 8343 9435
rect 8343 9401 8352 9435
rect 8300 9392 8352 9401
rect 17132 9528 17184 9580
rect 17960 9392 18012 9444
rect 10784 9324 10836 9376
rect 12348 9367 12400 9376
rect 12348 9333 12357 9367
rect 12357 9333 12391 9367
rect 12391 9333 12400 9367
rect 12348 9324 12400 9333
rect 17500 9324 17552 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 2320 9120 2372 9172
rect 4620 9120 4672 9172
rect 4896 9120 4948 9172
rect 3516 9052 3568 9104
rect 1676 9027 1728 9036
rect 1676 8993 1685 9027
rect 1685 8993 1719 9027
rect 1719 8993 1728 9027
rect 1676 8984 1728 8993
rect 4712 9052 4764 9104
rect 9128 9052 9180 9104
rect 9404 9163 9456 9172
rect 9404 9129 9413 9163
rect 9413 9129 9447 9163
rect 9447 9129 9456 9163
rect 9404 9120 9456 9129
rect 9956 9120 10008 9172
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 3516 8916 3568 8968
rect 5356 8916 5408 8968
rect 3792 8891 3844 8900
rect 3792 8857 3801 8891
rect 3801 8857 3835 8891
rect 3835 8857 3844 8891
rect 3792 8848 3844 8857
rect 4620 8891 4672 8900
rect 4620 8857 4629 8891
rect 4629 8857 4663 8891
rect 4663 8857 4672 8891
rect 4620 8848 4672 8857
rect 4712 8848 4764 8900
rect 5632 8891 5684 8900
rect 5632 8857 5641 8891
rect 5641 8857 5675 8891
rect 5675 8857 5684 8891
rect 5632 8848 5684 8857
rect 6184 9027 6236 9036
rect 6184 8993 6193 9027
rect 6193 8993 6227 9027
rect 6227 8993 6236 9027
rect 6184 8984 6236 8993
rect 6644 9027 6696 9036
rect 6644 8993 6653 9027
rect 6653 8993 6687 9027
rect 6687 8993 6696 9027
rect 6644 8984 6696 8993
rect 8024 9027 8076 9036
rect 8024 8993 8033 9027
rect 8033 8993 8067 9027
rect 8067 8993 8076 9027
rect 8024 8984 8076 8993
rect 12440 9163 12492 9172
rect 12440 9129 12449 9163
rect 12449 9129 12483 9163
rect 12483 9129 12492 9163
rect 12440 9120 12492 9129
rect 13820 9120 13872 9172
rect 10048 8984 10100 9036
rect 6092 8959 6144 8968
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 6276 8959 6328 8968
rect 6276 8925 6285 8959
rect 6285 8925 6319 8959
rect 6319 8925 6328 8959
rect 6276 8916 6328 8925
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 8300 8916 8352 8968
rect 8944 8848 8996 8900
rect 9220 8891 9272 8900
rect 9220 8857 9229 8891
rect 9229 8857 9263 8891
rect 9263 8857 9272 8891
rect 9220 8848 9272 8857
rect 9680 8916 9732 8968
rect 10140 8916 10192 8968
rect 10876 8916 10928 8968
rect 11888 8959 11940 8968
rect 11888 8925 11897 8959
rect 11897 8925 11931 8959
rect 11931 8925 11940 8959
rect 11888 8916 11940 8925
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 9496 8848 9548 8900
rect 10508 8891 10560 8900
rect 10508 8857 10517 8891
rect 10517 8857 10551 8891
rect 10551 8857 10560 8891
rect 10508 8848 10560 8857
rect 3884 8780 3936 8832
rect 4160 8823 4212 8832
rect 4160 8789 4169 8823
rect 4169 8789 4203 8823
rect 4203 8789 4212 8823
rect 4160 8780 4212 8789
rect 5172 8823 5224 8832
rect 5172 8789 5181 8823
rect 5181 8789 5215 8823
rect 5215 8789 5224 8823
rect 5172 8780 5224 8789
rect 5540 8780 5592 8832
rect 6368 8780 6420 8832
rect 7748 8823 7800 8832
rect 7748 8789 7757 8823
rect 7757 8789 7791 8823
rect 7791 8789 7800 8823
rect 7748 8780 7800 8789
rect 9588 8780 9640 8832
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 10784 8780 10836 8832
rect 11152 8848 11204 8900
rect 14188 8848 14240 8900
rect 12348 8780 12400 8832
rect 13912 8823 13964 8832
rect 13912 8789 13921 8823
rect 13921 8789 13955 8823
rect 13955 8789 13964 8823
rect 13912 8780 13964 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 1676 8576 1728 8628
rect 2228 8576 2280 8628
rect 5540 8576 5592 8628
rect 6276 8576 6328 8628
rect 8300 8576 8352 8628
rect 12440 8576 12492 8628
rect 4712 8440 4764 8492
rect 1584 8415 1636 8424
rect 1584 8381 1593 8415
rect 1593 8381 1627 8415
rect 1627 8381 1636 8415
rect 1584 8372 1636 8381
rect 2780 8372 2832 8424
rect 5632 8440 5684 8492
rect 6184 8508 6236 8560
rect 7748 8508 7800 8560
rect 9220 8508 9272 8560
rect 14096 8508 14148 8560
rect 6920 8440 6972 8492
rect 7564 8483 7616 8492
rect 7564 8449 7573 8483
rect 7573 8449 7607 8483
rect 7607 8449 7616 8483
rect 7564 8440 7616 8449
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 4804 8304 4856 8356
rect 9404 8372 9456 8424
rect 10048 8483 10100 8492
rect 10048 8449 10057 8483
rect 10057 8449 10091 8483
rect 10091 8449 10100 8483
rect 10048 8440 10100 8449
rect 12440 8440 12492 8492
rect 5448 8304 5500 8356
rect 4896 8236 4948 8288
rect 5632 8236 5684 8288
rect 7196 8236 7248 8288
rect 7748 8279 7800 8288
rect 7748 8245 7757 8279
rect 7757 8245 7791 8279
rect 7791 8245 7800 8279
rect 7748 8236 7800 8245
rect 12164 8372 12216 8424
rect 12348 8372 12400 8424
rect 11704 8304 11756 8356
rect 12992 8347 13044 8356
rect 12992 8313 13001 8347
rect 13001 8313 13035 8347
rect 13035 8313 13044 8347
rect 12992 8304 13044 8313
rect 12256 8279 12308 8288
rect 12256 8245 12265 8279
rect 12265 8245 12299 8279
rect 12299 8245 12308 8279
rect 12256 8236 12308 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 1124 7896 1176 7948
rect 4712 8007 4764 8016
rect 4712 7973 4721 8007
rect 4721 7973 4755 8007
rect 4755 7973 4764 8007
rect 4712 7964 4764 7973
rect 6920 8075 6972 8084
rect 6920 8041 6929 8075
rect 6929 8041 6963 8075
rect 6963 8041 6972 8075
rect 6920 8032 6972 8041
rect 8024 8075 8076 8084
rect 8024 8041 8033 8075
rect 8033 8041 8067 8075
rect 8067 8041 8076 8075
rect 8024 8032 8076 8041
rect 2136 7828 2188 7880
rect 3424 7828 3476 7880
rect 4896 7828 4948 7880
rect 6276 7871 6328 7880
rect 6276 7837 6285 7871
rect 6285 7837 6319 7871
rect 6319 7837 6328 7871
rect 6276 7828 6328 7837
rect 7104 7896 7156 7948
rect 6736 7828 6788 7880
rect 7288 7871 7340 7880
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 7748 7964 7800 8016
rect 10508 7964 10560 8016
rect 9036 7896 9088 7948
rect 10876 7828 10928 7880
rect 11244 7828 11296 7880
rect 6920 7760 6972 7812
rect 8116 7760 8168 7812
rect 18328 7803 18380 7812
rect 18328 7769 18337 7803
rect 18337 7769 18371 7803
rect 18371 7769 18380 7803
rect 18328 7760 18380 7769
rect 6644 7692 6696 7744
rect 6736 7692 6788 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 4160 7488 4212 7540
rect 4896 7488 4948 7540
rect 9128 7531 9180 7540
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 9496 7531 9548 7540
rect 9496 7497 9505 7531
rect 9505 7497 9539 7531
rect 9539 7497 9548 7531
rect 9496 7488 9548 7497
rect 12348 7488 12400 7540
rect 1308 7352 1360 7404
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 2228 7352 2280 7361
rect 2780 7395 2832 7404
rect 2780 7361 2789 7395
rect 2789 7361 2823 7395
rect 2823 7361 2832 7395
rect 2780 7352 2832 7361
rect 6184 7420 6236 7472
rect 6736 7420 6788 7472
rect 3884 7352 3936 7404
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 1124 7284 1176 7336
rect 3792 7284 3844 7336
rect 4712 7327 4764 7336
rect 4712 7293 4721 7327
rect 4721 7293 4755 7327
rect 4755 7293 4764 7327
rect 4712 7284 4764 7293
rect 6276 7352 6328 7404
rect 6644 7395 6696 7404
rect 6644 7361 6653 7395
rect 6653 7361 6687 7395
rect 6687 7361 6696 7395
rect 6644 7352 6696 7361
rect 7104 7420 7156 7472
rect 6920 7395 6972 7404
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 8024 7420 8076 7472
rect 8944 7463 8996 7472
rect 8944 7429 8953 7463
rect 8953 7429 8987 7463
rect 8987 7429 8996 7463
rect 8944 7420 8996 7429
rect 6920 7352 6972 7361
rect 7840 7395 7892 7404
rect 7840 7361 7849 7395
rect 7849 7361 7883 7395
rect 7883 7361 7892 7395
rect 7840 7352 7892 7361
rect 9220 7395 9272 7404
rect 9220 7361 9229 7395
rect 9229 7361 9263 7395
rect 9263 7361 9272 7395
rect 9220 7352 9272 7361
rect 9588 7352 9640 7404
rect 10692 7420 10744 7472
rect 10508 7395 10560 7404
rect 10508 7361 10517 7395
rect 10517 7361 10551 7395
rect 10551 7361 10560 7395
rect 10508 7352 10560 7361
rect 10876 7395 10928 7404
rect 10876 7361 10885 7395
rect 10885 7361 10919 7395
rect 10919 7361 10928 7395
rect 10876 7352 10928 7361
rect 11704 7395 11756 7404
rect 11704 7361 11713 7395
rect 11713 7361 11747 7395
rect 11747 7361 11756 7395
rect 11704 7352 11756 7361
rect 12900 7488 12952 7540
rect 15108 7488 15160 7540
rect 18236 7488 18288 7540
rect 13912 7420 13964 7472
rect 14648 7420 14700 7472
rect 2688 7216 2740 7268
rect 8944 7284 8996 7336
rect 9772 7284 9824 7336
rect 10784 7284 10836 7336
rect 11796 7327 11848 7336
rect 11796 7293 11805 7327
rect 11805 7293 11839 7327
rect 11839 7293 11848 7327
rect 11796 7284 11848 7293
rect 12256 7284 12308 7336
rect 13820 7395 13872 7404
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 14096 7395 14148 7404
rect 14096 7361 14105 7395
rect 14105 7361 14139 7395
rect 14139 7361 14148 7395
rect 14096 7352 14148 7361
rect 14188 7395 14240 7404
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14188 7352 14240 7361
rect 13912 7284 13964 7336
rect 5356 7216 5408 7268
rect 5632 7216 5684 7268
rect 7288 7216 7340 7268
rect 8116 7216 8168 7268
rect 11336 7216 11388 7268
rect 5172 7191 5224 7200
rect 5172 7157 5181 7191
rect 5181 7157 5215 7191
rect 5215 7157 5224 7191
rect 5172 7148 5224 7157
rect 6920 7148 6972 7200
rect 9128 7148 9180 7200
rect 9956 7148 10008 7200
rect 13084 7148 13136 7200
rect 14280 7148 14332 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 3884 6944 3936 6996
rect 4896 6876 4948 6928
rect 9128 6987 9180 6996
rect 9128 6953 9137 6987
rect 9137 6953 9171 6987
rect 9171 6953 9180 6987
rect 9128 6944 9180 6953
rect 9588 6944 9640 6996
rect 5448 6808 5500 6860
rect 2872 6740 2924 6792
rect 3424 6740 3476 6792
rect 5172 6740 5224 6792
rect 8760 6876 8812 6928
rect 9220 6876 9272 6928
rect 7748 6783 7800 6792
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 7748 6740 7800 6749
rect 8024 6740 8076 6792
rect 1584 6672 1636 6724
rect 5632 6672 5684 6724
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 9588 6783 9640 6792
rect 9588 6749 9597 6783
rect 9597 6749 9631 6783
rect 9631 6749 9640 6783
rect 9588 6740 9640 6749
rect 9772 6876 9824 6928
rect 13820 6944 13872 6996
rect 9956 6783 10008 6792
rect 9956 6749 9965 6783
rect 9965 6749 9999 6783
rect 9999 6749 10008 6783
rect 9956 6740 10008 6749
rect 11152 6740 11204 6792
rect 11336 6783 11388 6792
rect 11336 6749 11345 6783
rect 11345 6749 11379 6783
rect 11379 6749 11388 6783
rect 11336 6740 11388 6749
rect 11612 6740 11664 6792
rect 12164 6740 12216 6792
rect 12348 6808 12400 6860
rect 12900 6851 12952 6860
rect 12900 6817 12909 6851
rect 12909 6817 12943 6851
rect 12943 6817 12952 6851
rect 12900 6808 12952 6817
rect 12992 6808 13044 6860
rect 13912 6808 13964 6860
rect 2504 6604 2556 6656
rect 4528 6604 4580 6656
rect 6644 6604 6696 6656
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 14372 6783 14424 6792
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 14648 6783 14700 6792
rect 14648 6749 14657 6783
rect 14657 6749 14691 6783
rect 14691 6749 14700 6783
rect 14648 6740 14700 6749
rect 11060 6604 11112 6656
rect 11796 6604 11848 6656
rect 12256 6604 12308 6656
rect 13360 6604 13412 6656
rect 13636 6604 13688 6656
rect 14648 6604 14700 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 6460 6400 6512 6452
rect 9220 6400 9272 6452
rect 14372 6400 14424 6452
rect 1308 6264 1360 6316
rect 2688 6264 2740 6316
rect 5540 6264 5592 6316
rect 6828 6307 6880 6316
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 6920 6264 6972 6316
rect 8024 6264 8076 6316
rect 4712 6196 4764 6248
rect 8944 6264 8996 6316
rect 2780 6128 2832 6180
rect 3700 6128 3752 6180
rect 6644 6171 6696 6180
rect 6644 6137 6653 6171
rect 6653 6137 6687 6171
rect 6687 6137 6696 6171
rect 6644 6128 6696 6137
rect 6736 6171 6788 6180
rect 6736 6137 6745 6171
rect 6745 6137 6779 6171
rect 6779 6137 6788 6171
rect 6736 6128 6788 6137
rect 11060 6307 11112 6316
rect 11060 6273 11069 6307
rect 11069 6273 11103 6307
rect 11103 6273 11112 6307
rect 11060 6264 11112 6273
rect 11152 6307 11204 6316
rect 11152 6273 11161 6307
rect 11161 6273 11195 6307
rect 11195 6273 11204 6307
rect 11152 6264 11204 6273
rect 11336 6264 11388 6316
rect 11612 6307 11664 6316
rect 11612 6273 11621 6307
rect 11621 6273 11655 6307
rect 11655 6273 11664 6307
rect 11612 6264 11664 6273
rect 11796 6307 11848 6316
rect 11796 6273 11805 6307
rect 11805 6273 11839 6307
rect 11839 6273 11848 6307
rect 11796 6264 11848 6273
rect 12256 6264 12308 6316
rect 13084 6264 13136 6316
rect 14096 6332 14148 6384
rect 13360 6307 13412 6316
rect 13360 6273 13369 6307
rect 13369 6273 13403 6307
rect 13403 6273 13412 6307
rect 13360 6264 13412 6273
rect 13544 6307 13596 6316
rect 13544 6273 13553 6307
rect 13553 6273 13587 6307
rect 13587 6273 13596 6307
rect 13544 6264 13596 6273
rect 14188 6196 14240 6248
rect 2596 6060 2648 6112
rect 5356 6060 5408 6112
rect 9404 6128 9456 6180
rect 12440 6128 12492 6180
rect 6920 6060 6972 6112
rect 9220 6060 9272 6112
rect 12072 6103 12124 6112
rect 12072 6069 12081 6103
rect 12081 6069 12115 6103
rect 12115 6069 12124 6103
rect 12072 6060 12124 6069
rect 12532 6060 12584 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 1308 5856 1360 5908
rect 6644 5856 6696 5908
rect 6828 5856 6880 5908
rect 7288 5899 7340 5908
rect 7288 5865 7297 5899
rect 7297 5865 7331 5899
rect 7331 5865 7340 5899
rect 7288 5856 7340 5865
rect 9404 5899 9456 5908
rect 9404 5865 9413 5899
rect 9413 5865 9447 5899
rect 9447 5865 9456 5899
rect 9404 5856 9456 5865
rect 13544 5856 13596 5908
rect 1584 5652 1636 5704
rect 2872 5720 2924 5772
rect 2504 5695 2556 5704
rect 2504 5661 2513 5695
rect 2513 5661 2547 5695
rect 2547 5661 2556 5695
rect 2504 5652 2556 5661
rect 2688 5695 2740 5704
rect 2688 5661 2697 5695
rect 2697 5661 2731 5695
rect 2731 5661 2740 5695
rect 2688 5652 2740 5661
rect 2320 5559 2372 5568
rect 2320 5525 2329 5559
rect 2329 5525 2363 5559
rect 2363 5525 2372 5559
rect 2320 5516 2372 5525
rect 2688 5516 2740 5568
rect 4160 5652 4212 5704
rect 5356 5720 5408 5772
rect 4712 5652 4764 5704
rect 6276 5720 6328 5772
rect 6368 5652 6420 5704
rect 6552 5695 6604 5704
rect 6552 5661 6561 5695
rect 6561 5661 6595 5695
rect 6595 5661 6604 5695
rect 6552 5652 6604 5661
rect 6920 5720 6972 5772
rect 11520 5788 11572 5840
rect 7012 5652 7064 5704
rect 7564 5652 7616 5704
rect 9128 5652 9180 5704
rect 9588 5652 9640 5704
rect 7840 5627 7892 5636
rect 7840 5593 7849 5627
rect 7849 5593 7883 5627
rect 7883 5593 7892 5627
rect 7840 5584 7892 5593
rect 8944 5584 8996 5636
rect 12072 5652 12124 5704
rect 12624 5695 12676 5704
rect 12624 5661 12633 5695
rect 12633 5661 12667 5695
rect 12667 5661 12676 5695
rect 12624 5652 12676 5661
rect 12716 5695 12768 5704
rect 12716 5661 12725 5695
rect 12725 5661 12759 5695
rect 12759 5661 12768 5695
rect 12716 5652 12768 5661
rect 12808 5695 12860 5704
rect 12808 5661 12817 5695
rect 12817 5661 12851 5695
rect 12851 5661 12860 5695
rect 12808 5652 12860 5661
rect 12164 5584 12216 5636
rect 2964 5559 3016 5568
rect 2964 5525 2973 5559
rect 2973 5525 3007 5559
rect 3007 5525 3016 5559
rect 2964 5516 3016 5525
rect 5356 5516 5408 5568
rect 5448 5516 5500 5568
rect 5632 5516 5684 5568
rect 6552 5516 6604 5568
rect 9128 5516 9180 5568
rect 9772 5516 9824 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 5540 5312 5592 5364
rect 6736 5312 6788 5364
rect 2964 5244 3016 5296
rect 3700 5287 3752 5296
rect 3700 5253 3709 5287
rect 3709 5253 3743 5287
rect 3743 5253 3752 5287
rect 3700 5244 3752 5253
rect 1308 5176 1360 5228
rect 3424 5219 3476 5228
rect 3424 5185 3433 5219
rect 3433 5185 3467 5219
rect 3467 5185 3476 5219
rect 3424 5176 3476 5185
rect 5448 5244 5500 5296
rect 6920 5287 6972 5296
rect 6920 5253 6929 5287
rect 6929 5253 6963 5287
rect 6963 5253 6972 5287
rect 6920 5244 6972 5253
rect 7840 5244 7892 5296
rect 10600 5287 10652 5296
rect 10600 5253 10609 5287
rect 10609 5253 10643 5287
rect 10643 5253 10652 5287
rect 10600 5244 10652 5253
rect 2136 4972 2188 5024
rect 4712 5176 4764 5228
rect 4896 5176 4948 5228
rect 5908 5219 5960 5228
rect 5908 5185 5917 5219
rect 5917 5185 5951 5219
rect 5951 5185 5960 5219
rect 5908 5176 5960 5185
rect 6276 5176 6328 5228
rect 6552 5219 6604 5228
rect 6552 5185 6561 5219
rect 6561 5185 6595 5219
rect 6595 5185 6604 5219
rect 6552 5176 6604 5185
rect 6736 5176 6788 5228
rect 7012 5176 7064 5228
rect 7288 5176 7340 5228
rect 4712 4972 4764 5024
rect 4896 4972 4948 5024
rect 5540 4972 5592 5024
rect 9220 5219 9272 5228
rect 9220 5185 9229 5219
rect 9229 5185 9263 5219
rect 9263 5185 9272 5219
rect 9220 5176 9272 5185
rect 10692 5176 10744 5228
rect 7840 5151 7892 5160
rect 7840 5117 7849 5151
rect 7849 5117 7883 5151
rect 7883 5117 7892 5151
rect 7840 5108 7892 5117
rect 9128 5151 9180 5160
rect 9128 5117 9137 5151
rect 9137 5117 9171 5151
rect 9171 5117 9180 5151
rect 9128 5108 9180 5117
rect 10692 5040 10744 5092
rect 10876 5108 10928 5160
rect 11336 5219 11388 5228
rect 11336 5185 11345 5219
rect 11345 5185 11379 5219
rect 11379 5185 11388 5219
rect 11336 5176 11388 5185
rect 12624 5312 12676 5364
rect 12808 5244 12860 5296
rect 12900 5287 12952 5296
rect 12900 5253 12909 5287
rect 12909 5253 12943 5287
rect 12943 5253 12952 5287
rect 12900 5244 12952 5253
rect 11520 5176 11572 5228
rect 12348 5176 12400 5228
rect 12808 5108 12860 5160
rect 13084 5219 13136 5228
rect 13084 5185 13093 5219
rect 13093 5185 13127 5219
rect 13127 5185 13136 5219
rect 13084 5176 13136 5185
rect 14188 5176 14240 5228
rect 12532 5040 12584 5092
rect 12900 5040 12952 5092
rect 9772 4972 9824 5024
rect 13084 4972 13136 5024
rect 13176 5015 13228 5024
rect 13176 4981 13185 5015
rect 13185 4981 13219 5015
rect 13219 4981 13228 5015
rect 13176 4972 13228 4981
rect 14556 4972 14608 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 5908 4768 5960 4820
rect 9128 4768 9180 4820
rect 10784 4700 10836 4752
rect 6184 4632 6236 4684
rect 6736 4675 6788 4684
rect 6736 4641 6745 4675
rect 6745 4641 6779 4675
rect 6779 4641 6788 4675
rect 6736 4632 6788 4641
rect 8484 4675 8536 4684
rect 8484 4641 8493 4675
rect 8493 4641 8527 4675
rect 8527 4641 8536 4675
rect 8484 4632 8536 4641
rect 11336 4632 11388 4684
rect 12532 4675 12584 4684
rect 12532 4641 12541 4675
rect 12541 4641 12575 4675
rect 12575 4641 12584 4675
rect 12532 4632 12584 4641
rect 14556 4675 14608 4684
rect 14556 4641 14565 4675
rect 14565 4641 14599 4675
rect 14599 4641 14608 4675
rect 14556 4632 14608 4641
rect 14740 4675 14792 4684
rect 14740 4641 14749 4675
rect 14749 4641 14783 4675
rect 14783 4641 14792 4675
rect 14740 4632 14792 4641
rect 2044 4607 2096 4616
rect 2044 4573 2053 4607
rect 2053 4573 2087 4607
rect 2087 4573 2096 4607
rect 2044 4564 2096 4573
rect 2136 4564 2188 4616
rect 6920 4564 6972 4616
rect 2504 4496 2556 4548
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 10784 4607 10836 4616
rect 10784 4573 10793 4607
rect 10793 4573 10827 4607
rect 10827 4573 10836 4607
rect 10784 4564 10836 4573
rect 12808 4564 12860 4616
rect 13084 4564 13136 4616
rect 13176 4607 13228 4616
rect 13176 4573 13185 4607
rect 13185 4573 13219 4607
rect 13219 4573 13228 4607
rect 13176 4564 13228 4573
rect 14096 4564 14148 4616
rect 15108 4607 15160 4616
rect 15108 4573 15117 4607
rect 15117 4573 15151 4607
rect 15151 4573 15160 4607
rect 15108 4564 15160 4573
rect 6460 4428 6512 4480
rect 12348 4496 12400 4548
rect 11152 4471 11204 4480
rect 11152 4437 11161 4471
rect 11161 4437 11195 4471
rect 11195 4437 11204 4471
rect 11152 4428 11204 4437
rect 12900 4471 12952 4480
rect 12900 4437 12909 4471
rect 12909 4437 12943 4471
rect 12943 4437 12952 4471
rect 12900 4428 12952 4437
rect 13084 4471 13136 4480
rect 13084 4437 13093 4471
rect 13093 4437 13127 4471
rect 13127 4437 13136 4471
rect 13084 4428 13136 4437
rect 14096 4471 14148 4480
rect 14096 4437 14105 4471
rect 14105 4437 14139 4471
rect 14139 4437 14148 4471
rect 14096 4428 14148 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 1768 4224 1820 4276
rect 2136 4156 2188 4208
rect 2504 4267 2556 4276
rect 2504 4233 2513 4267
rect 2513 4233 2547 4267
rect 2547 4233 2556 4267
rect 2504 4224 2556 4233
rect 5356 4267 5408 4276
rect 5356 4233 5365 4267
rect 5365 4233 5399 4267
rect 5399 4233 5408 4267
rect 5356 4224 5408 4233
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 1952 4088 2004 4097
rect 1400 4020 1452 4072
rect 2044 4020 2096 4072
rect 3976 4088 4028 4140
rect 5080 4088 5132 4140
rect 5448 4131 5500 4140
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 5448 4088 5500 4097
rect 6460 4088 6512 4140
rect 10784 4088 10836 4140
rect 11152 4088 11204 4140
rect 12348 4088 12400 4140
rect 12624 4131 12676 4140
rect 12624 4097 12633 4131
rect 12633 4097 12667 4131
rect 12667 4097 12676 4131
rect 12624 4088 12676 4097
rect 5632 4063 5684 4072
rect 5632 4029 5641 4063
rect 5641 4029 5675 4063
rect 5675 4029 5684 4063
rect 5632 4020 5684 4029
rect 6828 4063 6880 4072
rect 6828 4029 6837 4063
rect 6837 4029 6871 4063
rect 6871 4029 6880 4063
rect 6828 4020 6880 4029
rect 12716 3952 12768 4004
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 5356 3884 5408 3936
rect 7196 3884 7248 3936
rect 18052 3884 18104 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 3332 3612 3384 3664
rect 3976 3612 4028 3664
rect 4252 3680 4304 3732
rect 4436 3680 4488 3732
rect 4712 3680 4764 3732
rect 9036 3723 9088 3732
rect 9036 3689 9045 3723
rect 9045 3689 9079 3723
rect 9079 3689 9088 3723
rect 9036 3680 9088 3689
rect 9772 3680 9824 3732
rect 12164 3723 12216 3732
rect 12164 3689 12173 3723
rect 12173 3689 12207 3723
rect 12207 3689 12216 3723
rect 12164 3680 12216 3689
rect 1584 3544 1636 3596
rect 1308 3476 1360 3528
rect 2044 3519 2096 3528
rect 2044 3485 2053 3519
rect 2053 3485 2087 3519
rect 2087 3485 2096 3519
rect 2044 3476 2096 3485
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 5080 3544 5132 3596
rect 8484 3587 8536 3596
rect 8484 3553 8493 3587
rect 8493 3553 8527 3587
rect 8527 3553 8536 3587
rect 8484 3544 8536 3553
rect 3332 3408 3384 3460
rect 3792 3408 3844 3460
rect 4160 3408 4212 3460
rect 4252 3340 4304 3392
rect 4436 3383 4488 3392
rect 4436 3349 4445 3383
rect 4445 3349 4479 3383
rect 4479 3349 4488 3383
rect 4436 3340 4488 3349
rect 4712 3408 4764 3460
rect 4988 3340 5040 3392
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 9220 3519 9272 3528
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 9772 3519 9824 3528
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 9772 3476 9824 3485
rect 10048 3476 10100 3528
rect 10692 3544 10744 3596
rect 11888 3544 11940 3596
rect 10876 3476 10928 3528
rect 12348 3519 12400 3528
rect 12348 3485 12357 3519
rect 12357 3485 12391 3519
rect 12391 3485 12400 3519
rect 12348 3476 12400 3485
rect 12624 3544 12676 3596
rect 18420 3544 18472 3596
rect 17500 3519 17552 3528
rect 17500 3485 17509 3519
rect 17509 3485 17543 3519
rect 17543 3485 17552 3519
rect 17500 3476 17552 3485
rect 18052 3519 18104 3528
rect 18052 3485 18061 3519
rect 18061 3485 18095 3519
rect 18095 3485 18104 3519
rect 18052 3476 18104 3485
rect 8484 3408 8536 3460
rect 8300 3340 8352 3392
rect 18328 3451 18380 3460
rect 18328 3417 18337 3451
rect 18337 3417 18371 3451
rect 18371 3417 18380 3451
rect 18328 3408 18380 3417
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 2596 3179 2648 3188
rect 2596 3145 2605 3179
rect 2605 3145 2639 3179
rect 2639 3145 2648 3179
rect 2596 3136 2648 3145
rect 4436 3136 4488 3188
rect 5356 3179 5408 3188
rect 5356 3145 5365 3179
rect 5365 3145 5399 3179
rect 5399 3145 5408 3179
rect 5356 3136 5408 3145
rect 9220 3136 9272 3188
rect 9772 3136 9824 3188
rect 10048 3136 10100 3188
rect 10876 3179 10928 3188
rect 10876 3145 10885 3179
rect 10885 3145 10919 3179
rect 10919 3145 10928 3179
rect 10876 3136 10928 3145
rect 11888 3179 11940 3188
rect 11888 3145 11897 3179
rect 11897 3145 11931 3179
rect 11931 3145 11940 3179
rect 11888 3136 11940 3145
rect 12348 3136 12400 3188
rect 12440 3136 12492 3188
rect 13084 3136 13136 3188
rect 1860 2975 1912 2984
rect 1860 2941 1869 2975
rect 1869 2941 1903 2975
rect 1903 2941 1912 2975
rect 1860 2932 1912 2941
rect 2596 2932 2648 2984
rect 2504 2864 2556 2916
rect 3608 2932 3660 2984
rect 4620 3068 4672 3120
rect 5448 3068 5500 3120
rect 6644 3068 6696 3120
rect 4252 3000 4304 3052
rect 4620 2975 4672 2984
rect 4620 2941 4629 2975
rect 4629 2941 4663 2975
rect 4663 2941 4672 2975
rect 4620 2932 4672 2941
rect 5632 3000 5684 3052
rect 8116 3068 8168 3120
rect 12532 3068 12584 3120
rect 12900 3068 12952 3120
rect 6368 2932 6420 2984
rect 8300 3000 8352 3052
rect 8484 2975 8536 2984
rect 8484 2941 8493 2975
rect 8493 2941 8527 2975
rect 8527 2941 8536 2975
rect 8484 2932 8536 2941
rect 17592 3000 17644 3052
rect 18512 3043 18564 3052
rect 18512 3009 18521 3043
rect 18521 3009 18555 3043
rect 18555 3009 18564 3043
rect 18512 3000 18564 3009
rect 14740 2932 14792 2984
rect 17408 2932 17460 2984
rect 17960 2932 18012 2984
rect 12532 2864 12584 2916
rect 3976 2796 4028 2848
rect 10324 2796 10376 2848
rect 11336 2796 11388 2848
rect 11520 2839 11572 2848
rect 11520 2805 11529 2839
rect 11529 2805 11563 2839
rect 11563 2805 11572 2839
rect 11520 2796 11572 2805
rect 12624 2796 12676 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 1952 2592 2004 2644
rect 3792 2592 3844 2644
rect 4620 2592 4672 2644
rect 2320 2499 2372 2508
rect 2320 2465 2329 2499
rect 2329 2465 2363 2499
rect 2363 2465 2372 2499
rect 2320 2456 2372 2465
rect 2596 2456 2648 2508
rect 1308 2388 1360 2440
rect 4068 2456 4120 2508
rect 4712 2456 4764 2508
rect 5264 2456 5316 2508
rect 1216 2320 1268 2372
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 3884 2388 3936 2440
rect 8116 2524 8168 2576
rect 5816 2456 5868 2508
rect 5724 2431 5776 2440
rect 5724 2397 5733 2431
rect 5733 2397 5767 2431
rect 5767 2397 5776 2431
rect 5724 2388 5776 2397
rect 7656 2431 7708 2440
rect 7656 2397 7665 2431
rect 7665 2397 7699 2431
rect 7699 2397 7708 2431
rect 7656 2388 7708 2397
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 8760 2431 8812 2440
rect 8760 2397 8769 2431
rect 8769 2397 8803 2431
rect 8803 2397 8812 2431
rect 8760 2388 8812 2397
rect 9772 2388 9824 2440
rect 11428 2456 11480 2508
rect 14740 2456 14792 2508
rect 15752 2456 15804 2508
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 11336 2431 11388 2440
rect 11336 2397 11345 2431
rect 11345 2397 11379 2431
rect 11379 2397 11388 2431
rect 11336 2388 11388 2397
rect 11520 2431 11572 2440
rect 11520 2397 11529 2431
rect 11529 2397 11563 2431
rect 11563 2397 11572 2431
rect 11520 2388 11572 2397
rect 12532 2431 12584 2440
rect 12532 2397 12541 2431
rect 12541 2397 12575 2431
rect 12575 2397 12584 2431
rect 12532 2388 12584 2397
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 13636 2431 13688 2440
rect 13636 2397 13645 2431
rect 13645 2397 13679 2431
rect 13679 2397 13688 2431
rect 13636 2388 13688 2397
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 14648 2431 14700 2440
rect 14648 2397 14657 2431
rect 14657 2397 14691 2431
rect 14691 2397 14700 2431
rect 14648 2388 14700 2397
rect 15568 2388 15620 2440
rect 16212 2431 16264 2440
rect 16212 2397 16221 2431
rect 16221 2397 16255 2431
rect 16255 2397 16264 2431
rect 16212 2388 16264 2397
rect 16672 2431 16724 2440
rect 16672 2397 16681 2431
rect 16681 2397 16715 2431
rect 16715 2397 16724 2431
rect 16672 2388 16724 2397
rect 17224 2431 17276 2440
rect 17224 2397 17233 2431
rect 17233 2397 17267 2431
rect 17267 2397 17276 2431
rect 17224 2388 17276 2397
rect 17776 2431 17828 2440
rect 17776 2397 17785 2431
rect 17785 2397 17819 2431
rect 17819 2397 17828 2431
rect 17776 2388 17828 2397
rect 3056 2320 3108 2372
rect 4160 2320 4212 2372
rect 4712 2320 4764 2372
rect 5264 2320 5316 2372
rect 5816 2320 5868 2372
rect 6920 2363 6972 2372
rect 6920 2329 6929 2363
rect 6929 2329 6963 2363
rect 6963 2329 6972 2363
rect 6920 2320 6972 2329
rect 7472 2320 7524 2372
rect 8024 2320 8076 2372
rect 8576 2320 8628 2372
rect 9128 2320 9180 2372
rect 10784 2320 10836 2372
rect 11888 2320 11940 2372
rect 12440 2320 12492 2372
rect 12992 2320 13044 2372
rect 13544 2320 13596 2372
rect 3424 2252 3476 2304
rect 3976 2252 4028 2304
rect 9680 2252 9732 2304
rect 10232 2252 10284 2304
rect 11336 2252 11388 2304
rect 14096 2252 14148 2304
rect 15200 2252 15252 2304
rect 16304 2320 16356 2372
rect 16856 2252 16908 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 1398 19200 1454 20000
rect 1950 19200 2006 20000
rect 2502 19200 2558 20000
rect 3054 19200 3110 20000
rect 3606 19200 3662 20000
rect 4158 19200 4214 20000
rect 4710 19200 4766 20000
rect 5262 19200 5318 20000
rect 5814 19200 5870 20000
rect 6366 19200 6422 20000
rect 6918 19200 6974 20000
rect 7470 19200 7526 20000
rect 8022 19200 8078 20000
rect 8574 19200 8630 20000
rect 9126 19200 9182 20000
rect 9678 19200 9734 20000
rect 10230 19200 10286 20000
rect 10782 19200 10838 20000
rect 11334 19200 11390 20000
rect 11886 19200 11942 20000
rect 12438 19200 12494 20000
rect 12990 19200 13046 20000
rect 13542 19200 13598 20000
rect 14094 19200 14150 20000
rect 14646 19200 14702 20000
rect 15198 19200 15254 20000
rect 15750 19200 15806 20000
rect 16302 19200 16358 20000
rect 16854 19200 16910 20000
rect 17406 19200 17462 20000
rect 17958 19200 18014 20000
rect 18510 19200 18566 20000
rect 1412 18170 1440 19200
rect 1412 18142 1532 18170
rect 1398 18048 1454 18057
rect 1398 17983 1454 17992
rect 1308 17128 1360 17134
rect 1308 17070 1360 17076
rect 1320 16969 1348 17070
rect 1306 16960 1362 16969
rect 1306 16895 1362 16904
rect 1320 16658 1348 16895
rect 1308 16652 1360 16658
rect 1308 16594 1360 16600
rect 1412 16590 1440 17983
rect 1504 17202 1532 18142
rect 1964 17270 1992 19200
rect 2516 17338 2544 19200
rect 3068 17338 3096 19200
rect 3620 17338 3648 19200
rect 2504 17332 2556 17338
rect 2504 17274 2556 17280
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 4172 17270 4200 19200
rect 1952 17264 2004 17270
rect 1952 17206 2004 17212
rect 4160 17264 4212 17270
rect 4160 17206 4212 17212
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 1400 16584 1452 16590
rect 1400 16526 1452 16532
rect 1504 16250 1532 17138
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1688 16726 1716 16934
rect 1964 16794 1992 17206
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 2044 16992 2096 16998
rect 2044 16934 2096 16940
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 1676 16720 1728 16726
rect 1676 16662 1728 16668
rect 1688 16574 1716 16662
rect 1688 16546 1808 16574
rect 1492 16244 1544 16250
rect 1492 16186 1544 16192
rect 1308 16108 1360 16114
rect 1308 16050 1360 16056
rect 1320 15881 1348 16050
rect 1306 15872 1362 15881
rect 1306 15807 1362 15816
rect 1308 15020 1360 15026
rect 1308 14962 1360 14968
rect 1320 14793 1348 14962
rect 1306 14784 1362 14793
rect 1306 14719 1362 14728
rect 1308 13932 1360 13938
rect 1308 13874 1360 13880
rect 1320 13705 1348 13874
rect 1584 13728 1636 13734
rect 1306 13696 1362 13705
rect 1584 13670 1636 13676
rect 1306 13631 1362 13640
rect 1308 12844 1360 12850
rect 1308 12786 1360 12792
rect 1320 12617 1348 12786
rect 1306 12608 1362 12617
rect 1306 12543 1362 12552
rect 1308 11756 1360 11762
rect 1308 11698 1360 11704
rect 1320 11529 1348 11698
rect 1306 11520 1362 11529
rect 1306 11455 1362 11464
rect 1596 11082 1624 13670
rect 1584 11076 1636 11082
rect 1584 11018 1636 11024
rect 1308 10668 1360 10674
rect 1308 10610 1360 10616
rect 1320 10441 1348 10610
rect 1306 10432 1362 10441
rect 1306 10367 1362 10376
rect 1308 10056 1360 10062
rect 1308 9998 1360 10004
rect 1320 9353 1348 9998
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1596 9586 1624 9862
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1306 9344 1362 9353
rect 1306 9279 1362 9288
rect 1596 8974 1624 9522
rect 1688 9042 1716 9522
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1688 8634 1716 8978
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1122 8256 1178 8265
rect 1122 8191 1178 8200
rect 1136 7954 1164 8191
rect 1124 7948 1176 7954
rect 1124 7890 1176 7896
rect 1136 7342 1164 7890
rect 1596 7546 1624 8366
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1308 7404 1360 7410
rect 1308 7346 1360 7352
rect 1124 7336 1176 7342
rect 1124 7278 1176 7284
rect 1320 7177 1348 7346
rect 1306 7168 1362 7177
rect 1306 7103 1362 7112
rect 1584 6724 1636 6730
rect 1584 6666 1636 6672
rect 1596 6458 1624 6666
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 1320 6089 1348 6258
rect 1306 6080 1362 6089
rect 1306 6015 1362 6024
rect 1320 5914 1348 6015
rect 1308 5908 1360 5914
rect 1308 5850 1360 5856
rect 1596 5710 1624 6394
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1308 5228 1360 5234
rect 1308 5170 1360 5176
rect 1320 5001 1348 5170
rect 1306 4992 1362 5001
rect 1306 4927 1362 4936
rect 1780 4282 1808 16546
rect 2056 4622 2084 16934
rect 2688 9648 2740 9654
rect 2740 9596 2912 9602
rect 2688 9590 2912 9596
rect 2700 9586 2912 9590
rect 3436 9586 3464 17138
rect 4172 17082 4200 17206
rect 4724 17202 4752 19200
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 5276 17202 5304 19200
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 5264 17196 5316 17202
rect 5828 17184 5856 19200
rect 6380 17270 6408 19200
rect 6736 17332 6788 17338
rect 6736 17274 6788 17280
rect 6368 17264 6420 17270
rect 6368 17206 6420 17212
rect 5908 17196 5960 17202
rect 5828 17156 5908 17184
rect 5264 17138 5316 17144
rect 5908 17138 5960 17144
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 4080 17054 4200 17082
rect 4620 17060 4672 17066
rect 3516 16992 3568 16998
rect 3516 16934 3568 16940
rect 3884 16992 3936 16998
rect 3884 16934 3936 16940
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2320 9580 2372 9586
rect 2700 9580 2924 9586
rect 2700 9574 2872 9580
rect 2320 9522 2372 9528
rect 2872 9522 2924 9528
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 2148 7886 2176 9522
rect 2332 9178 2360 9522
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2240 7410 2268 8570
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2792 7410 2820 8366
rect 3436 7886 3464 9522
rect 3528 9110 3556 16934
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3804 11694 3832 12174
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3528 8974 3556 9046
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2688 7268 2740 7274
rect 2688 7210 2740 7216
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2516 5710 2544 6598
rect 2700 6322 2728 7210
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2320 5568 2372 5574
rect 2320 5510 2372 5516
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2148 4622 2176 4966
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 1768 4276 1820 4282
rect 1768 4218 1820 4224
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1400 4072 1452 4078
rect 1400 4014 1452 4020
rect 1306 3904 1362 3913
rect 1306 3839 1362 3848
rect 1320 3534 1348 3839
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1306 2816 1362 2825
rect 1306 2751 1362 2760
rect 1320 2446 1348 2751
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 1216 2372 1268 2378
rect 1216 2314 1268 2320
rect 1228 1737 1256 2314
rect 1214 1728 1270 1737
rect 1214 1663 1270 1672
rect 1412 800 1440 4014
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 1596 2650 1624 3538
rect 1860 2984 1912 2990
rect 1860 2926 1912 2932
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1872 1578 1900 2926
rect 1964 2650 1992 4082
rect 2056 4078 2084 4558
rect 2148 4214 2176 4558
rect 2136 4208 2188 4214
rect 2136 4150 2188 4156
rect 2044 4072 2096 4078
rect 2044 4014 2096 4020
rect 2056 3534 2084 4014
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 2332 2514 2360 5510
rect 2504 4548 2556 4554
rect 2504 4490 2556 4496
rect 2516 4282 2544 4490
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2608 3194 2636 6054
rect 2700 5710 2728 6258
rect 2792 6186 2820 7346
rect 3436 6798 3464 7822
rect 3804 7342 3832 8842
rect 3896 8838 3924 16934
rect 4080 16776 4108 17054
rect 4620 17002 4672 17008
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4160 16788 4212 16794
rect 4080 16748 4160 16776
rect 4160 16730 4212 16736
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4080 14482 4108 14962
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 4528 14476 4580 14482
rect 4528 14418 4580 14424
rect 4540 14006 4568 14418
rect 4528 14000 4580 14006
rect 4528 13942 4580 13948
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4080 12434 4108 13330
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3988 12406 4108 12434
rect 3988 11694 4016 12406
rect 4080 12374 4108 12406
rect 4068 12368 4120 12374
rect 4068 12310 4120 12316
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 4264 11898 4292 12106
rect 4448 11898 4476 12242
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 3988 10810 4016 11630
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10266 4660 17002
rect 4724 16794 4752 17138
rect 6276 17060 6328 17066
rect 6276 17002 6328 17008
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4816 15722 4844 16934
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4988 16040 5040 16046
rect 4988 15982 5040 15988
rect 4724 15694 4844 15722
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9178 4660 9862
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4724 9110 4752 15694
rect 5000 15570 5028 15982
rect 4988 15564 5040 15570
rect 4816 15524 4988 15552
rect 4816 15026 4844 15524
rect 4988 15506 5040 15512
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 5276 14958 5304 15438
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4896 13796 4948 13802
rect 4896 13738 4948 13744
rect 4908 13530 4936 13738
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4816 12434 4844 13262
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 5368 12434 5396 16934
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5632 16516 5684 16522
rect 5632 16458 5684 16464
rect 5644 16114 5672 16458
rect 5828 16114 5856 16526
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5644 15502 5672 15846
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 5448 14884 5500 14890
rect 5448 14826 5500 14832
rect 5460 13326 5488 14826
rect 5552 14414 5580 15030
rect 5920 14770 5948 16934
rect 5920 14742 6040 14770
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5460 12850 5488 13262
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 4816 12406 5028 12434
rect 4816 11830 4844 12406
rect 5000 12102 5028 12406
rect 5276 12406 5396 12434
rect 5080 12368 5132 12374
rect 5080 12310 5132 12316
rect 5092 12102 5120 12310
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4896 10192 4948 10198
rect 4896 10134 4948 10140
rect 4908 10010 4936 10134
rect 4816 9982 5028 10010
rect 4712 9104 4764 9110
rect 4632 9052 4712 9058
rect 4632 9046 4764 9052
rect 4632 9030 4752 9046
rect 4632 8906 4660 9030
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 3896 7410 3924 8774
rect 4172 8378 4200 8774
rect 4724 8498 4752 8842
rect 4816 8616 4844 9982
rect 5000 9926 5028 9982
rect 5276 9926 5304 12406
rect 5552 12170 5580 13126
rect 5644 12306 5672 13670
rect 5736 13326 5764 14010
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5828 12434 5856 13670
rect 5920 13530 5948 13874
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 6012 12434 6040 14742
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 5736 12406 5856 12434
rect 5920 12406 6040 12434
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5368 10266 5396 10542
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5552 9722 5580 9930
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5644 9722 5672 9862
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 4908 9178 4936 9318
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 5170 8936 5226 8945
rect 5170 8871 5226 8880
rect 5184 8838 5212 8871
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4816 8588 4936 8616
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4080 8350 4200 8378
rect 4080 7970 4108 8350
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4724 8022 4752 8434
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 4712 8016 4764 8022
rect 4080 7942 4200 7970
rect 4712 7958 4764 7964
rect 4172 7546 4200 7942
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3896 7002 3924 7346
rect 4172 7256 4200 7482
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4080 7228 4200 7256
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 4080 6882 4108 7228
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4080 6854 4200 6882
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 2780 6180 2832 6186
rect 2780 6122 2832 6128
rect 2884 5778 2912 6734
rect 3700 6180 3752 6186
rect 3700 6122 3752 6128
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 2700 5574 2728 5646
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2976 5302 3004 5510
rect 3712 5302 3740 6122
rect 4172 6100 4200 6854
rect 4528 6656 4580 6662
rect 4580 6616 4660 6644
rect 4528 6598 4580 6604
rect 4080 6072 4200 6100
rect 4080 5794 4108 6072
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4080 5766 4200 5794
rect 4172 5710 4200 5766
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 2964 5296 3016 5302
rect 2964 5238 3016 5244
rect 3700 5296 3752 5302
rect 3700 5238 3752 5244
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3332 3664 3384 3670
rect 3332 3606 3384 3612
rect 3344 3466 3372 3606
rect 3332 3460 3384 3466
rect 3332 3402 3384 3408
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 2320 2508 2372 2514
rect 2320 2450 2372 2456
rect 1872 1550 1992 1578
rect 1964 800 1992 1550
rect 2516 800 2544 2858
rect 2608 2514 2636 2926
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 3056 2372 3108 2378
rect 3056 2314 3108 2320
rect 3068 800 3096 2314
rect 3436 2310 3464 5170
rect 4172 5080 4200 5646
rect 4080 5052 4200 5080
rect 4080 4706 4108 5052
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4080 4678 4200 4706
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3988 3670 4016 4082
rect 4172 3992 4200 4678
rect 4080 3964 4200 3992
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 4080 3618 4108 3964
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4264 3618 4292 3674
rect 3988 3534 4016 3606
rect 4080 3590 4292 3618
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3792 3460 3844 3466
rect 3792 3402 3844 3408
rect 3608 2984 3660 2990
rect 3608 2926 3660 2932
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3620 800 3648 2926
rect 3804 2650 3832 3402
rect 3988 3346 4016 3470
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 3896 3318 4016 3346
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3804 2446 3832 2586
rect 3896 2446 3924 3318
rect 3976 2848 4028 2854
rect 4172 2836 4200 3402
rect 4448 3398 4476 3674
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4264 3058 4292 3334
rect 4448 3194 4476 3334
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4632 3126 4660 6616
rect 4724 6254 4752 7278
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4724 5710 4752 6190
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4724 5030 4752 5170
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4724 3738 4752 4966
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4620 2984 4672 2990
rect 4724 2972 4752 3402
rect 4672 2944 4752 2972
rect 4620 2926 4672 2932
rect 3976 2790 4028 2796
rect 4080 2808 4200 2836
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 3988 2310 4016 2790
rect 4080 2514 4108 2808
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2650 4660 2926
rect 4816 2774 4844 8298
rect 4908 8294 4936 8588
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4908 7886 4936 8230
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4908 7410 4936 7482
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4908 6934 4936 7346
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 5184 6798 5212 7142
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4908 5030 4936 5170
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 5000 3398 5028 3878
rect 5092 3602 5120 4082
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4724 2746 4844 2774
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4724 2514 4752 2746
rect 5276 2514 5304 9318
rect 5356 8968 5408 8974
rect 5460 8945 5488 9454
rect 5356 8910 5408 8916
rect 5446 8936 5502 8945
rect 5368 7274 5396 8910
rect 5446 8871 5502 8880
rect 5632 8900 5684 8906
rect 5460 8480 5488 8871
rect 5632 8842 5684 8848
rect 5540 8832 5592 8838
rect 5644 8809 5672 8842
rect 5540 8774 5592 8780
rect 5630 8800 5686 8809
rect 5552 8634 5580 8774
rect 5630 8735 5686 8744
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5632 8492 5684 8498
rect 5460 8452 5632 8480
rect 5632 8434 5684 8440
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 5368 6118 5396 7210
rect 5460 6866 5488 8298
rect 5644 8294 5672 8434
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5632 7268 5684 7274
rect 5632 7210 5684 7216
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5368 5778 5396 6054
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5460 5574 5488 6802
rect 5644 6730 5672 7210
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5368 4282 5396 5510
rect 5552 5370 5580 6258
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5460 4146 5488 5238
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5552 4026 5580 4966
rect 5644 4078 5672 5510
rect 5460 3998 5580 4026
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5368 3194 5396 3878
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5460 3126 5488 3998
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5644 3058 5672 4014
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 5736 2446 5764 12406
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5828 2514 5856 11290
rect 5920 10742 5948 12406
rect 6104 12306 6132 12582
rect 6288 12434 6316 17002
rect 6564 15502 6592 17138
rect 6644 17128 6696 17134
rect 6644 17070 6696 17076
rect 6656 16590 6684 17070
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6748 15570 6776 17274
rect 6932 17270 6960 19200
rect 7012 17740 7064 17746
rect 7012 17682 7064 17688
rect 7024 17338 7052 17682
rect 7484 17338 7512 19200
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 7472 17332 7524 17338
rect 7472 17274 7524 17280
rect 6920 17264 6972 17270
rect 6920 17206 6972 17212
rect 6932 17082 6960 17206
rect 7024 17202 7052 17274
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 6932 17054 7052 17082
rect 6920 16992 6972 16998
rect 6920 16934 6972 16940
rect 6932 16658 6960 16934
rect 7024 16794 7052 17054
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 6932 16114 6960 16594
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 7024 16046 7052 16526
rect 7484 16250 7512 16526
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6460 15428 6512 15434
rect 6460 15370 6512 15376
rect 6472 14958 6500 15370
rect 6748 15162 6776 15506
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6472 14482 6500 14894
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6748 14414 6776 14962
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6748 12442 6776 14350
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6932 14006 6960 14214
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 6840 13530 6868 13874
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6736 12436 6788 12442
rect 6288 12406 6408 12434
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 6012 11286 6040 12242
rect 6000 11280 6052 11286
rect 6000 11222 6052 11228
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6092 9988 6144 9994
rect 6092 9930 6144 9936
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 6012 9586 6040 9862
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6104 8974 6132 9930
rect 6196 9586 6224 9998
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6288 9586 6316 9862
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6196 9042 6224 9522
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6182 8800 6238 8809
rect 6182 8735 6238 8744
rect 6196 8566 6224 8735
rect 6288 8634 6316 8910
rect 6380 8838 6408 12406
rect 6736 12378 6788 12384
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6184 8560 6236 8566
rect 6184 8502 6236 8508
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 5920 4826 5948 5170
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 6196 4690 6224 7414
rect 6288 7410 6316 7822
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6472 6458 6500 8910
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6564 5794 6592 12038
rect 6748 11762 6776 12378
rect 7208 12102 7236 13874
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 7208 11150 7236 12038
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7300 11218 7328 11494
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6840 10198 6868 10406
rect 6828 10192 6880 10198
rect 6828 10134 6880 10140
rect 6840 10062 6868 10134
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6656 9042 6684 9522
rect 6840 9518 6868 9998
rect 6932 9586 6960 10066
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 7576 8498 7604 16934
rect 7760 16658 7788 17478
rect 8036 17338 8064 19200
rect 8588 17338 8616 19200
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 8576 17332 8628 17338
rect 8576 17274 8628 17280
rect 9140 17202 9168 19200
rect 9692 17338 9720 19200
rect 10244 17338 10272 19200
rect 10796 17338 10824 19200
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 11348 17202 11376 19200
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11704 17128 11756 17134
rect 11702 17096 11704 17105
rect 11796 17128 11848 17134
rect 11756 17096 11758 17105
rect 10048 17060 10100 17066
rect 10048 17002 10100 17008
rect 10692 17060 10744 17066
rect 11796 17070 11848 17076
rect 11702 17031 11758 17040
rect 10692 17002 10744 17008
rect 7932 16992 7984 16998
rect 7932 16934 7984 16940
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 7748 16652 7800 16658
rect 7748 16594 7800 16600
rect 7944 12434 7972 16934
rect 8760 16652 8812 16658
rect 8760 16594 8812 16600
rect 8772 16250 8800 16594
rect 8760 16244 8812 16250
rect 8760 16186 8812 16192
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 7852 12406 7972 12434
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 6932 8090 6960 8434
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6748 7750 6776 7822
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6656 7410 6684 7686
rect 6748 7478 6776 7686
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6932 7410 6960 7754
rect 7116 7478 7144 7890
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6656 6662 6684 7346
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6932 6322 6960 7142
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6644 6180 6696 6186
rect 6644 6122 6696 6128
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6656 5914 6684 6122
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6276 5772 6328 5778
rect 6564 5766 6684 5794
rect 6276 5714 6328 5720
rect 6288 5234 6316 5714
rect 6368 5704 6420 5710
rect 6552 5704 6604 5710
rect 6420 5664 6552 5692
rect 6368 5646 6420 5652
rect 6552 5646 6604 5652
rect 6564 5574 6592 5646
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6564 5234 6592 5510
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6472 4146 6500 4422
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6656 3126 6684 5766
rect 6748 5370 6776 6122
rect 6840 5914 6868 6258
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6932 5778 6960 6054
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6748 4690 6776 5170
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6748 4026 6776 4626
rect 6932 4622 6960 5238
rect 7024 5234 7052 5646
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6828 4072 6880 4078
rect 6748 4020 6828 4026
rect 6748 4014 6880 4020
rect 6748 3998 6868 4014
rect 7208 3942 7236 8230
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7300 7274 7328 7822
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 7300 5914 7328 7210
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7300 5234 7328 5850
rect 7576 5710 7604 8434
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 4712 2372 4764 2378
rect 4712 2314 4764 2320
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 4172 800 4200 2314
rect 4724 800 4752 2314
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5276 800 5304 2314
rect 5828 800 5856 2314
rect 6380 800 6408 2926
rect 7668 2446 7696 11494
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7760 8566 7788 8774
rect 7748 8560 7800 8566
rect 7748 8502 7800 8508
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 8022 7788 8230
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7852 7410 7880 12406
rect 8220 11014 8248 15914
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8496 15366 8524 15846
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8668 15360 8720 15366
rect 8772 15337 8800 15846
rect 8852 15428 8904 15434
rect 8852 15370 8904 15376
rect 8668 15302 8720 15308
rect 8758 15328 8814 15337
rect 8496 15026 8524 15302
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8588 14958 8616 15302
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8392 14884 8444 14890
rect 8392 14826 8444 14832
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8312 12986 8340 13942
rect 8404 13326 8432 14826
rect 8680 13870 8708 15302
rect 8758 15263 8814 15272
rect 8864 15094 8892 15370
rect 8852 15088 8904 15094
rect 8852 15030 8904 15036
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8668 13456 8720 13462
rect 8668 13398 8720 13404
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8312 12374 8340 12786
rect 8496 12442 8524 13126
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8588 12102 8616 13262
rect 8680 12782 8708 13398
rect 8772 13190 8800 14826
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8680 12306 8708 12378
rect 8668 12300 8720 12306
rect 8668 12242 8720 12248
rect 8772 12170 8800 13126
rect 8864 12986 8892 13874
rect 8956 13841 8984 14214
rect 8942 13832 8998 13841
rect 8942 13767 8998 13776
rect 8944 13456 8996 13462
rect 8944 13398 8996 13404
rect 8852 12980 8904 12986
rect 8852 12922 8904 12928
rect 8852 12844 8904 12850
rect 8956 12834 8984 13398
rect 8852 12786 8904 12792
rect 8944 12828 8996 12834
rect 8864 12374 8892 12786
rect 8944 12770 8996 12776
rect 8852 12368 8904 12374
rect 8852 12310 8904 12316
rect 8760 12164 8812 12170
rect 8760 12106 8812 12112
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8588 11694 8616 12038
rect 8956 11898 8984 12038
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8772 11218 8800 11630
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 8404 10266 8432 10474
rect 9048 10470 9076 16934
rect 9220 16720 9272 16726
rect 9220 16662 9272 16668
rect 9232 16046 9260 16662
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9232 14482 9260 15982
rect 9324 15638 9352 16186
rect 9312 15632 9364 15638
rect 9312 15574 9364 15580
rect 9324 15026 9352 15574
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9128 12912 9180 12918
rect 9128 12854 9180 12860
rect 9140 12238 9168 12854
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9232 11694 9260 14418
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9508 14006 9536 14214
rect 9496 14000 9548 14006
rect 9496 13942 9548 13948
rect 9404 13456 9456 13462
rect 9404 13398 9456 13404
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 9324 12306 9352 12650
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9416 12238 9444 13398
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9508 11830 9536 12038
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9324 11218 9352 11562
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7760 5148 7788 6734
rect 7840 5636 7892 5642
rect 7840 5578 7892 5584
rect 7852 5302 7880 5578
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 7840 5160 7892 5166
rect 7760 5120 7840 5148
rect 7840 5102 7892 5108
rect 7944 4570 7972 9862
rect 8036 9586 8064 9862
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8036 9042 8064 9522
rect 8312 9450 8340 9930
rect 8404 9654 8432 10202
rect 9600 9994 9628 16934
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9784 16114 9812 16390
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9784 15638 9812 16050
rect 9864 15972 9916 15978
rect 9864 15914 9916 15920
rect 9772 15632 9824 15638
rect 9772 15574 9824 15580
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9692 14414 9720 15438
rect 9784 15162 9812 15438
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9784 14550 9812 15098
rect 9772 14544 9824 14550
rect 9772 14486 9824 14492
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9692 14074 9720 14350
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9692 11150 9720 11630
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9588 9988 9640 9994
rect 9588 9930 9640 9936
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 8404 9330 8432 9590
rect 8312 9302 8432 9330
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8036 8090 8064 8978
rect 8312 8974 8340 9302
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8312 8634 8340 8910
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8036 7478 8064 8026
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 8128 7274 8156 7754
rect 8956 7478 8984 8842
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 8944 7472 8996 7478
rect 8944 7414 8996 7420
rect 8956 7342 8984 7414
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8116 7268 8168 7274
rect 8116 7210 8168 7216
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8772 6798 8800 6870
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8036 6322 8064 6734
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8956 5642 8984 6258
rect 8944 5636 8996 5642
rect 8944 5578 8996 5584
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8392 4616 8444 4622
rect 8312 4576 8392 4604
rect 7944 4542 8064 4570
rect 8036 2774 8064 4542
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8128 3126 8156 3470
rect 8312 3398 8340 4576
rect 8392 4558 8444 4564
rect 8496 3602 8524 4626
rect 9048 3738 9076 7890
rect 9140 7546 9168 9046
rect 9232 8906 9260 9658
rect 9600 9586 9628 9930
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9220 8900 9272 8906
rect 9220 8842 9272 8848
rect 9232 8566 9260 8842
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 9416 8430 9444 9114
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9508 8498 9536 8842
rect 9600 8838 9628 9522
rect 9692 8974 9720 10678
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9508 7546 9536 8434
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9140 7206 9168 7482
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9140 6100 9168 6938
rect 9232 6934 9260 7346
rect 9600 7002 9628 7346
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9220 6928 9272 6934
rect 9220 6870 9272 6876
rect 9600 6798 9628 6938
rect 9784 6934 9812 7278
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9232 6458 9260 6734
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9220 6112 9272 6118
rect 9140 6072 9220 6100
rect 9220 6054 9272 6060
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9140 5574 9168 5646
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9140 5166 9168 5510
rect 9232 5234 9260 6054
rect 9416 5914 9444 6122
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9600 5710 9628 6734
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 9140 4826 9168 5102
rect 9784 5030 9812 5510
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 9784 3534 9812 3674
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 8484 3460 8536 3466
rect 8484 3402 8536 3408
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 8312 3058 8340 3334
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8496 2990 8524 3402
rect 9232 3194 9260 3470
rect 9784 3194 9812 3470
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 9876 2774 9904 15914
rect 9968 15502 9996 16594
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9968 14958 9996 15438
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 9968 14618 9996 14894
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9968 14414 9996 14554
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 10060 12434 10088 17002
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10060 12406 10180 12434
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 9968 7290 9996 9114
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 10060 8498 10088 8978
rect 10152 8974 10180 12406
rect 10244 10062 10272 16934
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10428 15502 10456 15846
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10508 15428 10560 15434
rect 10612 15416 10640 15982
rect 10560 15388 10640 15416
rect 10508 15370 10560 15376
rect 10612 14550 10640 15388
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10428 14074 10456 14350
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10336 11762 10364 12582
rect 10704 11762 10732 17002
rect 11336 16992 11388 16998
rect 11336 16934 11388 16940
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 11072 16538 11100 16594
rect 10888 16510 11100 16538
rect 10888 16454 10916 16510
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 11072 16046 11100 16510
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11150 16280 11206 16289
rect 11150 16215 11206 16224
rect 11164 16182 11192 16215
rect 11152 16176 11204 16182
rect 11152 16118 11204 16124
rect 11256 16114 11284 16390
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10796 15502 10824 15846
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10968 15428 11020 15434
rect 11072 15416 11100 15982
rect 11244 15972 11296 15978
rect 11244 15914 11296 15920
rect 11256 15706 11284 15914
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11072 15388 11284 15416
rect 10968 15370 11020 15376
rect 10784 15360 10836 15366
rect 10980 15314 11008 15370
rect 10836 15308 11008 15314
rect 10784 15302 11008 15308
rect 10796 15286 11008 15302
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11072 13938 11100 14214
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10980 13734 11008 13806
rect 10968 13728 11020 13734
rect 10968 13670 11020 13676
rect 10980 12866 11008 13670
rect 10888 12850 11192 12866
rect 10876 12844 11204 12850
rect 10928 12838 11152 12844
rect 10876 12786 10928 12792
rect 11152 12786 11204 12792
rect 10888 12442 10916 12786
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10336 10674 10364 11698
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10520 11218 10548 11630
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 10520 10810 10548 11154
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10704 10742 10732 11698
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10704 10606 10732 10678
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10520 8022 10548 8842
rect 10796 8838 10824 9318
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10508 8016 10560 8022
rect 10508 7958 10560 7964
rect 10520 7410 10548 7958
rect 10704 7478 10732 8774
rect 10692 7472 10744 7478
rect 10692 7414 10744 7420
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10796 7342 10824 8774
rect 10888 7886 10916 8910
rect 11164 8906 11192 10406
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 11256 7886 11284 15388
rect 11348 14414 11376 16934
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 16250 11744 16526
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11348 12782 11376 13126
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 10888 7410 10916 7822
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10784 7336 10836 7342
rect 9968 7262 10088 7290
rect 10784 7278 10836 7284
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9968 6798 9996 7142
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 10060 3534 10088 7262
rect 10600 5296 10652 5302
rect 10598 5264 10600 5273
rect 10652 5264 10654 5273
rect 10598 5199 10654 5208
rect 10692 5228 10744 5234
rect 10796 5216 10824 7278
rect 11336 7268 11388 7274
rect 11336 7210 11388 7216
rect 11348 6798 11376 7210
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11072 6322 11100 6598
rect 11164 6322 11192 6734
rect 11348 6322 11376 6734
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 10744 5188 10824 5216
rect 11334 5264 11390 5273
rect 11334 5199 11336 5208
rect 10692 5170 10744 5176
rect 10796 5148 10824 5188
rect 11388 5199 11390 5208
rect 11336 5170 11388 5176
rect 10876 5160 10928 5166
rect 10796 5120 10876 5148
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10704 3602 10732 5034
rect 10796 4758 10824 5120
rect 10876 5102 10928 5108
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 11348 4690 11376 5170
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10796 4146 10824 4558
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11164 4146 11192 4422
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10060 3194 10088 3470
rect 10888 3194 10916 3470
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 8036 2746 8156 2774
rect 8128 2582 8156 2746
rect 9784 2746 9904 2774
rect 8758 2680 8814 2689
rect 8758 2615 8814 2624
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 8206 2544 8262 2553
rect 8206 2479 8262 2488
rect 8220 2446 8248 2479
rect 8772 2446 8800 2615
rect 9784 2446 9812 2746
rect 10336 2446 10364 2790
rect 11348 2446 11376 2790
rect 11440 2514 11468 15302
rect 11520 14544 11572 14550
rect 11520 14486 11572 14492
rect 11532 13938 11560 14486
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11624 13938 11652 14418
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11624 13802 11652 13874
rect 11612 13796 11664 13802
rect 11612 13738 11664 13744
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11624 11830 11652 12038
rect 11612 11824 11664 11830
rect 11612 11766 11664 11772
rect 11808 11626 11836 17070
rect 11900 17066 11928 19200
rect 12256 17604 12308 17610
rect 12256 17546 12308 17552
rect 11888 17060 11940 17066
rect 11888 17002 11940 17008
rect 12268 16794 12296 17546
rect 12452 17202 12480 19200
rect 13004 17338 13032 19200
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 11888 16584 11940 16590
rect 12164 16584 12216 16590
rect 11940 16532 12020 16538
rect 11888 16526 12020 16532
rect 12164 16526 12216 16532
rect 11900 16510 12020 16526
rect 11992 16454 12020 16510
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 12176 16250 12204 16526
rect 12348 16516 12400 16522
rect 12348 16458 12400 16464
rect 12360 16425 12388 16458
rect 12346 16416 12402 16425
rect 12346 16351 12402 16360
rect 12452 16250 12480 17138
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12544 16232 12572 16594
rect 12728 16522 12756 16730
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12544 16204 12756 16232
rect 11992 16114 12480 16130
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11980 16108 12492 16114
rect 12032 16102 12440 16108
rect 11980 16050 12032 16056
rect 12440 16050 12492 16056
rect 11900 15638 11928 16050
rect 11888 15632 11940 15638
rect 11888 15574 11940 15580
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11992 10606 12020 15506
rect 12452 15502 12480 16050
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 12544 15434 12572 16204
rect 12728 16114 12756 16204
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12636 15570 12664 16050
rect 12820 15994 12848 17070
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12728 15966 12848 15994
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 12360 14278 12388 14758
rect 12728 14634 12756 15966
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12820 15162 12848 15846
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12912 15026 12940 16934
rect 13004 16522 13216 16538
rect 13004 16516 13228 16522
rect 13004 16510 13176 16516
rect 13004 16454 13032 16510
rect 13176 16458 13228 16464
rect 12992 16448 13044 16454
rect 13084 16448 13136 16454
rect 12992 16390 13044 16396
rect 13082 16416 13084 16425
rect 13136 16416 13138 16425
rect 13082 16351 13138 16360
rect 13096 15978 13124 16351
rect 13188 16114 13216 16458
rect 13280 16250 13308 17138
rect 13556 16522 13584 19200
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 13912 17196 13964 17202
rect 14016 17184 14044 17274
rect 14108 17202 14136 19200
rect 14660 17202 14688 19200
rect 15016 17740 15068 17746
rect 15016 17682 15068 17688
rect 13964 17156 14044 17184
rect 13912 17138 13964 17144
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13372 16182 13400 16390
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13084 15972 13136 15978
rect 13084 15914 13136 15920
rect 13464 15722 13492 16390
rect 13924 16114 13952 16934
rect 14016 16250 14044 17156
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14004 16244 14056 16250
rect 14004 16186 14056 16192
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 13372 15694 13492 15722
rect 13740 15706 13768 15846
rect 13728 15700 13780 15706
rect 13004 15366 13032 15642
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12636 14606 12756 14634
rect 12636 14550 12664 14606
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12256 13864 12308 13870
rect 12360 13852 12388 14214
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12452 13870 12480 14010
rect 12544 13938 12572 14214
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12308 13824 12388 13852
rect 12440 13864 12492 13870
rect 12256 13806 12308 13812
rect 12440 13806 12492 13812
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12268 12170 12296 12582
rect 12452 12434 12480 13806
rect 12636 13802 12664 14350
rect 12728 13870 12756 14606
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12624 13796 12676 13802
rect 12624 13738 12676 13744
rect 12912 13394 12940 14962
rect 13004 14414 13032 15302
rect 13096 14618 13124 15438
rect 13372 15434 13400 15694
rect 13728 15642 13780 15648
rect 13452 15632 13504 15638
rect 13452 15574 13504 15580
rect 13820 15632 13872 15638
rect 13820 15574 13872 15580
rect 13360 15428 13412 15434
rect 13360 15370 13412 15376
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 13004 13394 13032 13874
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 13004 12918 13032 13330
rect 13372 13326 13400 15370
rect 13464 15026 13492 15574
rect 13832 15026 13860 15574
rect 14476 15502 14504 17070
rect 15028 17066 15056 17682
rect 15212 17338 15240 19200
rect 15764 17542 15792 19200
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15016 17060 15068 17066
rect 15016 17002 15068 17008
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14660 16794 14688 16934
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 15120 16726 15148 17138
rect 15292 17060 15344 17066
rect 15292 17002 15344 17008
rect 15304 16794 15332 17002
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 15108 16720 15160 16726
rect 15108 16662 15160 16668
rect 14740 16516 14792 16522
rect 14740 16458 14792 16464
rect 15108 16516 15160 16522
rect 15108 16458 15160 16464
rect 14752 16289 14780 16458
rect 14738 16280 14794 16289
rect 15120 16250 15148 16458
rect 14738 16215 14794 16224
rect 15108 16244 15160 16250
rect 15160 16204 15240 16232
rect 15108 16186 15160 16192
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13636 14408 13688 14414
rect 13636 14350 13688 14356
rect 13648 13938 13676 14350
rect 14188 14340 14240 14346
rect 14188 14282 14240 14288
rect 14372 14340 14424 14346
rect 14372 14282 14424 14288
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 12992 12912 13044 12918
rect 12992 12854 13044 12860
rect 12452 12406 12572 12434
rect 12544 12238 12572 12406
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12256 12164 12308 12170
rect 12256 12106 12308 12112
rect 12544 11898 12572 12174
rect 13004 12102 13032 12854
rect 13648 12646 13676 13874
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 14016 13394 14044 13670
rect 14200 13530 14228 14282
rect 14384 13870 14412 14282
rect 14476 13938 14504 15438
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14280 13796 14332 13802
rect 14280 13738 14332 13744
rect 14292 13530 14320 13738
rect 14384 13530 14412 13806
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 14188 13252 14240 13258
rect 14292 13240 14320 13466
rect 14568 13258 14596 16050
rect 15212 15570 15240 16204
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 15304 15094 15332 16730
rect 15396 16590 15424 17478
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 16040 17202 16068 17274
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15396 15502 15424 16526
rect 15580 16522 15608 16934
rect 15672 16794 15700 17138
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15568 16516 15620 16522
rect 15568 16458 15620 16464
rect 15580 15502 15608 16458
rect 15672 16250 15700 16730
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15764 15978 15792 17138
rect 15948 16436 15976 17138
rect 16212 17128 16264 17134
rect 16118 17096 16174 17105
rect 16212 17070 16264 17076
rect 16118 17031 16174 17040
rect 16132 16998 16160 17031
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 16120 16992 16172 16998
rect 16120 16934 16172 16940
rect 16040 16658 16068 16934
rect 16224 16726 16252 17070
rect 16212 16720 16264 16726
rect 16212 16662 16264 16668
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 16316 16454 16344 19200
rect 16764 17604 16816 17610
rect 16764 17546 16816 17552
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16500 17270 16528 17478
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 16304 16448 16356 16454
rect 15948 16408 16068 16436
rect 16040 16182 16068 16408
rect 16304 16390 16356 16396
rect 16316 16182 16344 16390
rect 16028 16176 16080 16182
rect 16028 16118 16080 16124
rect 16304 16176 16356 16182
rect 16304 16118 16356 16124
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 15752 15972 15804 15978
rect 15752 15914 15804 15920
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 15292 15088 15344 15094
rect 15292 15030 15344 15036
rect 15396 15026 15424 15438
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15304 13938 15332 14758
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15304 13326 15332 13874
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 14240 13212 14320 13240
rect 14556 13252 14608 13258
rect 14188 13194 14240 13200
rect 14556 13194 14608 13200
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13648 12442 13676 12582
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13280 12170 13308 12378
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 13268 12164 13320 12170
rect 13268 12106 13320 12112
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13372 11898 13400 12038
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 14016 11762 14044 12310
rect 14384 12238 14412 12854
rect 14936 12850 14964 12922
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14936 12306 14964 12786
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 15212 11898 15240 13126
rect 15396 12986 15424 14962
rect 15580 14958 15608 15438
rect 15672 15026 15700 15506
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15476 13456 15528 13462
rect 15476 13398 15528 13404
rect 15488 13326 15516 13398
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15396 12850 15424 12922
rect 15580 12918 15608 14894
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15672 13326 15700 13466
rect 15764 13326 15792 13942
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15948 12918 15976 15982
rect 16040 15910 16068 16118
rect 16500 16114 16528 17206
rect 16776 17202 16804 17546
rect 16868 17338 16896 19200
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16592 16250 16620 16526
rect 16684 16522 16712 16934
rect 16776 16794 16804 17138
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16672 16516 16724 16522
rect 16672 16458 16724 16464
rect 16764 16516 16816 16522
rect 16764 16458 16816 16464
rect 16580 16244 16632 16250
rect 16580 16186 16632 16192
rect 16488 16108 16540 16114
rect 16488 16050 16540 16056
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 16028 15904 16080 15910
rect 16028 15846 16080 15852
rect 16028 15564 16080 15570
rect 16028 15506 16080 15512
rect 16040 13938 16068 15506
rect 16592 15502 16620 15914
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16132 15094 16160 15438
rect 16120 15088 16172 15094
rect 16120 15030 16172 15036
rect 16396 14408 16448 14414
rect 16396 14350 16448 14356
rect 16212 14340 16264 14346
rect 16212 14282 16264 14288
rect 16224 13938 16252 14282
rect 16408 14006 16436 14350
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 16040 13462 16068 13874
rect 16224 13462 16252 13874
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 16040 13326 16068 13398
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15384 12164 15436 12170
rect 15384 12106 15436 12112
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15304 11898 15332 12038
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15304 11762 15332 11834
rect 15396 11762 15424 12106
rect 15672 11762 15700 12582
rect 15764 11762 15792 12582
rect 16500 12306 16528 13806
rect 16580 13796 16632 13802
rect 16580 13738 16632 13744
rect 16488 12300 16540 12306
rect 16488 12242 16540 12248
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 14016 11082 14044 11698
rect 14200 11150 14228 11698
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14648 11620 14700 11626
rect 14648 11562 14700 11568
rect 14660 11354 14688 11562
rect 14844 11354 14872 11630
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 15304 11150 15332 11698
rect 15396 11558 15424 11698
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15396 11150 15424 11494
rect 15672 11286 15700 11698
rect 15660 11280 15712 11286
rect 15660 11222 15712 11228
rect 15764 11218 15792 11698
rect 16408 11558 16436 11698
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 14004 11076 14056 11082
rect 14004 11018 14056 11024
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12820 10674 12848 10950
rect 13464 10810 13492 11018
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 14016 10674 14044 11018
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 11992 9994 12020 10542
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12544 10198 12572 10406
rect 13004 10266 13032 10610
rect 13188 10538 13216 10610
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 13188 10266 13216 10474
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 15212 10130 15240 11018
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15304 10062 15332 10406
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11900 8974 11928 9522
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 12360 8838 12388 9318
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12360 8430 12388 8774
rect 12452 8634 12480 9114
rect 13556 8974 13584 9862
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12452 8498 12480 8570
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 11716 7410 11744 8298
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11624 6322 11652 6734
rect 11808 6662 11836 7278
rect 12176 6798 12204 8366
rect 12992 8356 13044 8362
rect 12992 8298 13044 8304
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12268 7342 12296 8230
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12164 6792 12216 6798
rect 12164 6734 12216 6740
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11808 6322 11836 6598
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11796 6316 11848 6322
rect 12176 6304 12204 6734
rect 12268 6662 12296 7278
rect 12360 6866 12388 7482
rect 12912 6866 12940 7482
rect 13004 6866 13032 8298
rect 13832 7410 13860 9114
rect 14188 8900 14240 8906
rect 14188 8842 14240 8848
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13924 7478 13952 8774
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 13912 7472 13964 7478
rect 13912 7414 13964 7420
rect 14108 7410 14136 8502
rect 14200 7410 14228 8842
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 14648 7472 14700 7478
rect 14648 7414 14700 7420
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 13096 6322 13124 7142
rect 13832 7002 13860 7346
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13924 6866 13952 7278
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13372 6322 13400 6598
rect 12256 6316 12308 6322
rect 12176 6276 12256 6304
rect 11796 6258 11848 6264
rect 12256 6258 12308 6264
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 12440 6180 12492 6186
rect 12440 6122 12492 6128
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 11520 5840 11572 5846
rect 11520 5782 11572 5788
rect 11532 5234 11560 5782
rect 12084 5710 12112 6054
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 12164 5636 12216 5642
rect 12164 5578 12216 5584
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 12176 3738 12204 5578
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12360 4554 12388 5170
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11900 3194 11928 3538
rect 12360 3534 12388 4082
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12360 3194 12388 3470
rect 12452 3194 12480 6122
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12544 5216 12572 6054
rect 13556 5914 13584 6258
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12636 5370 12664 5646
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12544 5188 12664 5216
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12544 4690 12572 5034
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12636 4298 12664 5188
rect 12544 4270 12664 4298
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12544 3126 12572 4270
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12636 3602 12664 4082
rect 12728 4010 12756 5646
rect 12820 5302 12848 5646
rect 12808 5296 12860 5302
rect 12808 5238 12860 5244
rect 12900 5296 12952 5302
rect 12900 5238 12952 5244
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12820 4622 12848 5102
rect 12912 5098 12940 5238
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 12900 5092 12952 5098
rect 12900 5034 12952 5040
rect 13096 5030 13124 5170
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 13176 5024 13228 5030
rect 13176 4966 13228 4972
rect 13096 4622 13124 4966
rect 13188 4622 13216 4966
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 12716 4004 12768 4010
rect 12716 3946 12768 3952
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12912 3126 12940 4422
rect 13096 3194 13124 4422
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12900 3120 12952 3126
rect 12900 3062 12952 3068
rect 12532 2916 12584 2922
rect 12532 2858 12584 2864
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 11532 2446 11560 2790
rect 12544 2446 12572 2858
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12636 2446 12664 2790
rect 13648 2446 13676 6598
rect 14108 6390 14136 7346
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 14108 4622 14136 6326
rect 14200 6254 14228 7346
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14292 6798 14320 7142
rect 14660 6798 14688 7414
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14384 6458 14412 6734
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14200 5234 14228 6190
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14568 4690 14596 4966
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 14108 2446 14136 4422
rect 14660 2446 14688 6598
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14752 2990 14780 4626
rect 15120 4622 15148 7482
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 11336 2440 11388 2446
rect 11336 2382 11388 2388
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 6920 2372 6972 2378
rect 6920 2314 6972 2320
rect 7472 2372 7524 2378
rect 7472 2314 7524 2320
rect 8024 2372 8076 2378
rect 8024 2314 8076 2320
rect 8576 2372 8628 2378
rect 8576 2314 8628 2320
rect 9128 2372 9180 2378
rect 9128 2314 9180 2320
rect 10784 2372 10836 2378
rect 10784 2314 10836 2320
rect 11888 2372 11940 2378
rect 11888 2314 11940 2320
rect 12440 2372 12492 2378
rect 12440 2314 12492 2320
rect 12992 2372 13044 2378
rect 12992 2314 13044 2320
rect 13544 2372 13596 2378
rect 13544 2314 13596 2320
rect 6932 800 6960 2314
rect 7484 800 7512 2314
rect 8036 800 8064 2314
rect 8588 800 8616 2314
rect 9140 800 9168 2314
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 9692 800 9720 2246
rect 10244 800 10272 2246
rect 10796 800 10824 2314
rect 11336 2304 11388 2310
rect 11336 2246 11388 2252
rect 11348 800 11376 2246
rect 11900 800 11928 2314
rect 12452 800 12480 2314
rect 13004 800 13032 2314
rect 13556 800 13584 2314
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 14108 800 14136 2246
rect 14752 1170 14780 2450
rect 15580 2446 15608 10134
rect 15764 10062 15792 10542
rect 16592 10538 16620 13738
rect 16776 10674 16804 16458
rect 16868 16250 16896 17274
rect 17420 16674 17448 19200
rect 17420 16646 17540 16674
rect 17512 16590 17540 16646
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 16856 16244 16908 16250
rect 16856 16186 16908 16192
rect 17236 16046 17264 16390
rect 17512 16250 17540 16526
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 16948 14272 17000 14278
rect 16948 14214 17000 14220
rect 16960 14074 16988 14214
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17052 13530 17080 13874
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 17144 12238 17172 15302
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17316 13796 17368 13802
rect 17316 13738 17368 13744
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17144 11898 17172 12174
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 16868 11286 16896 11630
rect 16948 11620 17000 11626
rect 16948 11562 17000 11568
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16960 10674 16988 11562
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16580 10532 16632 10538
rect 16580 10474 16632 10480
rect 16592 10062 16620 10474
rect 16672 10192 16724 10198
rect 16672 10134 16724 10140
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 15752 2508 15804 2514
rect 15752 2450 15804 2456
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 14660 1142 14780 1170
rect 14660 800 14688 1142
rect 15212 800 15240 2246
rect 15764 800 15792 2450
rect 16224 2446 16252 9862
rect 16684 2446 16712 10134
rect 16776 9994 16804 10610
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16868 10062 16896 10542
rect 16960 10130 16988 10610
rect 17132 10532 17184 10538
rect 17132 10474 17184 10480
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16764 9988 16816 9994
rect 16764 9930 16816 9936
rect 16776 9654 16804 9930
rect 16868 9722 16896 9998
rect 16948 9988 17000 9994
rect 16948 9930 17000 9936
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16764 9648 16816 9654
rect 16960 9602 16988 9930
rect 16764 9590 16816 9596
rect 16868 9586 16988 9602
rect 17144 9586 17172 10474
rect 16856 9580 16988 9586
rect 16908 9574 16988 9580
rect 17132 9580 17184 9586
rect 16856 9522 16908 9528
rect 17132 9522 17184 9528
rect 17236 2446 17264 11494
rect 17328 10810 17356 13738
rect 17512 12434 17540 14418
rect 17684 14068 17736 14074
rect 17684 14010 17736 14016
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17420 12406 17540 12434
rect 17420 11694 17448 12406
rect 17604 12238 17632 13126
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17408 11688 17460 11694
rect 17408 11630 17460 11636
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17420 10062 17448 11630
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17512 3534 17540 9318
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17604 3058 17632 10950
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 16304 2372 16356 2378
rect 16304 2314 16356 2320
rect 16316 800 16344 2314
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 16868 800 16896 2246
rect 17420 800 17448 2926
rect 17696 2774 17724 14010
rect 17788 13802 17816 16526
rect 17972 16250 18000 19200
rect 18326 17232 18382 17241
rect 18524 17202 18552 19200
rect 18326 17167 18382 17176
rect 18512 17196 18564 17202
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 18064 14498 18092 16662
rect 18340 16590 18368 17167
rect 18512 17138 18564 17144
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 18524 16250 18552 17138
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 17972 14470 18092 14498
rect 17776 13796 17828 13802
rect 17776 13738 17828 13744
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17880 13326 17908 13670
rect 17868 13320 17920 13326
rect 17868 13262 17920 13268
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17788 11762 17816 12038
rect 17880 11898 17908 12038
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17880 11150 17908 11834
rect 17972 11830 18000 14470
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17972 9926 18000 11766
rect 18064 11218 18092 13330
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18156 11370 18184 12786
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18340 12345 18368 12718
rect 18326 12336 18382 12345
rect 18326 12271 18382 12280
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 18248 11762 18276 12038
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 18156 11342 18276 11370
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 18156 10470 18184 11154
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 18156 9994 18184 10406
rect 18144 9988 18196 9994
rect 18144 9930 18196 9936
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17972 9450 18000 9862
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 18248 7546 18276 11342
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18328 7812 18380 7818
rect 18328 7754 18380 7760
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18340 7449 18368 7754
rect 18326 7440 18382 7449
rect 18326 7375 18382 7384
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18064 3534 18092 3878
rect 18420 3596 18472 3602
rect 18420 3538 18472 3544
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 18328 3460 18380 3466
rect 18328 3402 18380 3408
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 17696 2746 17816 2774
rect 17788 2446 17816 2746
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17972 800 18000 2926
rect 18340 2553 18368 3402
rect 18326 2544 18382 2553
rect 18326 2479 18382 2488
rect 18432 1714 18460 3538
rect 18524 3058 18552 9862
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18432 1686 18552 1714
rect 18524 800 18552 1686
rect 1398 0 1454 800
rect 1950 0 2006 800
rect 2502 0 2558 800
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4158 0 4214 800
rect 4710 0 4766 800
rect 5262 0 5318 800
rect 5814 0 5870 800
rect 6366 0 6422 800
rect 6918 0 6974 800
rect 7470 0 7526 800
rect 8022 0 8078 800
rect 8574 0 8630 800
rect 9126 0 9182 800
rect 9678 0 9734 800
rect 10230 0 10286 800
rect 10782 0 10838 800
rect 11334 0 11390 800
rect 11886 0 11942 800
rect 12438 0 12494 800
rect 12990 0 13046 800
rect 13542 0 13598 800
rect 14094 0 14150 800
rect 14646 0 14702 800
rect 15198 0 15254 800
rect 15750 0 15806 800
rect 16302 0 16358 800
rect 16854 0 16910 800
rect 17406 0 17462 800
rect 17958 0 18014 800
rect 18510 0 18566 800
<< via2 >>
rect 1398 17992 1454 18048
rect 1306 16904 1362 16960
rect 1306 15816 1362 15872
rect 1306 14728 1362 14784
rect 1306 13640 1362 13696
rect 1306 12552 1362 12608
rect 1306 11464 1362 11520
rect 1306 10376 1362 10432
rect 1306 9288 1362 9344
rect 1122 8200 1178 8256
rect 1306 7112 1362 7168
rect 1306 6024 1362 6080
rect 1306 4936 1362 4992
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 1306 3848 1362 3904
rect 1306 2760 1362 2816
rect 1214 1672 1270 1728
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 5170 8880 5226 8936
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 5446 8880 5502 8936
rect 5630 8744 5686 8800
rect 6182 8744 6238 8800
rect 11702 17076 11704 17096
rect 11704 17076 11756 17096
rect 11756 17076 11758 17096
rect 11702 17040 11758 17076
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 8758 15272 8814 15328
rect 8942 13776 8998 13832
rect 11150 16224 11206 16280
rect 10598 5244 10600 5264
rect 10600 5244 10652 5264
rect 10652 5244 10654 5264
rect 10598 5208 10654 5244
rect 11334 5228 11390 5264
rect 11334 5208 11336 5228
rect 11336 5208 11388 5228
rect 11388 5208 11390 5228
rect 8758 2624 8814 2680
rect 8206 2488 8262 2544
rect 12346 16360 12402 16416
rect 13082 16396 13084 16416
rect 13084 16396 13136 16416
rect 13136 16396 13138 16416
rect 13082 16360 13138 16396
rect 14738 16224 14794 16280
rect 16118 17040 16174 17096
rect 18326 17176 18382 17232
rect 18326 12280 18382 12336
rect 18326 7384 18382 7440
rect 18326 2488 18382 2544
<< metal3 >>
rect 0 18050 800 18080
rect 1393 18050 1459 18053
rect 0 18048 1459 18050
rect 0 17992 1398 18048
rect 1454 17992 1459 18048
rect 0 17990 1459 17992
rect 0 17960 800 17990
rect 1393 17987 1459 17990
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 18321 17234 18387 17237
rect 19200 17234 20000 17264
rect 18321 17232 20000 17234
rect 18321 17176 18326 17232
rect 18382 17176 20000 17232
rect 18321 17174 20000 17176
rect 18321 17171 18387 17174
rect 19200 17144 20000 17174
rect 11697 17098 11763 17101
rect 16113 17098 16179 17101
rect 11697 17096 16179 17098
rect 11697 17040 11702 17096
rect 11758 17040 16118 17096
rect 16174 17040 16179 17096
rect 11697 17038 16179 17040
rect 11697 17035 11763 17038
rect 16113 17035 16179 17038
rect 0 16962 800 16992
rect 1301 16962 1367 16965
rect 0 16960 1367 16962
rect 0 16904 1306 16960
rect 1362 16904 1367 16960
rect 0 16902 1367 16904
rect 0 16872 800 16902
rect 1301 16899 1367 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 12341 16418 12407 16421
rect 13077 16418 13143 16421
rect 12341 16416 13143 16418
rect 12341 16360 12346 16416
rect 12402 16360 13082 16416
rect 13138 16360 13143 16416
rect 12341 16358 13143 16360
rect 12341 16355 12407 16358
rect 13077 16355 13143 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 11145 16282 11211 16285
rect 14733 16282 14799 16285
rect 11145 16280 14799 16282
rect 11145 16224 11150 16280
rect 11206 16224 14738 16280
rect 14794 16224 14799 16280
rect 11145 16222 14799 16224
rect 11145 16219 11211 16222
rect 14733 16219 14799 16222
rect 0 15874 800 15904
rect 1301 15874 1367 15877
rect 0 15872 1367 15874
rect 0 15816 1306 15872
rect 1362 15816 1367 15872
rect 0 15814 1367 15816
rect 0 15784 800 15814
rect 1301 15811 1367 15814
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 8753 15330 8819 15333
rect 8886 15330 8892 15332
rect 8753 15328 8892 15330
rect 8753 15272 8758 15328
rect 8814 15272 8892 15328
rect 8753 15270 8892 15272
rect 8753 15267 8819 15270
rect 8886 15268 8892 15270
rect 8956 15268 8962 15332
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 0 14786 800 14816
rect 1301 14786 1367 14789
rect 0 14784 1367 14786
rect 0 14728 1306 14784
rect 1362 14728 1367 14784
rect 0 14726 1367 14728
rect 0 14696 800 14726
rect 1301 14723 1367 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 8937 13834 9003 13837
rect 9070 13834 9076 13836
rect 8937 13832 9076 13834
rect 8937 13776 8942 13832
rect 8998 13776 9076 13832
rect 8937 13774 9076 13776
rect 8937 13771 9003 13774
rect 9070 13772 9076 13774
rect 9140 13772 9146 13836
rect 0 13698 800 13728
rect 1301 13698 1367 13701
rect 0 13696 1367 13698
rect 0 13640 1306 13696
rect 1362 13640 1367 13696
rect 0 13638 1367 13640
rect 0 13608 800 13638
rect 1301 13635 1367 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 0 12610 800 12640
rect 1301 12610 1367 12613
rect 0 12608 1367 12610
rect 0 12552 1306 12608
rect 1362 12552 1367 12608
rect 0 12550 1367 12552
rect 0 12520 800 12550
rect 1301 12547 1367 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 18321 12338 18387 12341
rect 19200 12338 20000 12368
rect 18321 12336 20000 12338
rect 18321 12280 18326 12336
rect 18382 12280 20000 12336
rect 18321 12278 20000 12280
rect 18321 12275 18387 12278
rect 19200 12248 20000 12278
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 0 11522 800 11552
rect 1301 11522 1367 11525
rect 0 11520 1367 11522
rect 0 11464 1306 11520
rect 1362 11464 1367 11520
rect 0 11462 1367 11464
rect 0 11432 800 11462
rect 1301 11459 1367 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 0 10434 800 10464
rect 1301 10434 1367 10437
rect 0 10432 1367 10434
rect 0 10376 1306 10432
rect 1362 10376 1367 10432
rect 0 10374 1367 10376
rect 0 10344 800 10374
rect 1301 10371 1367 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 0 9346 800 9376
rect 1301 9346 1367 9349
rect 0 9344 1367 9346
rect 0 9288 1306 9344
rect 1362 9288 1367 9344
rect 0 9286 1367 9288
rect 0 9256 800 9286
rect 1301 9283 1367 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 5165 8938 5231 8941
rect 5441 8938 5507 8941
rect 5165 8936 5507 8938
rect 5165 8880 5170 8936
rect 5226 8880 5446 8936
rect 5502 8880 5507 8936
rect 5165 8878 5507 8880
rect 5165 8875 5231 8878
rect 5441 8875 5507 8878
rect 5625 8802 5691 8805
rect 6177 8802 6243 8805
rect 5625 8800 6243 8802
rect 5625 8744 5630 8800
rect 5686 8744 6182 8800
rect 6238 8744 6243 8800
rect 5625 8742 6243 8744
rect 5625 8739 5691 8742
rect 6177 8739 6243 8742
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 0 8258 800 8288
rect 1117 8258 1183 8261
rect 0 8256 1183 8258
rect 0 8200 1122 8256
rect 1178 8200 1183 8256
rect 0 8198 1183 8200
rect 0 8168 800 8198
rect 1117 8195 1183 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 18321 7442 18387 7445
rect 19200 7442 20000 7472
rect 18321 7440 20000 7442
rect 18321 7384 18326 7440
rect 18382 7384 20000 7440
rect 18321 7382 20000 7384
rect 18321 7379 18387 7382
rect 19200 7352 20000 7382
rect 0 7170 800 7200
rect 1301 7170 1367 7173
rect 0 7168 1367 7170
rect 0 7112 1306 7168
rect 1362 7112 1367 7168
rect 0 7110 1367 7112
rect 0 7080 800 7110
rect 1301 7107 1367 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 0 6082 800 6112
rect 1301 6082 1367 6085
rect 0 6080 1367 6082
rect 0 6024 1306 6080
rect 1362 6024 1367 6080
rect 0 6022 1367 6024
rect 0 5992 800 6022
rect 1301 6019 1367 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 10593 5266 10659 5269
rect 11329 5266 11395 5269
rect 10593 5264 11395 5266
rect 10593 5208 10598 5264
rect 10654 5208 11334 5264
rect 11390 5208 11395 5264
rect 10593 5206 11395 5208
rect 10593 5203 10659 5206
rect 11329 5203 11395 5206
rect 0 4994 800 5024
rect 1301 4994 1367 4997
rect 0 4992 1367 4994
rect 0 4936 1306 4992
rect 1362 4936 1367 4992
rect 0 4934 1367 4936
rect 0 4904 800 4934
rect 1301 4931 1367 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 0 3906 800 3936
rect 1301 3906 1367 3909
rect 0 3904 1367 3906
rect 0 3848 1306 3904
rect 1362 3848 1367 3904
rect 0 3846 1367 3848
rect 0 3816 800 3846
rect 1301 3843 1367 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 0 2818 800 2848
rect 1301 2818 1367 2821
rect 0 2816 1367 2818
rect 0 2760 1306 2816
rect 1362 2760 1367 2816
rect 0 2758 1367 2760
rect 0 2728 800 2758
rect 1301 2755 1367 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 8753 2682 8819 2685
rect 8886 2682 8892 2684
rect 8753 2680 8892 2682
rect 8753 2624 8758 2680
rect 8814 2624 8892 2680
rect 8753 2622 8892 2624
rect 8753 2619 8819 2622
rect 8886 2620 8892 2622
rect 8956 2620 8962 2684
rect 8201 2546 8267 2549
rect 9070 2546 9076 2548
rect 8201 2544 9076 2546
rect 8201 2488 8206 2544
rect 8262 2488 9076 2544
rect 8201 2486 9076 2488
rect 8201 2483 8267 2486
rect 9070 2484 9076 2486
rect 9140 2484 9146 2548
rect 18321 2546 18387 2549
rect 19200 2546 20000 2576
rect 18321 2544 20000 2546
rect 18321 2488 18326 2544
rect 18382 2488 20000 2544
rect 18321 2486 20000 2488
rect 18321 2483 18387 2486
rect 19200 2456 20000 2486
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 0 1730 800 1760
rect 1209 1730 1275 1733
rect 0 1728 1275 1730
rect 0 1672 1214 1728
rect 1270 1672 1275 1728
rect 0 1670 1275 1672
rect 0 1640 800 1670
rect 1209 1667 1275 1670
<< via3 >>
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 8892 15268 8956 15332
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 9076 13772 9140 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 8892 2620 8956 2684
rect 9076 2484 9140 2548
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 16896 4528 17456
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 17440 5188 17456
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 8891 15332 8957 15333
rect 8891 15268 8892 15332
rect 8956 15268 8957 15332
rect 8891 15267 8957 15268
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 8894 2685 8954 15267
rect 9075 13836 9141 13837
rect 9075 13772 9076 13836
rect 9140 13772 9141 13836
rect 9075 13771 9141 13772
rect 8891 2684 8957 2685
rect 8891 2620 8892 2684
rect 8956 2620 8957 2684
rect 8891 2619 8957 2620
rect 9078 2549 9138 13771
rect 9075 2548 9141 2549
rect 9075 2484 9076 2548
rect 9140 2484 9141 2548
rect 9075 2483 9141 2484
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _227_
timestamp -25199
transform -1 0 11960 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp -25199
transform 1 0 8740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp -25199
transform 1 0 9016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _230_
timestamp -25199
transform 1 0 11224 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp -25199
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _232_
timestamp -25199
transform -1 0 5888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _233_
timestamp -25199
transform -1 0 7084 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _234_
timestamp -25199
transform 1 0 5244 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _235_
timestamp -25199
transform 1 0 6624 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__nand3_1  _236_
timestamp -25199
transform 1 0 15456 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _237_
timestamp -25199
transform -1 0 15456 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _238_
timestamp -25199
transform 1 0 15732 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _239_
timestamp -25199
transform 1 0 9660 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _240_
timestamp -25199
transform 1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _241_
timestamp -25199
transform 1 0 8924 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _242_
timestamp -25199
transform -1 0 10764 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _243_
timestamp -25199
transform 1 0 13156 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _244_
timestamp -25199
transform -1 0 12512 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _245_
timestamp -25199
transform -1 0 16468 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _246_
timestamp -25199
transform 1 0 14996 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _247_
timestamp -25199
transform 1 0 12512 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp -25199
transform 1 0 14168 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _249_
timestamp -25199
transform 1 0 11040 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _250_
timestamp -25199
transform 1 0 6716 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _251_
timestamp -25199
transform 1 0 6440 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _252_
timestamp -25199
transform 1 0 10212 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _253_
timestamp -25199
transform 1 0 12512 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _254_
timestamp -25199
transform 1 0 12144 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _255_
timestamp -25199
transform 1 0 11500 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _256_
timestamp -25199
transform -1 0 13432 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _257_
timestamp -25199
transform 1 0 13432 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _258_
timestamp -25199
transform -1 0 14260 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _259_
timestamp -25199
transform 1 0 14904 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_2  _260_
timestamp -25199
transform 1 0 15272 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _261_
timestamp -25199
transform 1 0 15272 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _262_
timestamp -25199
transform 1 0 16192 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _263_
timestamp -25199
transform 1 0 13340 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_2  _264_
timestamp -25199
transform 1 0 12420 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _265_
timestamp -25199
transform 1 0 16376 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _266_
timestamp -25199
transform 1 0 15180 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _267_
timestamp -25199
transform 1 0 14812 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _268_
timestamp -25199
transform -1 0 14996 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _269_
timestamp -25199
transform 1 0 17664 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _270_
timestamp -25199
transform 1 0 17020 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _271_
timestamp -25199
transform 1 0 16560 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _272_
timestamp -25199
transform -1 0 16560 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _273_
timestamp -25199
transform -1 0 17664 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _274_
timestamp -25199
transform 1 0 15456 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _275_
timestamp -25199
transform -1 0 16008 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _276_
timestamp -25199
transform -1 0 17204 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _277_
timestamp -25199
transform 1 0 14076 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _278_
timestamp -25199
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _279_
timestamp -25199
transform 1 0 14168 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp -25199
transform 1 0 17296 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _281_
timestamp -25199
transform 1 0 17664 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _282_
timestamp -25199
transform -1 0 18308 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_2  _283_
timestamp -25199
transform 1 0 15732 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp -25199
transform 1 0 17296 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _285_
timestamp -25199
transform 1 0 14076 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _286_
timestamp -25199
transform -1 0 17296 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _287_
timestamp -25199
transform -1 0 17296 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _288_
timestamp -25199
transform 1 0 17756 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _289_
timestamp -25199
transform -1 0 14904 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _290_
timestamp -25199
transform -1 0 17112 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_1  _291_
timestamp -25199
transform -1 0 16284 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _292_
timestamp -25199
transform -1 0 15732 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _293_
timestamp -25199
transform -1 0 17480 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _294_
timestamp -25199
transform -1 0 17480 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _295_
timestamp -25199
transform 1 0 17572 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _296_
timestamp -25199
transform -1 0 18400 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _297_
timestamp -25199
transform 1 0 17572 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _298_
timestamp -25199
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _299_
timestamp -25199
transform 1 0 8004 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _300_
timestamp -25199
transform 1 0 8464 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _301_
timestamp -25199
transform 1 0 7176 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _302_
timestamp -25199
transform 1 0 2116 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _303_
timestamp -25199
transform 1 0 1932 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _304_
timestamp -25199
transform -1 0 8740 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _305_
timestamp -25199
transform 1 0 9016 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _306_
timestamp -25199
transform 1 0 1472 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _307_
timestamp -25199
transform -1 0 3496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _308_
timestamp -25199
transform 1 0 1380 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _309_
timestamp -25199
transform -1 0 2576 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _310_
timestamp -25199
transform 1 0 10580 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _311_
timestamp -25199
transform 1 0 2576 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _312_
timestamp -25199
transform 1 0 2392 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _313_
timestamp -25199
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _314_
timestamp -25199
transform 1 0 8924 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _315_
timestamp -25199
transform 1 0 8188 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _316_
timestamp -25199
transform -1 0 10580 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _317_
timestamp -25199
transform 1 0 11960 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _318_
timestamp -25199
transform 1 0 9200 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _319_
timestamp -25199
transform 1 0 9660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _320_
timestamp -25199
transform -1 0 13248 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _321_
timestamp -25199
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _322_
timestamp -25199
transform -1 0 11040 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _323_
timestamp -25199
transform 1 0 12512 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _324_
timestamp -25199
transform -1 0 13064 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _325_
timestamp -25199
transform -1 0 12696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _326_
timestamp -25199
transform 1 0 13064 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _327_
timestamp -25199
transform 1 0 8924 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_2  _328_
timestamp -25199
transform -1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _329_
timestamp -25199
transform -1 0 10304 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _330_
timestamp -25199
transform 1 0 10948 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _331_
timestamp -25199
transform 1 0 10488 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_2  _332_
timestamp -25199
transform 1 0 10120 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _333_
timestamp -25199
transform 1 0 12144 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _334_
timestamp -25199
transform -1 0 12144 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _335_
timestamp -25199
transform -1 0 13156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _336_
timestamp -25199
transform 1 0 12420 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _337_
timestamp -25199
transform 1 0 11776 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _338_
timestamp -25199
transform 1 0 11500 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _339_
timestamp -25199
transform -1 0 11776 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _340_
timestamp -25199
transform -1 0 12788 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _341_
timestamp -25199
transform 1 0 12788 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _342_
timestamp -25199
transform 1 0 9200 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _343_
timestamp -25199
transform -1 0 9844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _344_
timestamp -25199
transform -1 0 10304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _345_
timestamp -25199
transform 1 0 12236 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _346_
timestamp -25199
transform -1 0 12236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _347_
timestamp -25199
transform 1 0 12880 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp -25199
transform 1 0 13984 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _349_
timestamp -25199
transform 1 0 12972 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _350_
timestamp -25199
transform 1 0 13340 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _351_
timestamp -25199
transform 1 0 9660 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _352_
timestamp -25199
transform 1 0 13800 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _353_
timestamp -25199
transform 1 0 14076 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _354_
timestamp -25199
transform -1 0 10488 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp -25199
transform -1 0 11316 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _356_
timestamp -25199
transform 1 0 11500 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp -25199
transform 1 0 13156 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp -25199
transform 1 0 12328 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _359_
timestamp -25199
transform -1 0 13616 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _360_
timestamp -25199
transform 1 0 14076 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _361_
timestamp -25199
transform -1 0 15272 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _362_
timestamp -25199
transform 1 0 5152 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _363_
timestamp -25199
transform 1 0 3956 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _364_
timestamp -25199
transform 1 0 4416 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _365_
timestamp -25199
transform 1 0 4784 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _366_
timestamp -25199
transform 1 0 6348 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _367_
timestamp -25199
transform 1 0 6348 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _368_
timestamp -25199
transform 1 0 3864 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _369_
timestamp -25199
transform 1 0 3220 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _370_
timestamp -25199
transform -1 0 4600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _371_
timestamp -25199
transform -1 0 5428 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _372_
timestamp -25199
transform 1 0 6624 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _373_
timestamp -25199
transform 1 0 4140 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _374_
timestamp -25199
transform 1 0 4784 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _375_
timestamp -25199
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _376_
timestamp -25199
transform 1 0 6072 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _377_
timestamp -25199
transform 1 0 3956 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _378_
timestamp -25199
transform 1 0 3772 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _379_
timestamp -25199
transform 1 0 4508 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _380_
timestamp -25199
transform -1 0 5980 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _381_
timestamp -25199
transform 1 0 6624 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _382_
timestamp -25199
transform -1 0 11316 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _383_
timestamp -25199
transform 1 0 10396 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _384_
timestamp -25199
transform -1 0 9384 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _385_
timestamp -25199
transform -1 0 8832 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _386_
timestamp -25199
transform -1 0 8740 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _387_
timestamp -25199
transform 1 0 9384 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _388_
timestamp -25199
transform 1 0 7912 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _389_
timestamp -25199
transform 1 0 7268 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _390_
timestamp -25199
transform -1 0 8832 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_2  _391_
timestamp -25199
transform 1 0 7912 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _392_
timestamp -25199
transform -1 0 8832 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _393_
timestamp -25199
transform 1 0 12144 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_2  _394_
timestamp -25199
transform -1 0 12420 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _395_
timestamp -25199
transform 1 0 10764 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _396_
timestamp -25199
transform -1 0 10028 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _397_
timestamp -25199
transform 1 0 9752 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _398_
timestamp -25199
transform 1 0 8556 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _399_
timestamp -25199
transform 1 0 8188 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _400_
timestamp -25199
transform -1 0 11224 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _401_
timestamp -25199
transform 1 0 8188 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _402_
timestamp -25199
transform 1 0 9200 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _403_
timestamp -25199
transform -1 0 10120 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _404_
timestamp -25199
transform -1 0 12512 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _405_
timestamp -25199
transform -1 0 13340 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _406_
timestamp -25199
transform -1 0 12972 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp -25199
transform -1 0 12052 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _408_
timestamp -25199
transform 1 0 13432 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _409_
timestamp -25199
transform -1 0 13432 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _410_
timestamp -25199
transform 1 0 13432 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _411_
timestamp -25199
transform 1 0 10028 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _412_
timestamp -25199
transform 1 0 10580 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _413_
timestamp -25199
transform -1 0 13984 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _414_
timestamp -25199
transform -1 0 14720 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _415_
timestamp -25199
transform 1 0 12328 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _416_
timestamp -25199
transform -1 0 12328 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _417_
timestamp -25199
transform -1 0 5888 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _418_
timestamp -25199
transform -1 0 6624 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _419_
timestamp -25199
transform 1 0 6808 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _420_
timestamp -25199
transform 1 0 8096 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _421_
timestamp -25199
transform 1 0 8924 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _422_
timestamp -25199
transform 1 0 8740 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _423_
timestamp -25199
transform 1 0 10488 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _424_
timestamp -25199
transform -1 0 12420 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _425_
timestamp -25199
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _426_
timestamp -25199
transform 1 0 3220 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _427_
timestamp -25199
transform -1 0 4692 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _428_
timestamp -25199
transform 1 0 2484 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _429_
timestamp -25199
transform 1 0 1840 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _430_
timestamp -25199
transform -1 0 4416 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _431_
timestamp -25199
transform -1 0 8188 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _432_
timestamp -25199
transform 1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _433_
timestamp -25199
transform 1 0 1840 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _434_
timestamp -25199
transform 1 0 1380 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _435_
timestamp -25199
transform 1 0 2300 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _436_
timestamp -25199
transform -1 0 6992 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _437_
timestamp -25199
transform -1 0 7084 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _438_
timestamp -25199
transform 1 0 1748 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _439_
timestamp -25199
transform 1 0 2576 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _440_
timestamp -25199
transform -1 0 5060 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _441_
timestamp -25199
transform 1 0 1932 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _442_
timestamp -25199
transform -1 0 2760 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _443_
timestamp -25199
transform 1 0 2760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _444_
timestamp -25199
transform 1 0 3404 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _445_
timestamp -25199
transform 1 0 4232 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _446_
timestamp -25199
transform -1 0 8280 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _447_
timestamp -25199
transform -1 0 5060 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _448_
timestamp -25199
transform -1 0 5520 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _449_
timestamp -25199
transform -1 0 7544 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _450_
timestamp -25199
transform -1 0 7176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _451_
timestamp -25199
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _452_
timestamp -25199
transform -1 0 6440 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _453_
timestamp -25199
transform 1 0 5704 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _454_
timestamp -25199
transform -1 0 7084 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _455_
timestamp -25199
transform 1 0 3772 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_2  _456_
timestamp -25199
transform 1 0 7728 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _457_
timestamp -25199
transform -1 0 5152 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _458_
timestamp -25199
transform -1 0 5612 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _459_
timestamp -25199
transform -1 0 8648 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_2  _460_
timestamp -25199
transform 1 0 6992 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _461_
timestamp -25199
transform 1 0 6992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _462_
timestamp -25199
transform 1 0 6348 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _463_
timestamp -25199
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _464_
timestamp -25199
transform -1 0 8372 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _465_
timestamp -25199
transform -1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _466_
timestamp -25199
transform 1 0 4140 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _467_
timestamp -25199
transform -1 0 6992 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _468_
timestamp -25199
transform -1 0 6900 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _469_
timestamp -25199
transform 1 0 5428 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _470_
timestamp -25199
transform 1 0 4416 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _471_
timestamp -25199
transform -1 0 5244 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _472_
timestamp -25199
transform 1 0 5244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _473_
timestamp -25199
transform -1 0 9384 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _474_
timestamp -25199
transform -1 0 8372 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _475_
timestamp -25199
transform -1 0 8188 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _476_
timestamp -25199
transform -1 0 6256 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _477_
timestamp -25199
transform 1 0 5888 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _478_
timestamp -25199
transform -1 0 8832 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _479_
timestamp -25199
transform 1 0 5060 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _480_
timestamp -25199
transform -1 0 6900 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _481_
timestamp -25199
transform 1 0 6348 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _482_
timestamp -25199
transform 1 0 1840 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _483_
timestamp -25199
transform 1 0 2116 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _484_
timestamp -25199
transform 1 0 4876 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _485_
timestamp -25199
transform 1 0 4968 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _486_
timestamp -25199
transform 1 0 4140 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _487_
timestamp -25199
transform 1 0 4508 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _488_
timestamp -25199
transform -1 0 5060 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _489_
timestamp -25199
transform -1 0 7452 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__304__A1
timestamp -25199
transform 1 0 7912 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__488__S
timestamp -25199
transform 1 0 5060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout85_A
timestamp -25199
transform 1 0 5980 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout86_X
timestamp -25199
transform -1 0 6164 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout111_A
timestamp -25199
transform -1 0 4048 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp -25199
transform -1 0 3128 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp -25199
transform -1 0 1840 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp -25199
transform -1 0 1840 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp -25199
transform -1 0 1840 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp -25199
transform -1 0 1564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp -25199
transform -1 0 2024 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp -25199
transform -1 0 1840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp -25199
transform -1 0 1840 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp -25199
transform -1 0 1840 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp -25199
transform -1 0 1840 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp -25199
transform -1 0 1840 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp -25199
transform -1 0 1840 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp -25199
transform -1 0 1840 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp -25199
transform -1 0 1840 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp -25199
transform -1 0 2392 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp -25199
transform -1 0 1840 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp -25199
transform -1 0 2024 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_X
timestamp -25199
transform 1 0 2024 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp -25199
transform -1 0 2024 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp -25199
transform -1 0 2576 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp -25199
transform -1 0 3128 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp -25199
transform -1 0 3680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp -25199
transform -1 0 4232 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp -25199
transform -1 0 4784 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp -25199
transform -1 0 4784 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp -25199
transform -1 0 5336 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp -25199
transform -1 0 5888 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp -25199
transform -1 0 6624 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp -25199
transform -1 0 7544 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp -25199
transform -1 0 8096 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp -25199
transform -1 0 8648 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp -25199
transform -1 0 8832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp -25199
transform -1 0 9752 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp -25199
transform -1 0 10304 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp -25199
transform -1 0 11132 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp -25199
transform -1 0 10948 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp -25199
transform -1 0 13432 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp -25199
transform -1 0 13156 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp -25199
transform -1 0 14168 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp -25199
transform -1 0 14536 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp -25199
transform -1 0 15640 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp -25199
transform -1 0 15732 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp -25199
transform -1 0 16560 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp -25199
transform -1 0 17664 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp -25199
transform -1 0 17204 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp -25199
transform -1 0 17020 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp -25199
transform -1 0 17480 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp -25199
transform -1 0 18032 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp -25199
transform -1 0 18584 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output49_A
timestamp -25199
transform 1 0 17848 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  fanout85
timestamp -25199
transform -1 0 5704 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout86
timestamp -25199
transform -1 0 5980 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout87
timestamp -25199
transform -1 0 10212 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout88
timestamp -25199
transform -1 0 11776 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout89
timestamp -25199
transform -1 0 15272 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout90
timestamp -25199
transform -1 0 13524 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout91
timestamp -25199
transform -1 0 18308 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout92
timestamp -25199
transform -1 0 9200 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout93
timestamp -25199
transform 1 0 12144 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout94
timestamp -25199
transform -1 0 14904 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout95
timestamp -25199
transform -1 0 17020 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout96
timestamp -25199
transform -1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout97
timestamp -25199
transform -1 0 15364 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout98
timestamp -25199
transform -1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout99
timestamp -25199
transform -1 0 14904 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout100
timestamp -25199
transform -1 0 13984 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout101
timestamp -25199
transform 1 0 12696 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout102
timestamp -25199
transform -1 0 12696 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout103
timestamp -25199
transform 1 0 12788 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout104
timestamp -25199
transform -1 0 11500 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout105
timestamp -25199
transform -1 0 8832 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout106
timestamp -25199
transform -1 0 8004 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout107
timestamp -25199
transform 1 0 7544 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout108
timestamp -25199
transform 1 0 7544 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout109
timestamp -25199
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout110
timestamp -25199
transform -1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout111
timestamp -25199
transform -1 0 4968 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp -25199
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85
timestamp -25199
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -25199
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -25199
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp -25199
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp -25199
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp -25199
transform 1 0 3496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_39
timestamp -25199
transform 1 0 4692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_50
timestamp -25199
transform 1 0 5704 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp -25199
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_64
timestamp -25199
transform 1 0 6992 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_73
timestamp -25199
transform 1 0 7820 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_85
timestamp -25199
transform 1 0 8924 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -25199
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_140
timestamp 1636943256
transform 1 0 13984 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_152
timestamp 1636943256
transform 1 0 15088 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp -25199
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_169
timestamp -25199
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_177
timestamp -25199
transform 1 0 17388 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_20
timestamp -25199
transform 1 0 2944 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_43
timestamp 1636943256
transform 1 0 5060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_55
timestamp 1636943256
transform 1 0 6164 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_67
timestamp -25199
transform 1 0 7268 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_73
timestamp -25199
transform 1 0 7820 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_103
timestamp 1636943256
transform 1 0 10580 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_115
timestamp -25199
transform 1 0 11684 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_124
timestamp 1636943256
transform 1 0 12512 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp -25199
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636943256
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636943256
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636943256
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_177
timestamp -25199
transform 1 0 17388 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp -25199
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_10
timestamp -25199
transform 1 0 2024 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_16
timestamp 1636943256
transform 1 0 2576 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_28
timestamp -25199
transform 1 0 3680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp -25199
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -25199
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_64
timestamp 1636943256
transform 1 0 6992 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_76
timestamp 1636943256
transform 1 0 8096 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_88
timestamp 1636943256
transform 1 0 9200 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_100
timestamp 1636943256
transform 1 0 10304 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp -25199
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_121
timestamp -25199
transform 1 0 12236 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_126
timestamp 1636943256
transform 1 0 12696 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_138
timestamp 1636943256
transform 1 0 13800 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_150
timestamp 1636943256
transform 1 0 14904 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp -25199
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636943256
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_181
timestamp -25199
transform 1 0 17756 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_184
timestamp -25199
transform 1 0 18032 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp -25199
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_22
timestamp -25199
transform 1 0 3128 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636943256
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636943256
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp -25199
transform 1 0 5980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_57
timestamp -25199
transform 1 0 6348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_65
timestamp -25199
transform 1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_73
timestamp -25199
transform 1 0 7820 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -25199
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636943256
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_97
timestamp -25199
transform 1 0 10028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_113
timestamp -25199
transform 1 0 11500 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_121
timestamp -25199
transform 1 0 12236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_132
timestamp -25199
transform 1 0 13248 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_154
timestamp 1636943256
transform 1 0 15272 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_166
timestamp 1636943256
transform 1 0 16376 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_178
timestamp 1636943256
transform 1 0 17480 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_8
timestamp 1636943256
transform 1 0 1840 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_20
timestamp -25199
transform 1 0 2944 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_24
timestamp -25199
transform 1 0 3312 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_32
timestamp -25199
transform 1 0 4048 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_43
timestamp -25199
transform 1 0 5060 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_49
timestamp -25199
transform 1 0 5612 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp -25199
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_60
timestamp -25199
transform 1 0 6624 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_66
timestamp -25199
transform 1 0 7176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_77
timestamp -25199
transform 1 0 8188 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_85
timestamp -25199
transform 1 0 8924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_93
timestamp -25199
transform 1 0 9660 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_101
timestamp -25199
transform 1 0 10396 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp -25199
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_121
timestamp -25199
transform 1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_136
timestamp -25199
transform 1 0 13616 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_143
timestamp 1636943256
transform 1 0 14260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_155
timestamp 1636943256
transform 1 0 15364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -25199
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636943256
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_181
timestamp -25199
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp -25199
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_5
timestamp -25199
transform 1 0 1564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp -25199
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -25199
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp -25199
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_48
timestamp -25199
transform 1 0 5520 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_74
timestamp -25199
transform 1 0 7912 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp -25199
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp -25199
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636943256
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636943256
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_121
timestamp -25199
transform 1 0 12236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_131
timestamp -25199
transform 1 0 13156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp -25199
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636943256
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636943256
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636943256
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636943256
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_189
timestamp -25199
transform 1 0 18492 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_6
timestamp -25199
transform 1 0 1656 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_14
timestamp -25199
transform 1 0 2392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_23
timestamp 1636943256
transform 1 0 3220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_35
timestamp 1636943256
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp -25199
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -25199
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_65
timestamp -25199
transform 1 0 7084 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp -25199
transform 1 0 8280 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_82
timestamp -25199
transform 1 0 8648 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_89
timestamp 1636943256
transform 1 0 9292 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_101
timestamp -25199
transform 1 0 10396 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_123
timestamp -25199
transform 1 0 12420 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_138
timestamp 1636943256
transform 1 0 13800 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_150
timestamp 1636943256
transform 1 0 14904 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_162
timestamp -25199
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636943256
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_181
timestamp -25199
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_189
timestamp -25199
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp -25199
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_14
timestamp 1636943256
transform 1 0 2392 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp -25199
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_29
timestamp -25199
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_42
timestamp 1636943256
transform 1 0 4968 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_54
timestamp 1636943256
transform 1 0 6072 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_66
timestamp -25199
transform 1 0 7176 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_80
timestamp -25199
transform 1 0 8464 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_100
timestamp -25199
transform 1 0 10304 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_116
timestamp -25199
transform 1 0 11776 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_120
timestamp -25199
transform 1 0 12144 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp -25199
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_154
timestamp 1636943256
transform 1 0 15272 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_166
timestamp 1636943256
transform 1 0 16376 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_178
timestamp 1636943256
transform 1 0 17480 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_26
timestamp -25199
transform 1 0 3496 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_34
timestamp -25199
transform 1 0 4232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp -25199
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -25199
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_67
timestamp -25199
transform 1 0 7268 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_75
timestamp -25199
transform 1 0 8004 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_83
timestamp -25199
transform 1 0 8740 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_92
timestamp -25199
transform 1 0 9568 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp -25199
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_120
timestamp -25199
transform 1 0 12144 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_126
timestamp -25199
transform 1 0 12696 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_135
timestamp -25199
transform 1 0 13524 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_145
timestamp 1636943256
transform 1 0 14444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_157
timestamp -25199
transform 1 0 15548 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp -25199
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636943256
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_181
timestamp -25199
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_189
timestamp -25199
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_13
timestamp -25199
transform 1 0 2300 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -25199
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp -25199
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_40
timestamp 1636943256
transform 1 0 4784 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_52
timestamp -25199
transform 1 0 5888 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp -25199
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636943256
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1636943256
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1636943256
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1636943256
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp -25199
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp -25199
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636943256
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1636943256
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1636943256
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_177
timestamp -25199
transform 1 0 17388 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_183
timestamp -25199
transform 1 0 17940 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_16
timestamp 1636943256
transform 1 0 2576 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_28
timestamp -25199
transform 1 0 3680 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_36
timestamp -25199
transform 1 0 4416 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp -25199
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_63
timestamp -25199
transform 1 0 6900 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_69
timestamp -25199
transform 1 0 7452 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_73
timestamp 1636943256
transform 1 0 7820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_85
timestamp -25199
transform 1 0 8924 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_95
timestamp -25199
transform 1 0 9844 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_100
timestamp 1636943256
transform 1 0 10304 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp -25199
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_130
timestamp 1636943256
transform 1 0 13064 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_142
timestamp 1636943256
transform 1 0 14168 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_154
timestamp 1636943256
transform 1 0 15272 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp -25199
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1636943256
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_181
timestamp -25199
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_189
timestamp -25199
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_10
timestamp 1636943256
transform 1 0 2024 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_22
timestamp -25199
transform 1 0 3128 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_40
timestamp -25199
transform 1 0 4784 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_45
timestamp -25199
transform 1 0 5244 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_61
timestamp -25199
transform 1 0 6716 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_69
timestamp -25199
transform 1 0 7452 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp -25199
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp -25199
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_85
timestamp -25199
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_100
timestamp -25199
transform 1 0 10304 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_109
timestamp -25199
transform 1 0 11132 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_126
timestamp -25199
transform 1 0 12696 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1636943256
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1636943256
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1636943256
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1636943256
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp -25199
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp -25199
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_26
timestamp -25199
transform 1 0 3496 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_64
timestamp -25199
transform 1 0 6992 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_72
timestamp -25199
transform 1 0 7728 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_79
timestamp 1636943256
transform 1 0 8372 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_91
timestamp 1636943256
transform 1 0 9476 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_103
timestamp -25199
transform 1 0 10580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp -25199
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp -25199
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp -25199
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_124
timestamp 1636943256
transform 1 0 12512 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_136
timestamp 1636943256
transform 1 0 13616 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_148
timestamp 1636943256
transform 1 0 14720 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp -25199
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_182
timestamp -25199
transform 1 0 17848 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_8
timestamp 1636943256
transform 1 0 1840 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp -25199
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_29
timestamp -25199
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_35
timestamp -25199
transform 1 0 4324 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_48
timestamp -25199
transform 1 0 5520 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_52
timestamp -25199
transform 1 0 5888 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_55
timestamp -25199
transform 1 0 6164 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_69
timestamp -25199
transform 1 0 7452 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_90
timestamp 1636943256
transform 1 0 9384 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_102
timestamp 1636943256
transform 1 0 10488 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_114
timestamp -25199
transform 1 0 11592 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_122
timestamp -25199
transform 1 0 12328 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_130
timestamp -25199
transform 1 0 13064 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp -25199
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_174
timestamp -25199
transform 1 0 17112 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_188
timestamp -25199
transform 1 0 18400 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_8
timestamp 1636943256
transform 1 0 1840 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_20
timestamp 1636943256
transform 1 0 2944 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_32
timestamp -25199
transform 1 0 4048 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_40
timestamp -25199
transform 1 0 4784 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_50
timestamp -25199
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636943256
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_69
timestamp -25199
transform 1 0 7452 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_77
timestamp -25199
transform 1 0 8188 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_84
timestamp 1636943256
transform 1 0 8832 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_96
timestamp -25199
transform 1 0 9936 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp -25199
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_134
timestamp -25199
transform 1 0 13432 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_145
timestamp 1636943256
transform 1 0 14444 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_157
timestamp -25199
transform 1 0 15548 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp -25199
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_176
timestamp -25199
transform 1 0 17296 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp -25199
transform 1 0 17848 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_187
timestamp -25199
transform 1 0 18308 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636943256
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636943256
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp -25199
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636943256
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1636943256
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_53
timestamp -25199
transform 1 0 5980 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_61
timestamp -25199
transform 1 0 6716 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_71
timestamp 1636943256
transform 1 0 7636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp -25199
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_92
timestamp 1636943256
transform 1 0 9568 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_104
timestamp 1636943256
transform 1 0 10672 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_116
timestamp 1636943256
transform 1 0 11776 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_128
timestamp -25199
transform 1 0 12880 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp -25199
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp -25199
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_156
timestamp 1636943256
transform 1 0 15456 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_168
timestamp -25199
transform 1 0 16560 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_176
timestamp -25199
transform 1 0 17296 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_188
timestamp -25199
transform 1 0 18400 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_8
timestamp 1636943256
transform 1 0 1840 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_20
timestamp -25199
transform 1 0 2944 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_38
timestamp 1636943256
transform 1 0 4600 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_50
timestamp -25199
transform 1 0 5704 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_64
timestamp 1636943256
transform 1 0 6992 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_85
timestamp -25199
transform 1 0 8924 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp -25199
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp -25199
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1636943256
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1636943256
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_137
timestamp -25199
transform 1 0 13708 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp -25199
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_187
timestamp -25199
transform 1 0 18308 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636943256
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636943256
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp -25199
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp -25199
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_47
timestamp -25199
transform 1 0 5428 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_67
timestamp 1636943256
transform 1 0 7268 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_93
timestamp 1636943256
transform 1 0 9660 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_105
timestamp -25199
transform 1 0 10764 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_118
timestamp -25199
transform 1 0 11960 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp -25199
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1636943256
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1636943256
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_165
timestamp -25199
transform 1 0 16284 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_173
timestamp -25199
transform 1 0 17020 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_185
timestamp -25199
transform 1 0 18124 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp -25199
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_8
timestamp 1636943256
transform 1 0 1840 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_20
timestamp 1636943256
transform 1 0 2944 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_32
timestamp 1636943256
transform 1 0 4048 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_44
timestamp -25199
transform 1 0 5152 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_52
timestamp -25199
transform 1 0 5888 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636943256
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp -25199
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_73
timestamp -25199
transform 1 0 7820 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_89
timestamp 1636943256
transform 1 0 9292 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp -25199
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1636943256
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1636943256
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1636943256
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_149
timestamp -25199
transform 1 0 14812 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp -25199
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1636943256
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_181
timestamp -25199
transform 1 0 17756 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636943256
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1636943256
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp -25199
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_36
timestamp -25199
transform 1 0 4416 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_44
timestamp -25199
transform 1 0 5152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_53
timestamp -25199
transform 1 0 5980 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_59
timestamp 1636943256
transform 1 0 6532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_71
timestamp -25199
transform 1 0 7636 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp -25199
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1636943256
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1636943256
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1636943256
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_121
timestamp -25199
transform 1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_125
timestamp -25199
transform 1 0 12604 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_150
timestamp -25199
transform 1 0 14904 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_160
timestamp -25199
transform 1 0 15824 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_169
timestamp -25199
transform 1 0 16652 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_187
timestamp -25199
transform 1 0 18308 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_8
timestamp 1636943256
transform 1 0 1840 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_20
timestamp 1636943256
transform 1 0 2944 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_32
timestamp -25199
transform 1 0 4048 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_36
timestamp -25199
transform 1 0 4416 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp -25199
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_57
timestamp -25199
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_72
timestamp -25199
transform 1 0 7728 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_76
timestamp -25199
transform 1 0 8096 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_85
timestamp -25199
transform 1 0 8924 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_91
timestamp -25199
transform 1 0 9476 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_97
timestamp -25199
transform 1 0 10028 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_140
timestamp -25199
transform 1 0 13984 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_154
timestamp -25199
transform 1 0 15272 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_178
timestamp 1636943256
transform 1 0 17480 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636943256
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636943256
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp -25199
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp -25199
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_38
timestamp 1636943256
transform 1 0 4600 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_50
timestamp -25199
transform 1 0 5704 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_56
timestamp -25199
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_64
timestamp 1636943256
transform 1 0 6992 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_76
timestamp -25199
transform 1 0 8096 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_80
timestamp -25199
transform 1 0 8464 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_102
timestamp -25199
transform 1 0 10488 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_113
timestamp -25199
transform 1 0 11500 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_119
timestamp -25199
transform 1 0 12052 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp -25199
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_141
timestamp -25199
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_147
timestamp 1636943256
transform 1 0 14628 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_159
timestamp -25199
transform 1 0 15732 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_165
timestamp -25199
transform 1 0 16284 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_169
timestamp 1636943256
transform 1 0 16652 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_181
timestamp -25199
transform 1 0 17756 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_189
timestamp -25199
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_8
timestamp 1636943256
transform 1 0 1840 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_20
timestamp 1636943256
transform 1 0 2944 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_32
timestamp -25199
transform 1 0 4048 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_39
timestamp -25199
transform 1 0 4692 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp -25199
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp -25199
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1636943256
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_69
timestamp -25199
transform 1 0 7452 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_73
timestamp -25199
transform 1 0 7820 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_88
timestamp 1636943256
transform 1 0 9200 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_100
timestamp 1636943256
transform 1 0 10304 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp -25199
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_121
timestamp -25199
transform 1 0 12236 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_126
timestamp -25199
transform 1 0 12696 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1636943256
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_149
timestamp -25199
transform 1 0 14812 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_153
timestamp -25199
transform 1 0 15180 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp -25199
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp -25199
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1636943256
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_181
timestamp -25199
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_189
timestamp -25199
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636943256
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636943256
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp -25199
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_29
timestamp -25199
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_37
timestamp -25199
transform 1 0 4508 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp -25199
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_57
timestamp -25199
transform 1 0 6348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1636943256
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_85
timestamp -25199
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_89
timestamp -25199
transform 1 0 9292 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_98
timestamp -25199
transform 1 0 10120 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_102
timestamp -25199
transform 1 0 10488 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_111
timestamp -25199
transform 1 0 11316 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_123
timestamp -25199
transform 1 0 12420 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_129
timestamp -25199
transform 1 0 12972 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp -25199
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_148
timestamp -25199
transform 1 0 14720 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_164
timestamp -25199
transform 1 0 16192 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_175
timestamp 1636943256
transform 1 0 17204 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_187
timestamp -25199
transform 1 0 18308 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_10
timestamp 1636943256
transform 1 0 2024 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_22
timestamp -25199
transform 1 0 3128 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_30
timestamp -25199
transform 1 0 3864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_47
timestamp -25199
transform 1 0 5428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp -25199
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp -25199
transform 1 0 6348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_68
timestamp -25199
transform 1 0 7360 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_76
timestamp -25199
transform 1 0 8096 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_92
timestamp -25199
transform 1 0 9568 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_96
timestamp -25199
transform 1 0 9936 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp -25199
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp -25199
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_131
timestamp -25199
transform 1 0 13156 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_134
timestamp -25199
transform 1 0 13432 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_142
timestamp -25199
transform 1 0 14168 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_150
timestamp -25199
transform 1 0 14904 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_155
timestamp -25199
transform 1 0 15364 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp -25199
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp -25199
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp -25199
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_175
timestamp -25199
transform 1 0 17204 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_180
timestamp -25199
transform 1 0 17664 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_187
timestamp -25199
transform 1 0 18308 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_14
timestamp 1636943256
transform 1 0 2392 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp -25199
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_29
timestamp -25199
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_34
timestamp -25199
transform 1 0 4232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_40
timestamp -25199
transform 1 0 4784 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_44
timestamp -25199
transform 1 0 5152 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_73
timestamp -25199
transform 1 0 7820 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_85
timestamp -25199
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_99
timestamp -25199
transform 1 0 10212 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_105
timestamp -25199
transform 1 0 10764 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp -25199
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_19
timestamp -25199
transform 1 0 2852 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_25
timestamp -25199
transform 1 0 3404 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_33
timestamp -25199
transform 1 0 4140 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_43
timestamp -25199
transform 1 0 5060 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_49
timestamp -25199
transform 1 0 5612 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp -25199
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_73
timestamp -25199
transform 1 0 7820 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_91
timestamp -25199
transform 1 0 9476 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_97
timestamp -25199
transform 1 0 10028 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_104
timestamp -25199
transform 1 0 10672 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp -25199
transform 1 0 12420 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_141
timestamp -25199
transform 1 0 14076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp -25199
transform 1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp -25199
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp -25199
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp -25199
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp -25199
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp -25199
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp -25199
transform 1 0 1380 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp -25199
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp -25199
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp -25199
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp -25199
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp -25199
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp -25199
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp -25199
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp -25199
transform 1 0 1748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp -25199
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp -25199
transform -1 0 1748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp -25199
transform 1 0 2024 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input19
timestamp -25199
transform 1 0 2576 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp -25199
transform 1 0 3128 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp -25199
transform 1 0 3772 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp -25199
transform 1 0 4232 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input23
timestamp -25199
transform 1 0 4784 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp -25199
transform 1 0 5336 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp -25199
transform -1 0 6256 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp -25199
transform -1 0 6808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input27
timestamp -25199
transform 1 0 7084 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp -25199
transform 1 0 7544 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp -25199
transform 1 0 8096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input30
timestamp -25199
transform 1 0 8924 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp -25199
transform 1 0 9200 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp -25199
transform 1 0 9752 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp -25199
transform 1 0 10304 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp -25199
transform 1 0 11500 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp -25199
transform -1 0 11408 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp -25199
transform 1 0 13432 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp -25199
transform 1 0 12512 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input38
timestamp -25199
transform 1 0 13708 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp -25199
transform -1 0 14352 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp -25199
transform 1 0 14168 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp -25199
transform -1 0 15456 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp -25199
transform -1 0 16376 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input43
timestamp -25199
transform -1 0 17664 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp -25199
transform 1 0 17204 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp -25199
transform -1 0 17388 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp -25199
transform 1 0 17480 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp -25199
transform -1 0 18308 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp -25199
transform -1 0 18584 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  output49
timestamp -25199
transform 1 0 18032 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output50
timestamp -25199
transform 1 0 18032 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output51
timestamp -25199
transform 1 0 18032 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output52
timestamp -25199
transform 1 0 18032 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output53
timestamp -25199
transform -1 0 2024 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output54
timestamp -25199
transform -1 0 2116 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output55
timestamp -25199
transform -1 0 3496 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output56
timestamp -25199
transform -1 0 3680 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output57
timestamp -25199
transform -1 0 4232 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output58
timestamp -25199
transform -1 0 4600 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output59
timestamp -25199
transform -1 0 5152 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output60
timestamp -25199
transform -1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output61
timestamp -25199
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output62
timestamp -25199
transform 1 0 6440 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output63
timestamp -25199
transform 1 0 6624 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output64
timestamp -25199
transform -1 0 7728 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output65
timestamp -25199
transform -1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output66
timestamp -25199
transform -1 0 8832 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output67
timestamp -25199
transform -1 0 9752 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output68
timestamp -25199
transform -1 0 10304 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output69
timestamp -25199
transform 1 0 10304 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output70
timestamp -25199
transform -1 0 11408 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output71
timestamp -25199
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output72
timestamp -25199
transform -1 0 12604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output73
timestamp -25199
transform 1 0 12604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output74
timestamp -25199
transform -1 0 13708 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output75
timestamp -25199
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output76
timestamp -25199
transform 1 0 14628 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output77
timestamp -25199
transform 1 0 15180 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output78
timestamp -25199
transform -1 0 16284 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output79
timestamp -25199
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output80
timestamp -25199
transform 1 0 17204 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output81
timestamp -25199
transform 1 0 17756 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output82
timestamp -25199
transform 1 0 17480 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output83
timestamp -25199
transform -1 0 18584 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output84
timestamp -25199
transform 1 0 17480 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_28
timestamp -25199
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -25199
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_29
timestamp -25199
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -25199
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_30
timestamp -25199
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -25199
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_31
timestamp -25199
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -25199
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_32
timestamp -25199
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -25199
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_33
timestamp -25199
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -25199
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_34
timestamp -25199
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -25199
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_35
timestamp -25199
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -25199
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_36
timestamp -25199
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -25199
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_37
timestamp -25199
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -25199
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_38
timestamp -25199
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -25199
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_39
timestamp -25199
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -25199
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_40
timestamp -25199
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -25199
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_41
timestamp -25199
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -25199
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_42
timestamp -25199
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -25199
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_43
timestamp -25199
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -25199
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_44
timestamp -25199
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -25199
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_45
timestamp -25199
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -25199
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_46
timestamp -25199
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -25199
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_47
timestamp -25199
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -25199
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_48
timestamp -25199
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -25199
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_49
timestamp -25199
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -25199
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_50
timestamp -25199
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -25199
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_51
timestamp -25199
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -25199
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_52
timestamp -25199
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -25199
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_53
timestamp -25199
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp -25199
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_54
timestamp -25199
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp -25199
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_55
timestamp -25199
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp -25199
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_56
timestamp -25199
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_57
timestamp -25199
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp -25199
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp -25199
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp -25199
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_61
timestamp -25199
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_62
timestamp -25199
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_63
timestamp -25199
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_64
timestamp -25199
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_65
timestamp -25199
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_66
timestamp -25199
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_67
timestamp -25199
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_68
timestamp -25199
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_69
timestamp -25199
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_70
timestamp -25199
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_71
timestamp -25199
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_72
timestamp -25199
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_73
timestamp -25199
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_74
timestamp -25199
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_75
timestamp -25199
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp -25199
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp -25199
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp -25199
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp -25199
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp -25199
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp -25199
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp -25199
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_83
timestamp -25199
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_84
timestamp -25199
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_85
timestamp -25199
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_86
timestamp -25199
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_87
timestamp -25199
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp -25199
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_89
timestamp -25199
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_90
timestamp -25199
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp -25199
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_92
timestamp -25199
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_93
timestamp -25199
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_94
timestamp -25199
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_95
timestamp -25199
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_96
timestamp -25199
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_97
timestamp -25199
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_98
timestamp -25199
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_99
timestamp -25199
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_100
timestamp -25199
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_101
timestamp -25199
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_102
timestamp -25199
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_103
timestamp -25199
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_104
timestamp -25199
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_105
timestamp -25199
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_106
timestamp -25199
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_107
timestamp -25199
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_108
timestamp -25199
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_109
timestamp -25199
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_110
timestamp -25199
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_111
timestamp -25199
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_112
timestamp -25199
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_113
timestamp -25199
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_114
timestamp -25199
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_115
timestamp -25199
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_116
timestamp -25199
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_117
timestamp -25199
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_118
timestamp -25199
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_119
timestamp -25199
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_120
timestamp -25199
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_121
timestamp -25199
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_122
timestamp -25199
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_123
timestamp -25199
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_124
timestamp -25199
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_125
timestamp -25199
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_126
timestamp -25199
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_127
timestamp -25199
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_128
timestamp -25199
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_129
timestamp -25199
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_130
timestamp -25199
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_131
timestamp -25199
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_132
timestamp -25199
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_133
timestamp -25199
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_134
timestamp -25199
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_135
timestamp -25199
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_136
timestamp -25199
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_137
timestamp -25199
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_138
timestamp -25199
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_139
timestamp -25199
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_140
timestamp -25199
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_141
timestamp -25199
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_142
timestamp -25199
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_143
timestamp -25199
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_144
timestamp -25199
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_145
timestamp -25199
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 bm_s0_s0_i[0]
port 0 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 bm_s0_s0_i[1]
port 1 nsew signal input
flabel metal3 s 0 3816 800 3936 0 FreeSans 480 0 0 0 bm_s0_s2_i[0]
port 2 nsew signal input
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 bm_s0_s2_i[1]
port 3 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 bm_s1_s0_i[0]
port 4 nsew signal input
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 bm_s1_s0_i[1]
port 5 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 bm_s1_s2_i[0]
port 6 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 bm_s1_s2_i[1]
port 7 nsew signal input
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 bm_s2_s1_i[0]
port 8 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 bm_s2_s1_i[1]
port 9 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 bm_s2_s3_i[0]
port 10 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 bm_s2_s3_i[1]
port 11 nsew signal input
flabel metal3 s 0 14696 800 14816 0 FreeSans 480 0 0 0 bm_s3_s1_i[0]
port 12 nsew signal input
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 bm_s3_s1_i[1]
port 13 nsew signal input
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 bm_s3_s3_i[0]
port 14 nsew signal input
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 bm_s3_s3_i[1]
port 15 nsew signal input
flabel metal3 s 19200 2456 20000 2576 0 FreeSans 480 0 0 0 dec_bits_o[0]
port 16 nsew signal output
flabel metal3 s 19200 7352 20000 7472 0 FreeSans 480 0 0 0 dec_bits_o[1]
port 17 nsew signal output
flabel metal3 s 19200 12248 20000 12368 0 FreeSans 480 0 0 0 dec_bits_o[2]
port 18 nsew signal output
flabel metal3 s 19200 17144 20000 17264 0 FreeSans 480 0 0 0 dec_bits_o[3]
port 19 nsew signal output
flabel metal2 s 1398 19200 1454 20000 0 FreeSans 224 90 0 0 pm_s0_i[0]
port 20 nsew signal input
flabel metal2 s 1950 19200 2006 20000 0 FreeSans 224 90 0 0 pm_s0_i[1]
port 21 nsew signal input
flabel metal2 s 2502 19200 2558 20000 0 FreeSans 224 90 0 0 pm_s0_i[2]
port 22 nsew signal input
flabel metal2 s 3054 19200 3110 20000 0 FreeSans 224 90 0 0 pm_s0_i[3]
port 23 nsew signal input
flabel metal2 s 3606 19200 3662 20000 0 FreeSans 224 90 0 0 pm_s0_i[4]
port 24 nsew signal input
flabel metal2 s 4158 19200 4214 20000 0 FreeSans 224 90 0 0 pm_s0_i[5]
port 25 nsew signal input
flabel metal2 s 4710 19200 4766 20000 0 FreeSans 224 90 0 0 pm_s0_i[6]
port 26 nsew signal input
flabel metal2 s 5262 19200 5318 20000 0 FreeSans 224 90 0 0 pm_s0_i[7]
port 27 nsew signal input
flabel metal2 s 1398 0 1454 800 0 FreeSans 224 90 0 0 pm_s0_o[0]
port 28 nsew signal output
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 pm_s0_o[1]
port 29 nsew signal output
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 pm_s0_o[2]
port 30 nsew signal output
flabel metal2 s 3054 0 3110 800 0 FreeSans 224 90 0 0 pm_s0_o[3]
port 31 nsew signal output
flabel metal2 s 3606 0 3662 800 0 FreeSans 224 90 0 0 pm_s0_o[4]
port 32 nsew signal output
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 pm_s0_o[5]
port 33 nsew signal output
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 pm_s0_o[6]
port 34 nsew signal output
flabel metal2 s 5262 0 5318 800 0 FreeSans 224 90 0 0 pm_s0_o[7]
port 35 nsew signal output
flabel metal2 s 5814 19200 5870 20000 0 FreeSans 224 90 0 0 pm_s1_i[0]
port 36 nsew signal input
flabel metal2 s 6366 19200 6422 20000 0 FreeSans 224 90 0 0 pm_s1_i[1]
port 37 nsew signal input
flabel metal2 s 6918 19200 6974 20000 0 FreeSans 224 90 0 0 pm_s1_i[2]
port 38 nsew signal input
flabel metal2 s 7470 19200 7526 20000 0 FreeSans 224 90 0 0 pm_s1_i[3]
port 39 nsew signal input
flabel metal2 s 8022 19200 8078 20000 0 FreeSans 224 90 0 0 pm_s1_i[4]
port 40 nsew signal input
flabel metal2 s 8574 19200 8630 20000 0 FreeSans 224 90 0 0 pm_s1_i[5]
port 41 nsew signal input
flabel metal2 s 9126 19200 9182 20000 0 FreeSans 224 90 0 0 pm_s1_i[6]
port 42 nsew signal input
flabel metal2 s 9678 19200 9734 20000 0 FreeSans 224 90 0 0 pm_s1_i[7]
port 43 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 pm_s1_o[0]
port 44 nsew signal output
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 pm_s1_o[1]
port 45 nsew signal output
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 pm_s1_o[2]
port 46 nsew signal output
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 pm_s1_o[3]
port 47 nsew signal output
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 pm_s1_o[4]
port 48 nsew signal output
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 pm_s1_o[5]
port 49 nsew signal output
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 pm_s1_o[6]
port 50 nsew signal output
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 pm_s1_o[7]
port 51 nsew signal output
flabel metal2 s 10230 19200 10286 20000 0 FreeSans 224 90 0 0 pm_s2_i[0]
port 52 nsew signal input
flabel metal2 s 10782 19200 10838 20000 0 FreeSans 224 90 0 0 pm_s2_i[1]
port 53 nsew signal input
flabel metal2 s 11334 19200 11390 20000 0 FreeSans 224 90 0 0 pm_s2_i[2]
port 54 nsew signal input
flabel metal2 s 11886 19200 11942 20000 0 FreeSans 224 90 0 0 pm_s2_i[3]
port 55 nsew signal input
flabel metal2 s 12438 19200 12494 20000 0 FreeSans 224 90 0 0 pm_s2_i[4]
port 56 nsew signal input
flabel metal2 s 12990 19200 13046 20000 0 FreeSans 224 90 0 0 pm_s2_i[5]
port 57 nsew signal input
flabel metal2 s 13542 19200 13598 20000 0 FreeSans 224 90 0 0 pm_s2_i[6]
port 58 nsew signal input
flabel metal2 s 14094 19200 14150 20000 0 FreeSans 224 90 0 0 pm_s2_i[7]
port 59 nsew signal input
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 pm_s2_o[0]
port 60 nsew signal output
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 pm_s2_o[1]
port 61 nsew signal output
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 pm_s2_o[2]
port 62 nsew signal output
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 pm_s2_o[3]
port 63 nsew signal output
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 pm_s2_o[4]
port 64 nsew signal output
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 pm_s2_o[5]
port 65 nsew signal output
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 pm_s2_o[6]
port 66 nsew signal output
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 pm_s2_o[7]
port 67 nsew signal output
flabel metal2 s 14646 19200 14702 20000 0 FreeSans 224 90 0 0 pm_s3_i[0]
port 68 nsew signal input
flabel metal2 s 15198 19200 15254 20000 0 FreeSans 224 90 0 0 pm_s3_i[1]
port 69 nsew signal input
flabel metal2 s 15750 19200 15806 20000 0 FreeSans 224 90 0 0 pm_s3_i[2]
port 70 nsew signal input
flabel metal2 s 16302 19200 16358 20000 0 FreeSans 224 90 0 0 pm_s3_i[3]
port 71 nsew signal input
flabel metal2 s 16854 19200 16910 20000 0 FreeSans 224 90 0 0 pm_s3_i[4]
port 72 nsew signal input
flabel metal2 s 17406 19200 17462 20000 0 FreeSans 224 90 0 0 pm_s3_i[5]
port 73 nsew signal input
flabel metal2 s 17958 19200 18014 20000 0 FreeSans 224 90 0 0 pm_s3_i[6]
port 74 nsew signal input
flabel metal2 s 18510 19200 18566 20000 0 FreeSans 224 90 0 0 pm_s3_i[7]
port 75 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 pm_s3_o[0]
port 76 nsew signal output
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 pm_s3_o[1]
port 77 nsew signal output
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 pm_s3_o[2]
port 78 nsew signal output
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 pm_s3_o[3]
port 79 nsew signal output
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 pm_s3_o[4]
port 80 nsew signal output
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 pm_s3_o[5]
port 81 nsew signal output
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 pm_s3_o[6]
port 82 nsew signal output
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 pm_s3_o[7]
port 83 nsew signal output
flabel metal4 s 4208 2128 4528 17456 0 FreeSans 1920 90 0 0 vccd1
port 84 nsew power bidirectional
flabel metal4 s 4868 2128 5188 17456 0 FreeSans 1920 90 0 0 vssd1
port 85 nsew ground bidirectional
rlabel metal1 9982 16864 9982 16864 0 vccd1
rlabel metal1 9982 17408 9982 17408 0 vssd1
rlabel metal1 13110 14042 13110 14042 0 _000_
rlabel metal2 15318 11900 15318 11900 0 _001_
rlabel metal2 15410 11934 15410 11934 0 _002_
rlabel metal1 16652 11798 16652 11798 0 _003_
rlabel metal1 14766 11764 14766 11764 0 _004_
rlabel metal2 14030 12036 14030 12036 0 _005_
rlabel metal2 15318 10234 15318 10234 0 _006_
rlabel metal1 13938 11118 13938 11118 0 _007_
rlabel metal1 12834 10608 12834 10608 0 _008_
rlabel metal1 13524 9962 13524 9962 0 _009_
rlabel metal1 13662 10166 13662 10166 0 _010_
rlabel metal2 13018 10438 13018 10438 0 _011_
rlabel metal1 12834 10438 12834 10438 0 _012_
rlabel metal2 13202 10438 13202 10438 0 _013_
rlabel metal1 13432 10778 13432 10778 0 _014_
rlabel metal2 14674 11458 14674 11458 0 _015_
rlabel metal1 14398 11594 14398 11594 0 _016_
rlabel metal1 15594 16762 15594 16762 0 _017_
rlabel metal1 16330 15538 16330 15538 0 _018_
rlabel metal1 15594 13906 15594 13906 0 _019_
rlabel metal1 16836 13498 16836 13498 0 _020_
rlabel metal1 14766 13328 14766 13328 0 _021_
rlabel metal1 16146 13940 16146 13940 0 _022_
rlabel metal2 16974 14144 16974 14144 0 _023_
rlabel metal1 14858 11866 14858 11866 0 _024_
rlabel metal2 14858 11492 14858 11492 0 _025_
rlabel metal1 17112 11730 17112 11730 0 _026_
rlabel metal1 18170 13362 18170 13362 0 _027_
rlabel metal1 17756 12206 17756 12206 0 _028_
rlabel metal1 17802 12138 17802 12138 0 _029_
rlabel metal1 17434 12240 17434 12240 0 _030_
rlabel metal1 17848 11730 17848 11730 0 _031_
rlabel metal1 16751 16558 16751 16558 0 _032_
rlabel metal1 17158 16592 17158 16592 0 _033_
rlabel metal2 18032 14484 18032 14484 0 _034_
rlabel metal2 14398 14076 14398 14076 0 _035_
rlabel metal2 14214 13906 14214 13906 0 _036_
rlabel metal1 16054 14450 16054 14450 0 _037_
rlabel metal1 17894 10098 17894 10098 0 _038_
rlabel metal2 18262 11900 18262 11900 0 _039_
rlabel metal2 16974 11118 16974 11118 0 _040_
rlabel metal1 16836 16490 16836 16490 0 _041_
rlabel metal1 17802 9588 17802 9588 0 _042_
rlabel metal1 15916 13770 15916 13770 0 _043_
rlabel metal2 16882 9860 16882 9860 0 _044_
rlabel metal1 16882 13804 16882 13804 0 _045_
rlabel metal1 16284 10030 16284 10030 0 _046_
rlabel metal1 8418 3468 8418 3468 0 _047_
rlabel metal1 8556 3026 8556 3026 0 _048_
rlabel metal1 9476 3026 9476 3026 0 _049_
rlabel metal2 9246 3332 9246 3332 0 _050_
rlabel metal2 2530 4386 2530 4386 0 _051_
rlabel metal1 8510 4692 8510 4692 0 _052_
rlabel metal2 9154 4964 9154 4964 0 _053_
rlabel metal1 11362 3570 11362 3570 0 _054_
rlabel metal1 1932 9554 1932 9554 0 _055_
rlabel metal1 2806 9588 2806 9588 0 _056_
rlabel metal2 2346 9350 2346 9350 0 _057_
rlabel metal1 8234 9384 8234 9384 0 _058_
rlabel metal2 11178 4284 11178 4284 0 _059_
rlabel metal1 10028 3502 10028 3502 0 _060_
rlabel metal2 9062 5814 9062 5814 0 _061_
rlabel metal1 10028 3570 10028 3570 0 _062_
rlabel metal1 9706 3434 9706 3434 0 _063_
rlabel metal1 10350 3502 10350 3502 0 _064_
rlabel metal2 12650 3842 12650 3842 0 _065_
rlabel metal1 12926 5644 12926 5644 0 _066_
rlabel metal2 13110 5100 13110 5100 0 _067_
rlabel metal1 12466 5201 12466 5201 0 _068_
rlabel metal1 13340 3162 13340 3162 0 _069_
rlabel metal2 12926 5168 12926 5168 0 _070_
rlabel metal1 13018 5168 13018 5168 0 _071_
rlabel metal1 13294 3094 13294 3094 0 _072_
rlabel metal1 12696 5270 12696 5270 0 _073_
rlabel metal1 12696 3978 12696 3978 0 _074_
rlabel metal2 12650 5508 12650 5508 0 _075_
rlabel metal2 9522 7990 9522 7990 0 _076_
rlabel metal1 11270 6732 11270 6732 0 _077_
rlabel metal1 11086 6800 11086 6800 0 _078_
rlabel metal1 12604 3162 12604 3162 0 _079_
rlabel metal2 11914 9248 11914 9248 0 _080_
rlabel metal2 11362 7004 11362 7004 0 _081_
rlabel metal1 12696 3094 12696 3094 0 _082_
rlabel metal2 12098 5882 12098 5882 0 _083_
rlabel metal1 13340 5882 13340 5882 0 _084_
rlabel metal1 13064 6834 13064 6834 0 _085_
rlabel metal1 13018 7344 13018 7344 0 _086_
rlabel metal1 13018 6766 13018 6766 0 _087_
rlabel metal1 12558 6732 12558 6732 0 _088_
rlabel metal2 13386 6460 13386 6460 0 _089_
rlabel metal1 13064 6290 13064 6290 0 _090_
rlabel metal1 9798 9044 9798 9044 0 _091_
rlabel metal1 10258 8432 10258 8432 0 _092_
rlabel metal2 14122 7956 14122 7956 0 _093_
rlabel metal1 13110 8976 13110 8976 0 _094_
rlabel metal1 12190 9010 12190 9010 0 _095_
rlabel metal2 14214 8126 14214 8126 0 _096_
rlabel metal2 14582 4828 14582 4828 0 _097_
rlabel metal1 14076 6426 14076 6426 0 _098_
rlabel metal1 13984 7446 13984 7446 0 _099_
rlabel metal2 13846 8262 13846 8262 0 _100_
rlabel metal2 14306 6970 14306 6970 0 _101_
rlabel metal2 5658 15674 5658 15674 0 _102_
rlabel metal2 5014 15776 5014 15776 0 _103_
rlabel metal1 5198 14926 5198 14926 0 _104_
rlabel via1 6486 14926 6486 14926 0 _105_
rlabel metal2 7314 11356 7314 11356 0 _106_
rlabel metal2 6946 14110 6946 14110 0 _107_
rlabel metal2 4278 12002 4278 12002 0 _108_
rlabel metal1 4094 12206 4094 12206 0 _109_
rlabel metal2 4462 12070 4462 12070 0 _110_
rlabel metal2 12558 14076 12558 14076 0 _111_
rlabel metal1 7268 13906 7268 13906 0 _112_
rlabel metal1 6302 13192 6302 13192 0 _113_
rlabel metal2 5474 14076 5474 14076 0 _114_
rlabel metal2 6118 12444 6118 12444 0 _115_
rlabel metal1 6670 13498 6670 13498 0 _116_
rlabel metal2 4554 14212 4554 14212 0 _117_
rlabel metal1 4968 13770 4968 13770 0 _118_
rlabel metal2 5750 13668 5750 13668 0 _119_
rlabel metal2 5934 13702 5934 13702 0 _120_
rlabel metal1 8602 14008 8602 14008 0 _121_
rlabel viali 9064 12821 9064 12821 0 _122_
rlabel metal1 9246 12852 9246 12852 0 _123_
rlabel metal1 8740 11866 8740 11866 0 _124_
rlabel metal1 9016 12342 9016 12342 0 _125_
rlabel metal1 9062 13430 9062 13430 0 _126_
rlabel metal1 9062 11798 9062 11798 0 _127_
rlabel metal1 8142 12954 8142 12954 0 _128_
rlabel metal1 8050 13906 8050 13906 0 _129_
rlabel metal1 9200 14994 9200 14994 0 _130_
rlabel metal1 9292 15130 9292 15130 0 _131_
rlabel metal1 9062 14314 9062 14314 0 _132_
rlabel metal2 13110 15028 13110 15028 0 _133_
rlabel metal1 11270 14450 11270 14450 0 _134_
rlabel metal2 10442 14212 10442 14212 0 _135_
rlabel metal1 9522 14382 9522 14382 0 _136_
rlabel metal1 8786 13940 8786 13940 0 _137_
rlabel metal1 8740 12954 8740 12954 0 _138_
rlabel metal1 8234 13804 8234 13804 0 _139_
rlabel metal1 10350 16014 10350 16014 0 _140_
rlabel metal1 9016 16218 9016 16218 0 _141_
rlabel metal1 10028 16082 10028 16082 0 _142_
rlabel metal1 10996 15470 10996 15470 0 _143_
rlabel metal1 13662 16694 13662 16694 0 _144_
rlabel metal1 13018 16490 13018 16490 0 _145_
rlabel metal2 12558 16014 12558 16014 0 _146_
rlabel metal1 11132 16082 11132 16082 0 _147_
rlabel metal1 14122 15606 14122 15606 0 _148_
rlabel metal2 13478 15300 13478 15300 0 _149_
rlabel metal2 12834 15504 12834 15504 0 _150_
rlabel metal1 10534 15470 10534 15470 0 _151_
rlabel metal2 11270 15810 11270 15810 0 _152_
rlabel metal1 12558 16116 12558 16116 0 _153_
rlabel metal2 12650 15810 12650 15810 0 _154_
rlabel metal1 12236 16150 12236 16150 0 _155_
rlabel metal1 4278 2618 4278 2618 0 _156_
rlabel metal1 4370 3026 4370 3026 0 _157_
rlabel metal1 3128 2278 3128 2278 0 _158_
rlabel metal1 3404 3502 3404 3502 0 _159_
rlabel metal1 4462 3570 4462 3570 0 _160_
rlabel metal2 4922 7446 4922 7446 0 _161_
rlabel metal1 5750 5066 5750 5066 0 _162_
rlabel metal1 3174 7412 3174 7412 0 _163_
rlabel metal2 2714 5984 2714 5984 0 _164_
rlabel metal1 2415 6222 2415 6222 0 _165_
rlabel metal1 6900 7854 6900 7854 0 _166_
rlabel metal2 5382 3536 5382 3536 0 _167_
rlabel metal1 5796 5202 5796 5202 0 _168_
rlabel metal2 2622 4624 2622 4624 0 _169_
rlabel metal2 3726 5712 3726 5712 0 _170_
rlabel metal1 2645 3094 2645 3094 0 _171_
rlabel metal2 2530 6154 2530 6154 0 _172_
rlabel metal2 2346 4012 2346 4012 0 _173_
rlabel metal1 3312 5270 3312 5270 0 _174_
rlabel metal1 4140 5202 4140 5202 0 _175_
rlabel metal1 5290 5338 5290 5338 0 _176_
rlabel metal1 6762 5712 6762 5712 0 _177_
rlabel metal1 5750 5644 5750 5644 0 _178_
rlabel metal2 5382 4896 5382 4896 0 _179_
rlabel metal2 6578 5610 6578 5610 0 _180_
rlabel metal1 6394 5168 6394 5168 0 _181_
rlabel metal2 5474 4692 5474 4692 0 _182_
rlabel metal1 6532 5882 6532 5882 0 _183_
rlabel metal1 6440 5338 6440 5338 0 _184_
rlabel metal1 6946 5882 6946 5882 0 _185_
rlabel via1 4654 9894 4654 9894 0 _186_
rlabel metal2 6670 7004 6670 7004 0 _187_
rlabel metal1 5382 7344 5382 7344 0 _188_
rlabel metal1 4876 6766 4876 6766 0 _189_
rlabel metal2 8050 9724 8050 9724 0 _190_
rlabel metal1 6578 7820 6578 7820 0 _191_
rlabel metal1 5152 6698 5152 6698 0 _192_
rlabel metal1 6992 6290 6992 6290 0 _193_
rlabel metal1 6440 6426 6440 6426 0 _194_
rlabel metal1 7130 8534 7130 8534 0 _195_
rlabel metal1 5428 8534 5428 8534 0 _196_
rlabel metal1 4830 8466 4830 8466 0 _197_
rlabel metal2 6946 8262 6946 8262 0 _198_
rlabel metal1 6578 8602 6578 8602 0 _199_
rlabel metal1 5888 8942 5888 8942 0 _200_
rlabel metal1 5428 10030 5428 10030 0 _201_
rlabel metal1 5244 10030 5244 10030 0 _202_
rlabel metal1 5980 9962 5980 9962 0 _203_
rlabel metal1 8694 10132 8694 10132 0 _204_
rlabel metal2 8326 9690 8326 9690 0 _205_
rlabel metal1 6532 10030 6532 10030 0 _206_
rlabel metal1 5336 9622 5336 9622 0 _207_
rlabel metal2 6670 9282 6670 9282 0 _208_
rlabel metal1 7406 10132 7406 10132 0 _209_
rlabel metal2 6854 10234 6854 10234 0 _210_
rlabel metal1 6440 9554 6440 9554 0 _211_
rlabel metal1 11270 12172 11270 12172 0 _212_
rlabel metal1 9062 6426 9062 6426 0 _213_
rlabel metal1 9200 6086 9200 6086 0 _214_
rlabel metal2 10810 4352 10810 4352 0 _215_
rlabel metal1 8832 6698 8832 6698 0 _216_
rlabel metal1 6624 16218 6624 16218 0 _217_
rlabel metal1 6900 16626 6900 16626 0 _218_
rlabel metal1 6900 16558 6900 16558 0 _219_
rlabel metal1 15364 16558 15364 16558 0 _220_
rlabel metal1 15502 11764 15502 11764 0 _221_
rlabel metal1 15548 12614 15548 12614 0 _222_
rlabel metal1 16606 11866 16606 11866 0 _223_
rlabel metal1 10166 11662 10166 11662 0 _224_
rlabel metal1 11730 10676 11730 10676 0 _225_
rlabel metal1 11822 10642 11822 10642 0 _226_
rlabel metal1 2714 2380 2714 2380 0 bm_s0_s0_i[0]
rlabel metal1 1380 2414 1380 2414 0 bm_s0_s0_i[1]
rlabel metal1 1380 3502 1380 3502 0 bm_s0_s2_i[0]
rlabel metal1 1380 5202 1380 5202 0 bm_s0_s2_i[1]
rlabel metal1 1380 5882 1380 5882 0 bm_s1_s0_i[0]
rlabel metal1 1380 7378 1380 7378 0 bm_s1_s0_i[1]
rlabel metal1 1288 7922 1288 7922 0 bm_s1_s2_i[0]
rlabel metal1 1380 10030 1380 10030 0 bm_s1_s2_i[1]
rlabel metal1 1380 10642 1380 10642 0 bm_s2_s1_i[0]
rlabel metal1 1380 11730 1380 11730 0 bm_s2_s1_i[1]
rlabel metal1 1380 12818 1380 12818 0 bm_s2_s3_i[0]
rlabel metal1 1380 13906 1380 13906 0 bm_s2_s3_i[1]
rlabel metal1 1380 14994 1380 14994 0 bm_s3_s1_i[0]
rlabel metal1 1380 16082 1380 16082 0 bm_s3_s1_i[1]
rlabel metal1 1794 17136 1794 17136 0 bm_s3_s3_i[0]
rlabel metal3 1050 18020 1050 18020 0 bm_s3_s3_i[1]
rlabel metal3 18868 2516 18868 2516 0 dec_bits_o[0]
rlabel metal2 18354 7599 18354 7599 0 dec_bits_o[1]
rlabel metal3 18868 12308 18868 12308 0 dec_bits_o[2]
rlabel metal2 18354 16881 18354 16881 0 dec_bits_o[3]
rlabel metal1 3358 2618 3358 2618 0 net1
rlabel metal1 3358 11628 3358 11628 0 net10
rlabel metal2 14306 13634 14306 13634 0 net100
rlabel metal1 13294 13906 13294 13906 0 net101
rlabel metal2 12374 14518 12374 14518 0 net102
rlabel metal2 13662 13260 13662 13260 0 net103
rlabel metal1 12650 13940 12650 13940 0 net104
rlabel metal2 12466 8874 12466 8874 0 net105
rlabel metal1 7452 5202 7452 5202 0 net106
rlabel metal2 7866 5440 7866 5440 0 net107
rlabel metal2 10534 8126 10534 8126 0 net108
rlabel metal1 3726 8874 3726 8874 0 net109
rlabel metal1 6578 12648 6578 12648 0 net11
rlabel metal1 4462 8976 4462 8976 0 net110
rlabel metal1 3956 2414 3956 2414 0 net111
rlabel metal2 1610 12376 1610 12376 0 net12
rlabel metal1 2185 15130 2185 15130 0 net13
rlabel metal1 4186 15980 4186 15980 0 net14
rlabel metal1 1978 17068 1978 17068 0 net15
rlabel metal1 1610 16456 1610 16456 0 net16
rlabel metal1 1886 16694 1886 16694 0 net17
rlabel metal1 2116 4046 2116 4046 0 net18
rlabel metal2 4784 15708 4784 15708 0 net19
rlabel metal1 1794 3570 1794 3570 0 net2
rlabel metal1 3450 16966 3450 16966 0 net20
rlabel metal1 3956 16966 3956 16966 0 net21
rlabel metal1 4600 17034 4600 17034 0 net22
rlabel metal1 5198 16966 5198 16966 0 net23
rlabel metal2 5980 14756 5980 14756 0 net24
rlabel metal1 2162 5712 2162 5712 0 net25
rlabel metal1 1886 8534 1886 8534 0 net26
rlabel metal1 7452 16966 7452 16966 0 net27
rlabel metal1 7866 16966 7866 16966 0 net28
rlabel metal1 9246 17034 9246 17034 0 net29
rlabel metal1 6486 3502 6486 3502 0 net3
rlabel metal1 9108 16966 9108 16966 0 net30
rlabel metal1 9522 16966 9522 16966 0 net31
rlabel metal2 13570 9418 13570 9418 0 net32
rlabel metal1 4416 13294 4416 13294 0 net33
rlabel metal1 9890 11662 9890 11662 0 net34
rlabel metal1 11408 14382 11408 14382 0 net35
rlabel metal1 12788 14994 12788 14994 0 net36
rlabel metal2 12650 14569 12650 14569 0 net37
rlabel metal1 14214 16082 14214 16082 0 net38
rlabel metal2 13386 15555 13386 15555 0 net39
rlabel metal2 2162 4794 2162 4794 0 net4
rlabel metal2 14490 16286 14490 16286 0 net40
rlabel metal1 15088 17034 15088 17034 0 net41
rlabel metal1 6348 16558 6348 16558 0 net42
rlabel metal2 14766 16371 14766 16371 0 net43
rlabel metal1 15318 16048 15318 16048 0 net44
rlabel metal1 15778 15028 15778 15028 0 net45
rlabel metal1 16836 17170 16836 17170 0 net46
rlabel metal1 15778 16150 15778 16150 0 net47
rlabel metal1 15870 16626 15870 16626 0 net48
rlabel metal1 6164 9486 6164 9486 0 net49
rlabel metal2 1610 6562 1610 6562 0 net5
rlabel metal2 11730 16388 11730 16388 0 net50
rlabel metal1 14030 6834 14030 6834 0 net51
rlabel metal1 17986 16558 17986 16558 0 net52
rlabel metal1 1932 2618 1932 2618 0 net53
rlabel metal1 2116 3026 2116 3026 0 net54
rlabel metal1 3450 2958 3450 2958 0 net55
rlabel metal1 3634 2448 3634 2448 0 net56
rlabel metal1 4186 3060 4186 3060 0 net57
rlabel metal1 4738 2448 4738 2448 0 net58
rlabel metal1 5290 2448 5290 2448 0 net59
rlabel metal2 1610 7956 1610 7956 0 net6
rlabel metal1 5658 2482 5658 2482 0 net60
rlabel metal2 5842 13061 5842 13061 0 net61
rlabel metal1 6578 3026 6578 3026 0 net62
rlabel metal1 5842 2448 5842 2448 0 net63
rlabel metal1 7912 11526 7912 11526 0 net64
rlabel metal3 8671 2516 8671 2516 0 net65
rlabel metal3 8855 2652 8855 2652 0 net66
rlabel metal1 9752 2414 9752 2414 0 net67
rlabel metal1 10856 2482 10856 2482 0 net68
rlabel metal1 10396 2822 10396 2822 0 net69
rlabel metal1 2116 7854 2116 7854 0 net7
rlabel metal1 11316 2822 11316 2822 0 net70
rlabel metal2 11546 2618 11546 2618 0 net71
rlabel metal1 12880 2890 12880 2890 0 net72
rlabel metal2 12650 2618 12650 2618 0 net73
rlabel metal1 13616 6630 13616 6630 0 net74
rlabel metal2 14122 3434 14122 3434 0 net75
rlabel metal1 14720 6630 14720 6630 0 net76
rlabel metal1 15410 2414 15410 2414 0 net77
rlabel metal1 16146 9894 16146 9894 0 net78
rlabel metal1 16192 10166 16192 10166 0 net79
rlabel metal2 1610 9724 1610 9724 0 net8
rlabel metal1 17342 11526 17342 11526 0 net80
rlabel metal1 17572 14042 17572 14042 0 net81
rlabel metal1 17572 3026 17572 3026 0 net82
rlabel metal2 18538 6460 18538 6460 0 net83
rlabel metal2 17526 6426 17526 6426 0 net84
rlabel metal1 2668 2958 2668 2958 0 net85
rlabel metal2 18078 3706 18078 3706 0 net86
rlabel metal1 9384 14450 9384 14450 0 net87
rlabel metal2 11086 15708 11086 15708 0 net88
rlabel metal1 14858 4658 14858 4658 0 net89
rlabel metal2 4094 12891 4094 12891 0 net9
rlabel metal1 18124 12818 18124 12818 0 net90
rlabel metal1 15042 10064 15042 10064 0 net91
rlabel metal1 9890 16626 9890 16626 0 net92
rlabel metal2 12374 9078 12374 9078 0 net93
rlabel metal2 16238 13668 16238 13668 0 net94
rlabel via2 13110 16405 13110 16405 0 net95
rlabel viali 15216 12818 15216 12818 0 net96
rlabel metal2 15134 16354 15134 16354 0 net97
rlabel metal1 6670 14382 6670 14382 0 net98
rlabel metal1 14720 12886 14720 12886 0 net99
rlabel metal2 1472 18156 1472 18156 0 pm_s0_i[0]
rlabel metal1 2070 17238 2070 17238 0 pm_s0_i[1]
rlabel metal2 2530 18268 2530 18268 0 pm_s0_i[2]
rlabel metal2 3082 18268 3082 18268 0 pm_s0_i[3]
rlabel metal2 3634 18268 3634 18268 0 pm_s0_i[4]
rlabel metal1 4278 17238 4278 17238 0 pm_s0_i[5]
rlabel metal1 4784 17170 4784 17170 0 pm_s0_i[6]
rlabel metal1 5336 17170 5336 17170 0 pm_s0_i[7]
rlabel metal2 1426 2404 1426 2404 0 pm_s0_o[0]
rlabel metal2 1978 1163 1978 1163 0 pm_s0_o[1]
rlabel metal2 2530 1826 2530 1826 0 pm_s0_o[2]
rlabel metal2 3082 1554 3082 1554 0 pm_s0_o[3]
rlabel metal1 3772 2958 3772 2958 0 pm_s0_o[4]
rlabel metal2 4186 1554 4186 1554 0 pm_s0_o[5]
rlabel metal2 4738 1554 4738 1554 0 pm_s0_o[6]
rlabel metal2 5290 1554 5290 1554 0 pm_s0_o[7]
rlabel metal1 6026 17170 6026 17170 0 pm_s1_i[0]
rlabel metal1 6532 17238 6532 17238 0 pm_s1_i[1]
rlabel metal1 7130 17204 7130 17204 0 pm_s1_i[2]
rlabel metal2 7498 18268 7498 18268 0 pm_s1_i[3]
rlabel metal2 8050 18268 8050 18268 0 pm_s1_i[4]
rlabel metal2 8602 18268 8602 18268 0 pm_s1_i[5]
rlabel metal1 9200 17170 9200 17170 0 pm_s1_i[6]
rlabel metal2 9706 18268 9706 18268 0 pm_s1_i[7]
rlabel metal2 5842 1554 5842 1554 0 pm_s1_o[0]
rlabel metal1 6532 2958 6532 2958 0 pm_s1_o[1]
rlabel metal2 6946 1554 6946 1554 0 pm_s1_o[2]
rlabel metal2 7498 1554 7498 1554 0 pm_s1_o[3]
rlabel metal2 8050 1554 8050 1554 0 pm_s1_o[4]
rlabel metal2 8602 1554 8602 1554 0 pm_s1_o[5]
rlabel metal2 9154 1554 9154 1554 0 pm_s1_o[6]
rlabel metal2 9706 1520 9706 1520 0 pm_s1_o[7]
rlabel metal2 10258 18268 10258 18268 0 pm_s2_i[0]
rlabel metal1 10948 17306 10948 17306 0 pm_s2_i[1]
rlabel metal1 11270 17170 11270 17170 0 pm_s2_i[2]
rlabel via1 13294 17170 13294 17170 0 pm_s2_i[3]
rlabel metal1 12512 17170 12512 17170 0 pm_s2_i[4]
rlabel metal2 14030 16762 14030 16762 0 pm_s2_i[5]
rlabel metal1 13984 16490 13984 16490 0 pm_s2_i[6]
rlabel metal1 14168 17170 14168 17170 0 pm_s2_i[7]
rlabel metal2 10258 1520 10258 1520 0 pm_s2_o[0]
rlabel metal2 10810 1554 10810 1554 0 pm_s2_o[1]
rlabel metal2 11362 1520 11362 1520 0 pm_s2_o[2]
rlabel metal2 11914 1554 11914 1554 0 pm_s2_o[3]
rlabel metal2 12466 1554 12466 1554 0 pm_s2_o[4]
rlabel metal2 13018 1554 13018 1554 0 pm_s2_o[5]
rlabel metal2 13570 1554 13570 1554 0 pm_s2_o[6]
rlabel metal2 14122 1520 14122 1520 0 pm_s2_o[7]
rlabel metal1 14996 17170 14996 17170 0 pm_s3_i[0]
rlabel metal1 15824 17306 15824 17306 0 pm_s3_i[1]
rlabel metal1 17296 17170 17296 17170 0 pm_s3_i[2]
rlabel metal1 16698 16150 16698 16150 0 pm_s3_i[3]
rlabel metal1 17250 17272 17250 17272 0 pm_s3_i[4]
rlabel metal1 17618 16558 17618 16558 0 pm_s3_i[5]
rlabel metal2 17986 17724 17986 17724 0 pm_s3_i[6]
rlabel metal2 18538 18200 18538 18200 0 pm_s3_i[7]
rlabel metal2 14674 959 14674 959 0 pm_s3_o[0]
rlabel metal2 15226 1520 15226 1520 0 pm_s3_o[1]
rlabel metal1 16882 2414 16882 2414 0 pm_s3_o[2]
rlabel metal2 16330 1554 16330 1554 0 pm_s3_o[3]
rlabel metal2 16882 1520 16882 1520 0 pm_s3_o[4]
rlabel metal1 17572 2958 17572 2958 0 pm_s3_o[5]
rlabel metal1 18124 2958 18124 2958 0 pm_s3_o[6]
rlabel metal2 18538 1231 18538 1231 0 pm_s3_o[7]
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
