magic
tech sky130A
magscale 1 2
timestamp 1769196221
<< viali >>
rect 2145 11849 2179 11883
rect 1593 11781 1627 11815
rect 3433 11781 3467 11815
rect 10701 11781 10735 11815
rect 1869 11713 1903 11747
rect 2053 11713 2087 11747
rect 2513 11713 2547 11747
rect 2697 11713 2731 11747
rect 2973 11713 3007 11747
rect 3249 11713 3283 11747
rect 10977 11713 11011 11747
rect 2881 11577 2915 11611
rect 2421 11509 2455 11543
rect 3157 11509 3191 11543
rect 10977 11305 11011 11339
rect 6469 11237 6503 11271
rect 3157 11169 3191 11203
rect 4629 11169 4663 11203
rect 3249 11101 3283 11135
rect 3433 11101 3467 11135
rect 6653 11101 6687 11135
rect 8309 11101 8343 11135
rect 9229 11101 9263 11135
rect 2881 11033 2915 11067
rect 3341 11033 3375 11067
rect 4905 11033 4939 11067
rect 7849 11033 7883 11067
rect 8033 11033 8067 11067
rect 9505 11033 9539 11067
rect 1409 10965 1443 10999
rect 6377 10965 6411 10999
rect 8401 10965 8435 10999
rect 2605 10761 2639 10795
rect 5181 10761 5215 10795
rect 5549 10761 5583 10795
rect 9597 10761 9631 10795
rect 3617 10693 3651 10727
rect 1409 10625 1443 10659
rect 1685 10625 1719 10659
rect 1869 10625 1903 10659
rect 2053 10625 2087 10659
rect 2145 10625 2179 10659
rect 3341 10625 3375 10659
rect 9137 10625 9171 10659
rect 9229 10625 9263 10659
rect 9413 10625 9447 10659
rect 2697 10557 2731 10591
rect 5641 10557 5675 10591
rect 5733 10557 5767 10591
rect 6377 10557 6411 10591
rect 6653 10557 6687 10591
rect 8217 10557 8251 10591
rect 8493 10557 8527 10591
rect 2421 10489 2455 10523
rect 2973 10489 3007 10523
rect 1593 10421 1627 10455
rect 2053 10421 2087 10455
rect 3157 10421 3191 10455
rect 5089 10421 5123 10455
rect 8125 10421 8159 10455
rect 2513 10217 2547 10251
rect 3801 10217 3835 10251
rect 5273 10217 5307 10251
rect 7297 10217 7331 10251
rect 1869 10149 1903 10183
rect 1961 10081 1995 10115
rect 4445 10081 4479 10115
rect 7849 10081 7883 10115
rect 1409 10013 1443 10047
rect 1685 10013 1719 10047
rect 4169 10013 4203 10047
rect 4629 10013 4663 10047
rect 4905 10013 4939 10047
rect 5089 10013 5123 10047
rect 7665 10013 7699 10047
rect 8125 10013 8159 10047
rect 8401 10013 8435 10047
rect 8493 10013 8527 10047
rect 8585 10013 8619 10047
rect 2145 9945 2179 9979
rect 2697 9945 2731 9979
rect 2881 9945 2915 9979
rect 4767 9945 4801 9979
rect 4997 9945 5031 9979
rect 5457 9945 5491 9979
rect 8263 9945 8297 9979
rect 1593 9877 1627 9911
rect 4261 9877 4295 9911
rect 6745 9877 6779 9911
rect 7757 9877 7791 9911
rect 8769 9877 8803 9911
rect 7021 9673 7055 9707
rect 1685 9605 1719 9639
rect 3341 9605 3375 9639
rect 3617 9605 3651 9639
rect 5707 9605 5741 9639
rect 5825 9605 5859 9639
rect 5916 9605 5950 9639
rect 6515 9605 6549 9639
rect 1409 9537 1443 9571
rect 3111 9537 3145 9571
rect 3249 9537 3283 9571
rect 3433 9537 3467 9571
rect 3893 9537 3927 9571
rect 4077 9537 4111 9571
rect 4905 9537 4939 9571
rect 4997 9537 5031 9571
rect 5365 9537 5399 9571
rect 6008 9537 6042 9571
rect 6653 9537 6687 9571
rect 6745 9537 6779 9571
rect 6837 9537 6871 9571
rect 2973 9469 3007 9503
rect 5549 9469 5583 9503
rect 6377 9469 6411 9503
rect 1593 9401 1627 9435
rect 4261 9401 4295 9435
rect 3801 9333 3835 9367
rect 5273 9333 5307 9367
rect 6193 9333 6227 9367
rect 7021 9061 7055 9095
rect 1685 8993 1719 9027
rect 8953 8993 8987 9027
rect 1409 8925 1443 8959
rect 8769 8925 8803 8959
rect 9229 8925 9263 8959
rect 1961 8857 1995 8891
rect 8493 8857 8527 8891
rect 1593 8789 1627 8823
rect 3433 8789 3467 8823
rect 1593 8585 1627 8619
rect 2421 8585 2455 8619
rect 2789 8585 2823 8619
rect 8125 8585 8159 8619
rect 8309 8585 8343 8619
rect 8953 8585 8987 8619
rect 1685 8517 1719 8551
rect 5457 8517 5491 8551
rect 1409 8449 1443 8483
rect 1869 8449 1903 8483
rect 5227 8449 5261 8483
rect 5365 8449 5399 8483
rect 5549 8449 5583 8483
rect 6377 8449 6411 8483
rect 8217 8449 8251 8483
rect 8493 8449 8527 8483
rect 8769 8449 8803 8483
rect 2881 8381 2915 8415
rect 2973 8381 3007 8415
rect 5089 8381 5123 8415
rect 6653 8381 6687 8415
rect 8677 8313 8711 8347
rect 5733 8245 5767 8279
rect 2513 8041 2547 8075
rect 6837 8041 6871 8075
rect 4077 7905 4111 7939
rect 6285 7905 6319 7939
rect 6377 7905 6411 7939
rect 1409 7837 1443 7871
rect 1777 7837 1811 7871
rect 2697 7837 2731 7871
rect 2789 7837 2823 7871
rect 3157 7837 3191 7871
rect 6469 7837 6503 7871
rect 2881 7769 2915 7803
rect 2999 7769 3033 7803
rect 4353 7769 4387 7803
rect 1593 7701 1627 7735
rect 5825 7701 5859 7735
rect 4721 7497 4755 7531
rect 5089 7497 5123 7531
rect 6035 7429 6069 7463
rect 9505 7429 9539 7463
rect 1409 7361 1443 7395
rect 3433 7361 3467 7395
rect 3525 7361 3559 7395
rect 3617 7361 3651 7395
rect 3735 7361 3769 7395
rect 5181 7361 5215 7395
rect 5549 7361 5583 7395
rect 5733 7361 5767 7395
rect 5825 7361 5859 7395
rect 5917 7361 5951 7395
rect 6193 7361 6227 7395
rect 9229 7361 9263 7395
rect 1685 7293 1719 7327
rect 3893 7293 3927 7327
rect 5273 7293 5307 7327
rect 3249 7225 3283 7259
rect 3157 7157 3191 7191
rect 10977 7157 11011 7191
rect 2237 6953 2271 6987
rect 3249 6953 3283 6987
rect 1593 6885 1627 6919
rect 2789 6817 2823 6851
rect 6653 6817 6687 6851
rect 10793 6817 10827 6851
rect 1409 6749 1443 6783
rect 1685 6749 1719 6783
rect 3157 6749 3191 6783
rect 10977 6749 11011 6783
rect 1961 6681 1995 6715
rect 2605 6681 2639 6715
rect 4813 6681 4847 6715
rect 6929 6681 6963 6715
rect 1869 6613 1903 6647
rect 2697 6613 2731 6647
rect 4629 6613 4663 6647
rect 6101 6613 6135 6647
rect 8401 6613 8435 6647
rect 1593 6409 1627 6443
rect 7389 6409 7423 6443
rect 1685 6341 1719 6375
rect 8769 6341 8803 6375
rect 9321 6341 9355 6375
rect 1409 6273 1443 6307
rect 1869 6273 1903 6307
rect 6377 6273 6411 6307
rect 6653 6273 6687 6307
rect 7573 6273 7607 6307
rect 7849 6273 7883 6307
rect 8033 6273 8067 6307
rect 8217 6273 8251 6307
rect 8493 6273 8527 6307
rect 8953 6273 8987 6307
rect 2145 6205 2179 6239
rect 2421 6205 2455 6239
rect 4445 6205 4479 6239
rect 4721 6205 4755 6239
rect 7665 6205 7699 6239
rect 8125 6205 8159 6239
rect 8585 6205 8619 6239
rect 7757 6137 7791 6171
rect 3893 6069 3927 6103
rect 6193 6069 6227 6103
rect 8309 6069 8343 6103
rect 8769 6069 8803 6103
rect 9321 6069 9355 6103
rect 9505 6069 9539 6103
rect 2605 5865 2639 5899
rect 4997 5865 5031 5899
rect 1593 5797 1627 5831
rect 7941 5797 7975 5831
rect 3249 5729 3283 5763
rect 5549 5729 5583 5763
rect 6469 5729 6503 5763
rect 8033 5729 8067 5763
rect 8953 5729 8987 5763
rect 1409 5661 1443 5695
rect 1685 5661 1719 5695
rect 2973 5661 3007 5695
rect 5365 5661 5399 5695
rect 6009 5661 6043 5695
rect 7573 5661 7607 5695
rect 8125 5661 8159 5695
rect 8217 5661 8251 5695
rect 8401 5661 8435 5695
rect 8585 5661 8619 5695
rect 6101 5593 6135 5627
rect 6193 5593 6227 5627
rect 6311 5593 6345 5627
rect 8493 5593 8527 5627
rect 9229 5593 9263 5627
rect 3065 5525 3099 5559
rect 5457 5525 5491 5559
rect 5825 5525 5859 5559
rect 8769 5525 8803 5559
rect 10701 5525 10735 5559
rect 3249 5321 3283 5355
rect 7757 5321 7791 5355
rect 8401 5321 8435 5355
rect 8585 5321 8619 5355
rect 10977 5321 11011 5355
rect 2763 5253 2797 5287
rect 2973 5253 3007 5287
rect 6745 5253 6779 5287
rect 6863 5253 6897 5287
rect 9505 5253 9539 5287
rect 1409 5185 1443 5219
rect 1685 5185 1719 5219
rect 2881 5185 2915 5219
rect 3065 5185 3099 5219
rect 6561 5185 6595 5219
rect 6653 5185 6687 5219
rect 7481 5185 7515 5219
rect 7941 5185 7975 5219
rect 8953 5185 8987 5219
rect 2605 5117 2639 5151
rect 4445 5117 4479 5151
rect 4721 5117 4755 5151
rect 7021 5117 7055 5151
rect 8125 5117 8159 5151
rect 9229 5117 9263 5151
rect 7665 5049 7699 5083
rect 1593 4981 1627 5015
rect 6193 4981 6227 5015
rect 6377 4981 6411 5015
rect 8585 4981 8619 5015
rect 3157 4777 3191 4811
rect 8125 4777 8159 4811
rect 4169 4709 4203 4743
rect 8309 4709 8343 4743
rect 7389 4641 7423 4675
rect 7573 4641 7607 4675
rect 8677 4641 8711 4675
rect 1409 4573 1443 4607
rect 4629 4573 4663 4607
rect 5089 4573 5123 4607
rect 6745 4573 6779 4607
rect 7481 4573 7515 4607
rect 7665 4573 7699 4607
rect 8493 4573 8527 4607
rect 8585 4573 8619 4607
rect 1685 4505 1719 4539
rect 4353 4505 4387 4539
rect 8033 4505 8067 4539
rect 7205 4437 7239 4471
rect 2145 4233 2179 4267
rect 2513 4233 2547 4267
rect 5089 4233 5123 4267
rect 5549 4233 5583 4267
rect 8493 4233 8527 4267
rect 3459 4165 3493 4199
rect 4445 4165 4479 4199
rect 5457 4165 5491 4199
rect 7021 4165 7055 4199
rect 1409 4097 1443 4131
rect 1685 4097 1719 4131
rect 2605 4097 2639 4131
rect 2973 4097 3007 4131
rect 3157 4097 3191 4131
rect 3249 4097 3283 4131
rect 3341 4097 3375 4131
rect 4215 4097 4249 4131
rect 4353 4097 4387 4131
rect 4537 4097 4571 4131
rect 6745 4097 6779 4131
rect 1961 4029 1995 4063
rect 2697 4029 2731 4063
rect 3617 4029 3651 4063
rect 4077 4029 4111 4063
rect 5641 4029 5675 4063
rect 1593 3961 1627 3995
rect 1869 3893 1903 3927
rect 4721 3893 4755 3927
rect 1685 3689 1719 3723
rect 3893 3689 3927 3723
rect 1593 3621 1627 3655
rect 4169 3621 4203 3655
rect 5273 3553 5307 3587
rect 5365 3553 5399 3587
rect 1409 3485 1443 3519
rect 2053 3485 2087 3519
rect 2421 3485 2455 3519
rect 2513 3485 2547 3519
rect 2697 3485 2731 3519
rect 2881 3485 2915 3519
rect 5181 3485 5215 3519
rect 2145 3417 2179 3451
rect 2237 3417 2271 3451
rect 2789 3417 2823 3451
rect 3249 3417 3283 3451
rect 3985 3417 4019 3451
rect 4353 3417 4387 3451
rect 1869 3349 1903 3383
rect 3065 3349 3099 3383
rect 3341 3349 3375 3383
rect 4813 3349 4847 3383
rect 1593 3145 1627 3179
rect 4353 3145 4387 3179
rect 6193 3145 6227 3179
rect 1685 3077 1719 3111
rect 2881 3077 2915 3111
rect 4721 3077 4755 3111
rect 9505 3077 9539 3111
rect 1409 3009 1443 3043
rect 1869 3009 1903 3043
rect 9229 3009 9263 3043
rect 2605 2941 2639 2975
rect 4445 2941 4479 2975
rect 10977 2805 11011 2839
rect 3157 2601 3191 2635
rect 1409 2465 1443 2499
rect 10977 2397 11011 2431
rect 1685 2329 1719 2363
rect 10701 2329 10735 2363
<< metal1 >>
rect 1104 11994 11316 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 11316 11994
rect 1104 11920 11316 11942
rect 2133 11883 2191 11889
rect 2133 11849 2145 11883
rect 2179 11880 2191 11883
rect 4798 11880 4804 11892
rect 2179 11852 4804 11880
rect 2179 11849 2191 11852
rect 2133 11843 2191 11849
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 1302 11772 1308 11824
rect 1360 11812 1366 11824
rect 1581 11815 1639 11821
rect 1581 11812 1593 11815
rect 1360 11784 1593 11812
rect 1360 11772 1366 11784
rect 1581 11781 1593 11784
rect 1627 11781 1639 11815
rect 3421 11815 3479 11821
rect 3421 11812 3433 11815
rect 1581 11775 1639 11781
rect 1780 11784 3433 11812
rect 1118 11704 1124 11756
rect 1176 11744 1182 11756
rect 1780 11744 1808 11784
rect 1176 11716 1808 11744
rect 1176 11704 1182 11716
rect 1854 11704 1860 11756
rect 1912 11704 1918 11756
rect 2041 11747 2099 11753
rect 2041 11713 2053 11747
rect 2087 11744 2099 11747
rect 2406 11744 2412 11756
rect 2087 11716 2412 11744
rect 2087 11713 2099 11716
rect 2041 11707 2099 11713
rect 2406 11704 2412 11716
rect 2464 11704 2470 11756
rect 2498 11704 2504 11756
rect 2556 11704 2562 11756
rect 2700 11753 2728 11784
rect 3421 11781 3433 11784
rect 3467 11781 3479 11815
rect 3421 11775 3479 11781
rect 10686 11772 10692 11824
rect 10744 11772 10750 11824
rect 2685 11747 2743 11753
rect 2685 11713 2697 11747
rect 2731 11713 2743 11747
rect 2685 11707 2743 11713
rect 2961 11747 3019 11753
rect 2961 11713 2973 11747
rect 3007 11744 3019 11747
rect 3237 11747 3295 11753
rect 3237 11744 3249 11747
rect 3007 11716 3249 11744
rect 3007 11713 3019 11716
rect 2961 11707 3019 11713
rect 3237 11713 3249 11716
rect 3283 11713 3295 11747
rect 3237 11707 3295 11713
rect 1210 11636 1216 11688
rect 1268 11676 1274 11688
rect 2976 11676 3004 11707
rect 10962 11704 10968 11756
rect 11020 11704 11026 11756
rect 1268 11648 3004 11676
rect 1268 11636 1274 11648
rect 2869 11611 2927 11617
rect 2869 11577 2881 11611
rect 2915 11608 2927 11611
rect 5718 11608 5724 11620
rect 2915 11580 5724 11608
rect 2915 11577 2927 11580
rect 2869 11571 2927 11577
rect 5718 11568 5724 11580
rect 5776 11568 5782 11620
rect 2406 11500 2412 11552
rect 2464 11540 2470 11552
rect 3050 11540 3056 11552
rect 2464 11512 3056 11540
rect 2464 11500 2470 11512
rect 3050 11500 3056 11512
rect 3108 11500 3114 11552
rect 3142 11500 3148 11552
rect 3200 11500 3206 11552
rect 1104 11450 11316 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 11316 11450
rect 1104 11376 11316 11398
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 2832 11308 6040 11336
rect 2832 11296 2838 11308
rect 3145 11203 3203 11209
rect 3145 11169 3157 11203
rect 3191 11200 3203 11203
rect 3326 11200 3332 11212
rect 3191 11172 3332 11200
rect 3191 11169 3203 11172
rect 3145 11163 3203 11169
rect 3326 11160 3332 11172
rect 3384 11200 3390 11212
rect 4617 11203 4675 11209
rect 4617 11200 4629 11203
rect 3384 11172 4629 11200
rect 3384 11160 3390 11172
rect 4617 11169 4629 11172
rect 4663 11200 4675 11203
rect 5442 11200 5448 11212
rect 4663 11172 5448 11200
rect 4663 11169 4675 11172
rect 4617 11163 4675 11169
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 6012 11200 6040 11308
rect 10962 11296 10968 11348
rect 11020 11296 11026 11348
rect 6454 11228 6460 11280
rect 6512 11228 6518 11280
rect 7466 11200 7472 11212
rect 6012 11172 7472 11200
rect 3234 11092 3240 11144
rect 3292 11092 3298 11144
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11101 3479 11135
rect 6012 11118 6040 11172
rect 7466 11160 7472 11172
rect 7524 11160 7530 11212
rect 3421 11095 3479 11101
rect 2774 11064 2780 11076
rect 2438 11036 2780 11064
rect 2774 11024 2780 11036
rect 2832 11024 2838 11076
rect 2869 11067 2927 11073
rect 2869 11033 2881 11067
rect 2915 11064 2927 11067
rect 3329 11067 3387 11073
rect 3329 11064 3341 11067
rect 2915 11036 3341 11064
rect 2915 11033 2927 11036
rect 2869 11027 2927 11033
rect 3329 11033 3341 11036
rect 3375 11033 3387 11067
rect 3436 11064 3464 11095
rect 6638 11092 6644 11144
rect 6696 11132 6702 11144
rect 8297 11135 8355 11141
rect 8297 11132 8309 11135
rect 6696 11104 8309 11132
rect 6696 11092 6702 11104
rect 8297 11101 8309 11104
rect 8343 11101 8355 11135
rect 8297 11095 8355 11101
rect 8754 11092 8760 11144
rect 8812 11132 8818 11144
rect 9217 11135 9275 11141
rect 9217 11132 9229 11135
rect 8812 11104 9229 11132
rect 8812 11092 8818 11104
rect 9217 11101 9229 11104
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 4798 11064 4804 11076
rect 3436 11036 4804 11064
rect 3329 11027 3387 11033
rect 4798 11024 4804 11036
rect 4856 11024 4862 11076
rect 4893 11067 4951 11073
rect 4893 11033 4905 11067
rect 4939 11033 4951 11067
rect 4893 11027 4951 11033
rect 1397 10999 1455 11005
rect 1397 10965 1409 10999
rect 1443 10996 1455 10999
rect 1854 10996 1860 11008
rect 1443 10968 1860 10996
rect 1443 10965 1455 10968
rect 1397 10959 1455 10965
rect 1854 10956 1860 10968
rect 1912 10956 1918 11008
rect 4908 10996 4936 11027
rect 7742 11024 7748 11076
rect 7800 11064 7806 11076
rect 7837 11067 7895 11073
rect 7837 11064 7849 11067
rect 7800 11036 7849 11064
rect 7800 11024 7806 11036
rect 7837 11033 7849 11036
rect 7883 11033 7895 11067
rect 7837 11027 7895 11033
rect 8021 11067 8079 11073
rect 8021 11033 8033 11067
rect 8067 11064 8079 11067
rect 8662 11064 8668 11076
rect 8067 11036 8668 11064
rect 8067 11033 8079 11036
rect 8021 11027 8079 11033
rect 8662 11024 8668 11036
rect 8720 11024 8726 11076
rect 9490 11024 9496 11076
rect 9548 11024 9554 11076
rect 9950 11024 9956 11076
rect 10008 11024 10014 11076
rect 5258 10996 5264 11008
rect 4908 10968 5264 10996
rect 5258 10956 5264 10968
rect 5316 10956 5322 11008
rect 6362 10956 6368 11008
rect 6420 10956 6426 11008
rect 8110 10956 8116 11008
rect 8168 10996 8174 11008
rect 8389 10999 8447 11005
rect 8389 10996 8401 10999
rect 8168 10968 8401 10996
rect 8168 10956 8174 10968
rect 8389 10965 8401 10968
rect 8435 10965 8447 10999
rect 8389 10959 8447 10965
rect 1104 10906 11316 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 11316 10906
rect 1104 10832 11316 10854
rect 2593 10795 2651 10801
rect 2593 10761 2605 10795
rect 2639 10792 2651 10795
rect 5169 10795 5227 10801
rect 2639 10764 5120 10792
rect 2639 10761 2651 10764
rect 2593 10755 2651 10761
rect 3602 10684 3608 10736
rect 3660 10684 3666 10736
rect 3878 10684 3884 10736
rect 3936 10724 3942 10736
rect 3936 10696 4094 10724
rect 3936 10684 3942 10696
rect 4890 10684 4896 10736
rect 4948 10684 4954 10736
rect 5092 10724 5120 10764
rect 5169 10761 5181 10795
rect 5215 10792 5227 10795
rect 5258 10792 5264 10804
rect 5215 10764 5264 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 5537 10795 5595 10801
rect 5537 10761 5549 10795
rect 5583 10792 5595 10795
rect 5810 10792 5816 10804
rect 5583 10764 5816 10792
rect 5583 10761 5595 10764
rect 5537 10755 5595 10761
rect 5810 10752 5816 10764
rect 5868 10792 5874 10804
rect 6362 10792 6368 10804
rect 5868 10764 6368 10792
rect 5868 10752 5874 10764
rect 6362 10752 6368 10764
rect 6420 10752 6426 10804
rect 9490 10752 9496 10804
rect 9548 10792 9554 10804
rect 9585 10795 9643 10801
rect 9585 10792 9597 10795
rect 9548 10764 9597 10792
rect 9548 10752 9554 10764
rect 9585 10761 9597 10764
rect 9631 10761 9643 10795
rect 9585 10755 9643 10761
rect 6638 10724 6644 10736
rect 5092 10696 6644 10724
rect 6638 10684 6644 10696
rect 6696 10684 6702 10736
rect 8018 10724 8024 10736
rect 7866 10696 8024 10724
rect 8018 10684 8024 10696
rect 8076 10684 8082 10736
rect 1302 10616 1308 10668
rect 1360 10656 1366 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 1360 10628 1409 10656
rect 1360 10616 1366 10628
rect 1397 10625 1409 10628
rect 1443 10656 1455 10659
rect 1673 10659 1731 10665
rect 1673 10656 1685 10659
rect 1443 10628 1685 10656
rect 1443 10625 1455 10628
rect 1397 10619 1455 10625
rect 1673 10625 1685 10628
rect 1719 10625 1731 10659
rect 1673 10619 1731 10625
rect 1854 10616 1860 10668
rect 1912 10616 1918 10668
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 2133 10659 2191 10665
rect 2133 10656 2145 10659
rect 2087 10628 2145 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 2133 10625 2145 10628
rect 2179 10656 2191 10659
rect 2179 10628 3004 10656
rect 2179 10625 2191 10628
rect 2133 10619 2191 10625
rect 1872 10520 1900 10616
rect 2682 10588 2688 10600
rect 2424 10560 2688 10588
rect 2424 10529 2452 10560
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 2976 10532 3004 10628
rect 3326 10616 3332 10668
rect 3384 10616 3390 10668
rect 4908 10656 4936 10684
rect 9125 10659 9183 10665
rect 9125 10656 9137 10659
rect 4908 10628 5764 10656
rect 3068 10560 5212 10588
rect 2409 10523 2467 10529
rect 2409 10520 2421 10523
rect 1872 10492 2421 10520
rect 2409 10489 2421 10492
rect 2455 10489 2467 10523
rect 2409 10483 2467 10489
rect 2958 10480 2964 10532
rect 3016 10480 3022 10532
rect 1581 10455 1639 10461
rect 1581 10421 1593 10455
rect 1627 10452 1639 10455
rect 1854 10452 1860 10464
rect 1627 10424 1860 10452
rect 1627 10421 1639 10424
rect 1581 10415 1639 10421
rect 1854 10412 1860 10424
rect 1912 10412 1918 10464
rect 2038 10412 2044 10464
rect 2096 10412 2102 10464
rect 2498 10412 2504 10464
rect 2556 10452 2562 10464
rect 3068 10452 3096 10560
rect 2556 10424 3096 10452
rect 3145 10455 3203 10461
rect 2556 10412 2562 10424
rect 3145 10421 3157 10455
rect 3191 10452 3203 10455
rect 4062 10452 4068 10464
rect 3191 10424 4068 10452
rect 3191 10421 3203 10424
rect 3145 10415 3203 10421
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 4890 10412 4896 10464
rect 4948 10452 4954 10464
rect 5077 10455 5135 10461
rect 5077 10452 5089 10455
rect 4948 10424 5089 10452
rect 4948 10412 4954 10424
rect 5077 10421 5089 10424
rect 5123 10421 5135 10455
rect 5184 10452 5212 10560
rect 5258 10548 5264 10600
rect 5316 10588 5322 10600
rect 5736 10597 5764 10628
rect 8588 10628 9137 10656
rect 8588 10600 8616 10628
rect 9125 10625 9137 10628
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 9214 10616 9220 10668
rect 9272 10616 9278 10668
rect 9306 10616 9312 10668
rect 9364 10656 9370 10668
rect 9401 10659 9459 10665
rect 9401 10656 9413 10659
rect 9364 10628 9413 10656
rect 9364 10616 9370 10628
rect 9401 10625 9413 10628
rect 9447 10625 9459 10659
rect 9401 10619 9459 10625
rect 5629 10591 5687 10597
rect 5629 10588 5641 10591
rect 5316 10560 5641 10588
rect 5316 10548 5322 10560
rect 5629 10557 5641 10560
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10557 5779 10591
rect 5721 10551 5779 10557
rect 6365 10591 6423 10597
rect 6365 10557 6377 10591
rect 6411 10557 6423 10591
rect 6365 10551 6423 10557
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10588 6699 10591
rect 7282 10588 7288 10600
rect 6687 10560 7288 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 5534 10480 5540 10532
rect 5592 10520 5598 10532
rect 6380 10520 6408 10551
rect 7282 10548 7288 10560
rect 7340 10548 7346 10600
rect 7926 10548 7932 10600
rect 7984 10588 7990 10600
rect 8205 10591 8263 10597
rect 8205 10588 8217 10591
rect 7984 10560 8217 10588
rect 7984 10548 7990 10560
rect 8205 10557 8217 10560
rect 8251 10557 8263 10591
rect 8205 10551 8263 10557
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10588 8539 10591
rect 8570 10588 8576 10600
rect 8527 10560 8576 10588
rect 8527 10557 8539 10560
rect 8481 10551 8539 10557
rect 8570 10548 8576 10560
rect 8628 10548 8634 10600
rect 5592 10492 6408 10520
rect 5592 10480 5598 10492
rect 6270 10452 6276 10464
rect 5184 10424 6276 10452
rect 5077 10415 5135 10421
rect 6270 10412 6276 10424
rect 6328 10412 6334 10464
rect 6380 10452 6408 10492
rect 6730 10452 6736 10464
rect 6380 10424 6736 10452
rect 6730 10412 6736 10424
rect 6788 10412 6794 10464
rect 8113 10455 8171 10461
rect 8113 10421 8125 10455
rect 8159 10452 8171 10455
rect 8386 10452 8392 10464
rect 8159 10424 8392 10452
rect 8159 10421 8171 10424
rect 8113 10415 8171 10421
rect 8386 10412 8392 10424
rect 8444 10412 8450 10464
rect 1104 10362 11316 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 11316 10362
rect 1104 10288 11316 10310
rect 2498 10208 2504 10260
rect 2556 10208 2562 10260
rect 3602 10208 3608 10260
rect 3660 10248 3666 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 3660 10220 3801 10248
rect 3660 10208 3666 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 3789 10211 3847 10217
rect 5258 10208 5264 10260
rect 5316 10208 5322 10260
rect 7282 10208 7288 10260
rect 7340 10208 7346 10260
rect 1857 10183 1915 10189
rect 1857 10149 1869 10183
rect 1903 10180 1915 10183
rect 1903 10152 5580 10180
rect 1903 10149 1915 10152
rect 1857 10143 1915 10149
rect 1118 10072 1124 10124
rect 1176 10112 1182 10124
rect 1949 10115 2007 10121
rect 1949 10112 1961 10115
rect 1176 10084 1961 10112
rect 1176 10072 1182 10084
rect 1210 10004 1216 10056
rect 1268 10044 1274 10056
rect 1688 10053 1716 10084
rect 1949 10081 1961 10084
rect 1995 10081 2007 10115
rect 1949 10075 2007 10081
rect 4430 10072 4436 10124
rect 4488 10072 4494 10124
rect 4540 10084 4936 10112
rect 1397 10047 1455 10053
rect 1397 10044 1409 10047
rect 1268 10016 1409 10044
rect 1268 10004 1274 10016
rect 1397 10013 1409 10016
rect 1443 10013 1455 10047
rect 1397 10007 1455 10013
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10013 1731 10047
rect 1673 10007 1731 10013
rect 1412 9976 1440 10007
rect 1854 10004 1860 10056
rect 1912 10044 1918 10056
rect 4157 10047 4215 10053
rect 1912 10016 3740 10044
rect 1912 10004 1918 10016
rect 2133 9979 2191 9985
rect 2133 9976 2145 9979
rect 1412 9948 2145 9976
rect 2133 9945 2145 9948
rect 2179 9945 2191 9979
rect 2133 9939 2191 9945
rect 2682 9936 2688 9988
rect 2740 9936 2746 9988
rect 2869 9979 2927 9985
rect 2869 9945 2881 9979
rect 2915 9976 2927 9979
rect 2958 9976 2964 9988
rect 2915 9948 2964 9976
rect 2915 9945 2927 9948
rect 2869 9939 2927 9945
rect 1578 9868 1584 9920
rect 1636 9868 1642 9920
rect 2884 9908 2912 9939
rect 2958 9936 2964 9948
rect 3016 9936 3022 9988
rect 3712 9976 3740 10016
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4540 10044 4568 10084
rect 4908 10056 4936 10084
rect 4203 10016 4568 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 4614 10004 4620 10056
rect 4672 10004 4678 10056
rect 4890 10004 4896 10056
rect 4948 10004 4954 10056
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10044 5135 10047
rect 5258 10044 5264 10056
rect 5123 10016 5264 10044
rect 5123 10013 5135 10016
rect 5077 10007 5135 10013
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 4755 9979 4813 9985
rect 4755 9976 4767 9979
rect 3712 9948 4767 9976
rect 4755 9945 4767 9948
rect 4801 9945 4813 9979
rect 4755 9939 4813 9945
rect 4985 9979 5043 9985
rect 4985 9945 4997 9979
rect 5031 9945 5043 9979
rect 4985 9939 5043 9945
rect 4154 9908 4160 9920
rect 2884 9880 4160 9908
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 4246 9868 4252 9920
rect 4304 9868 4310 9920
rect 4522 9868 4528 9920
rect 4580 9908 4586 9920
rect 5000 9908 5028 9939
rect 5442 9936 5448 9988
rect 5500 9936 5506 9988
rect 5552 9976 5580 10152
rect 6638 10140 6644 10192
rect 6696 10180 6702 10192
rect 7742 10180 7748 10192
rect 6696 10152 7748 10180
rect 6696 10140 6702 10152
rect 7742 10140 7748 10152
rect 7800 10180 7806 10192
rect 7800 10152 8524 10180
rect 7800 10140 7806 10152
rect 6270 10072 6276 10124
rect 6328 10112 6334 10124
rect 7837 10115 7895 10121
rect 7837 10112 7849 10115
rect 6328 10084 7849 10112
rect 6328 10072 6334 10084
rect 7837 10081 7849 10084
rect 7883 10081 7895 10115
rect 7837 10075 7895 10081
rect 8036 10084 8432 10112
rect 7653 10047 7711 10053
rect 7653 10013 7665 10047
rect 7699 10044 7711 10047
rect 8036 10044 8064 10084
rect 8404 10056 8432 10084
rect 7699 10016 8064 10044
rect 7699 10013 7711 10016
rect 7653 10007 7711 10013
rect 8110 10004 8116 10056
rect 8168 10004 8174 10056
rect 8386 10004 8392 10056
rect 8444 10004 8450 10056
rect 8496 10053 8524 10152
rect 8481 10047 8539 10053
rect 8481 10013 8493 10047
rect 8527 10013 8539 10047
rect 8481 10007 8539 10013
rect 8570 10004 8576 10056
rect 8628 10044 8634 10056
rect 9030 10044 9036 10056
rect 8628 10016 9036 10044
rect 8628 10004 8634 10016
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 8251 9979 8309 9985
rect 8251 9976 8263 9979
rect 5552 9948 8263 9976
rect 8251 9945 8263 9948
rect 8297 9945 8309 9979
rect 8251 9939 8309 9945
rect 5534 9908 5540 9920
rect 4580 9880 5540 9908
rect 4580 9868 4586 9880
rect 5534 9868 5540 9880
rect 5592 9908 5598 9920
rect 6638 9908 6644 9920
rect 5592 9880 6644 9908
rect 5592 9868 5598 9880
rect 6638 9868 6644 9880
rect 6696 9868 6702 9920
rect 6730 9868 6736 9920
rect 6788 9868 6794 9920
rect 7742 9868 7748 9920
rect 7800 9868 7806 9920
rect 7834 9868 7840 9920
rect 7892 9908 7898 9920
rect 8110 9908 8116 9920
rect 7892 9880 8116 9908
rect 7892 9868 7898 9880
rect 8110 9868 8116 9880
rect 8168 9868 8174 9920
rect 8757 9911 8815 9917
rect 8757 9877 8769 9911
rect 8803 9908 8815 9911
rect 9398 9908 9404 9920
rect 8803 9880 9404 9908
rect 8803 9877 8815 9880
rect 8757 9871 8815 9877
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 1104 9818 11316 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 11316 9818
rect 1104 9744 11316 9766
rect 1578 9664 1584 9716
rect 1636 9704 1642 9716
rect 1636 9676 6132 9704
rect 1636 9664 1642 9676
rect 6104 9674 6132 9676
rect 1673 9639 1731 9645
rect 1673 9636 1685 9639
rect 1412 9608 1685 9636
rect 1302 9528 1308 9580
rect 1360 9568 1366 9580
rect 1412 9577 1440 9608
rect 1673 9605 1685 9608
rect 1719 9605 1731 9639
rect 1673 9599 1731 9605
rect 2774 9596 2780 9648
rect 2832 9636 2838 9648
rect 3329 9639 3387 9645
rect 3329 9636 3341 9639
rect 2832 9608 3341 9636
rect 2832 9596 2838 9608
rect 3329 9605 3341 9608
rect 3375 9636 3387 9639
rect 3510 9636 3516 9648
rect 3375 9608 3516 9636
rect 3375 9605 3387 9608
rect 3329 9599 3387 9605
rect 3510 9596 3516 9608
rect 3568 9596 3574 9648
rect 3605 9639 3663 9645
rect 3605 9605 3617 9639
rect 3651 9636 3663 9639
rect 4246 9636 4252 9648
rect 3651 9608 4252 9636
rect 3651 9605 3663 9608
rect 3605 9599 3663 9605
rect 4246 9596 4252 9608
rect 4304 9596 4310 9648
rect 5718 9645 5724 9648
rect 5695 9639 5724 9645
rect 5695 9605 5707 9639
rect 5695 9599 5724 9605
rect 5718 9596 5724 9599
rect 5776 9596 5782 9648
rect 5810 9596 5816 9648
rect 5868 9596 5874 9648
rect 5902 9596 5908 9648
rect 5960 9596 5966 9648
rect 6104 9646 6224 9674
rect 6638 9664 6644 9716
rect 6696 9664 6702 9716
rect 6730 9664 6736 9716
rect 6788 9704 6794 9716
rect 7009 9707 7067 9713
rect 6788 9676 6868 9704
rect 6788 9664 6794 9676
rect 6196 9636 6224 9646
rect 6503 9639 6561 9645
rect 6503 9636 6515 9639
rect 6196 9608 6515 9636
rect 6503 9605 6515 9608
rect 6549 9605 6561 9639
rect 6656 9636 6684 9664
rect 6840 9636 6868 9676
rect 7009 9673 7021 9707
rect 7055 9704 7067 9707
rect 7742 9704 7748 9716
rect 7055 9676 7748 9704
rect 7055 9673 7067 9676
rect 7009 9667 7067 9673
rect 7742 9664 7748 9676
rect 7800 9664 7806 9716
rect 8754 9636 8760 9648
rect 6656 9608 6776 9636
rect 6840 9608 8760 9636
rect 6503 9599 6561 9605
rect 1397 9571 1455 9577
rect 1397 9568 1409 9571
rect 1360 9540 1409 9568
rect 1360 9528 1366 9540
rect 1397 9537 1409 9540
rect 1443 9537 1455 9571
rect 3099 9571 3157 9577
rect 3099 9568 3111 9571
rect 1397 9531 1455 9537
rect 1596 9540 3111 9568
rect 1596 9441 1624 9540
rect 3099 9537 3111 9540
rect 3145 9537 3157 9571
rect 3099 9531 3157 9537
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9537 3295 9571
rect 3237 9531 3295 9537
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9568 3479 9571
rect 3786 9568 3792 9580
rect 3467 9540 3792 9568
rect 3467 9537 3479 9540
rect 3421 9531 3479 9537
rect 2961 9503 3019 9509
rect 2961 9469 2973 9503
rect 3007 9469 3019 9503
rect 3252 9500 3280 9531
rect 3786 9528 3792 9540
rect 3844 9528 3850 9580
rect 3881 9571 3939 9577
rect 3881 9537 3893 9571
rect 3927 9537 3939 9571
rect 3881 9531 3939 9537
rect 3896 9500 3924 9531
rect 4062 9528 4068 9580
rect 4120 9528 4126 9580
rect 4154 9528 4160 9580
rect 4212 9568 4218 9580
rect 4890 9568 4896 9580
rect 4212 9540 4896 9568
rect 4212 9528 4218 9540
rect 4890 9528 4896 9540
rect 4948 9528 4954 9580
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 5350 9568 5356 9580
rect 5031 9540 5356 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5350 9528 5356 9540
rect 5408 9528 5414 9580
rect 5996 9571 6054 9577
rect 5736 9566 5948 9568
rect 5996 9566 6008 9571
rect 5736 9540 6008 9566
rect 5736 9512 5764 9540
rect 5920 9538 6008 9540
rect 5996 9537 6008 9538
rect 6042 9537 6054 9571
rect 5996 9531 6054 9537
rect 6638 9528 6644 9580
rect 6696 9528 6702 9580
rect 6748 9577 6776 9608
rect 8754 9596 8760 9608
rect 8812 9596 8818 9648
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9537 6791 9571
rect 6733 9531 6791 9537
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9568 6883 9571
rect 6914 9568 6920 9580
rect 6871 9540 6920 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 6914 9528 6920 9540
rect 6972 9568 6978 9580
rect 7926 9568 7932 9580
rect 6972 9540 7932 9568
rect 6972 9528 6978 9540
rect 7926 9528 7932 9540
rect 7984 9528 7990 9580
rect 5258 9500 5264 9512
rect 3252 9472 3464 9500
rect 3896 9472 5264 9500
rect 2961 9463 3019 9469
rect 1581 9435 1639 9441
rect 1581 9401 1593 9435
rect 1627 9401 1639 9435
rect 2976 9432 3004 9463
rect 3436 9444 3464 9472
rect 3142 9432 3148 9444
rect 2976 9404 3148 9432
rect 1581 9395 1639 9401
rect 3142 9392 3148 9404
rect 3200 9392 3206 9444
rect 3418 9392 3424 9444
rect 3476 9392 3482 9444
rect 3510 9392 3516 9444
rect 3568 9432 3574 9444
rect 4264 9441 4292 9472
rect 5258 9460 5264 9472
rect 5316 9460 5322 9512
rect 5537 9503 5595 9509
rect 5537 9469 5549 9503
rect 5583 9500 5595 9503
rect 5626 9500 5632 9512
rect 5583 9472 5632 9500
rect 5583 9469 5595 9472
rect 5537 9463 5595 9469
rect 5626 9460 5632 9472
rect 5684 9460 5690 9512
rect 5718 9460 5724 9512
rect 5776 9460 5782 9512
rect 6178 9460 6184 9512
rect 6236 9500 6242 9512
rect 6365 9503 6423 9509
rect 6365 9500 6377 9503
rect 6236 9472 6377 9500
rect 6236 9460 6242 9472
rect 6365 9469 6377 9472
rect 6411 9469 6423 9503
rect 6365 9463 6423 9469
rect 6454 9460 6460 9512
rect 6512 9500 6518 9512
rect 9306 9500 9312 9512
rect 6512 9472 9312 9500
rect 6512 9460 6518 9472
rect 9306 9460 9312 9472
rect 9364 9460 9370 9512
rect 4249 9435 4307 9441
rect 3568 9404 4200 9432
rect 3568 9392 3574 9404
rect 3786 9324 3792 9376
rect 3844 9324 3850 9376
rect 4172 9364 4200 9404
rect 4249 9401 4261 9435
rect 4295 9401 4307 9435
rect 4249 9395 4307 9401
rect 5902 9392 5908 9444
rect 5960 9432 5966 9444
rect 8294 9432 8300 9444
rect 5960 9404 8300 9432
rect 5960 9392 5966 9404
rect 8294 9392 8300 9404
rect 8352 9432 8358 9444
rect 9214 9432 9220 9444
rect 8352 9404 9220 9432
rect 8352 9392 8358 9404
rect 9214 9392 9220 9404
rect 9272 9392 9278 9444
rect 4522 9364 4528 9376
rect 4172 9336 4528 9364
rect 4522 9324 4528 9336
rect 4580 9324 4586 9376
rect 4614 9324 4620 9376
rect 4672 9364 4678 9376
rect 5261 9367 5319 9373
rect 5261 9364 5273 9367
rect 4672 9336 5273 9364
rect 4672 9324 4678 9336
rect 5261 9333 5273 9336
rect 5307 9364 5319 9367
rect 5626 9364 5632 9376
rect 5307 9336 5632 9364
rect 5307 9333 5319 9336
rect 5261 9327 5319 9333
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 6181 9367 6239 9373
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 8110 9364 8116 9376
rect 6227 9336 8116 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 1104 9274 11316 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 11316 9274
rect 1104 9200 11316 9222
rect 5258 9120 5264 9172
rect 5316 9160 5322 9172
rect 6914 9160 6920 9172
rect 5316 9132 6920 9160
rect 5316 9120 5322 9132
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 3786 9052 3792 9104
rect 3844 9092 3850 9104
rect 3844 9064 4200 9092
rect 3844 9052 3850 9064
rect 1670 8984 1676 9036
rect 1728 9024 1734 9036
rect 4062 9024 4068 9036
rect 1728 8996 4068 9024
rect 1728 8984 1734 8996
rect 4062 8984 4068 8996
rect 4120 8984 4126 9036
rect 4172 9024 4200 9064
rect 4890 9052 4896 9104
rect 4948 9092 4954 9104
rect 7009 9095 7067 9101
rect 7009 9092 7021 9095
rect 4948 9064 7021 9092
rect 4948 9052 4954 9064
rect 7009 9061 7021 9064
rect 7055 9061 7067 9095
rect 7009 9055 7067 9061
rect 5718 9024 5724 9036
rect 4172 8996 5724 9024
rect 5718 8984 5724 8996
rect 5776 8984 5782 9036
rect 7466 8984 7472 9036
rect 7524 9024 7530 9036
rect 8941 9027 8999 9033
rect 8941 9024 8953 9027
rect 7524 8996 8953 9024
rect 7524 8984 7530 8996
rect 8941 8993 8953 8996
rect 8987 8993 8999 9027
rect 8941 8987 8999 8993
rect 1026 8916 1032 8968
rect 1084 8956 1090 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 1084 8928 1409 8956
rect 1084 8916 1090 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 5350 8916 5356 8968
rect 5408 8956 5414 8968
rect 5994 8956 6000 8968
rect 5408 8928 6000 8956
rect 5408 8916 5414 8928
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 8754 8916 8760 8968
rect 8812 8916 8818 8968
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8956 9275 8959
rect 9950 8956 9956 8968
rect 9263 8928 9956 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 1946 8848 1952 8900
rect 2004 8848 2010 8900
rect 3878 8888 3884 8900
rect 3174 8860 3884 8888
rect 3878 8848 3884 8860
rect 3936 8848 3942 8900
rect 8018 8848 8024 8900
rect 8076 8888 8082 8900
rect 8076 8860 8156 8888
rect 8076 8848 8082 8860
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 3326 8820 3332 8832
rect 1627 8792 3332 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 3326 8780 3332 8792
rect 3384 8780 3390 8832
rect 3418 8780 3424 8832
rect 3476 8780 3482 8832
rect 8128 8820 8156 8860
rect 8202 8848 8208 8900
rect 8260 8888 8266 8900
rect 8481 8891 8539 8897
rect 8481 8888 8493 8891
rect 8260 8860 8493 8888
rect 8260 8848 8266 8860
rect 8481 8857 8493 8860
rect 8527 8857 8539 8891
rect 8481 8851 8539 8857
rect 9232 8820 9260 8919
rect 9950 8916 9956 8928
rect 10008 8916 10014 8968
rect 8128 8792 9260 8820
rect 1104 8730 11316 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 11316 8730
rect 1104 8656 11316 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 1627 8588 1900 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 1026 8508 1032 8560
rect 1084 8548 1090 8560
rect 1673 8551 1731 8557
rect 1673 8548 1685 8551
rect 1084 8520 1685 8548
rect 1084 8508 1090 8520
rect 1673 8517 1685 8520
rect 1719 8517 1731 8551
rect 1872 8548 1900 8588
rect 1946 8576 1952 8628
rect 2004 8616 2010 8628
rect 2409 8619 2467 8625
rect 2409 8616 2421 8619
rect 2004 8588 2421 8616
rect 2004 8576 2010 8588
rect 2409 8585 2421 8588
rect 2455 8585 2467 8619
rect 2409 8579 2467 8585
rect 2777 8619 2835 8625
rect 2777 8585 2789 8619
rect 2823 8616 2835 8619
rect 3418 8616 3424 8628
rect 2823 8588 3424 8616
rect 2823 8585 2835 8588
rect 2777 8579 2835 8585
rect 3418 8576 3424 8588
rect 3476 8576 3482 8628
rect 5534 8576 5540 8628
rect 5592 8576 5598 8628
rect 6638 8576 6644 8628
rect 6696 8616 6702 8628
rect 8113 8619 8171 8625
rect 8113 8616 8125 8619
rect 6696 8588 8125 8616
rect 6696 8576 6702 8588
rect 8113 8585 8125 8588
rect 8159 8585 8171 8619
rect 8113 8579 8171 8585
rect 8294 8576 8300 8628
rect 8352 8616 8358 8628
rect 8941 8619 8999 8625
rect 8941 8616 8953 8619
rect 8352 8588 8953 8616
rect 8352 8576 8358 8588
rect 8941 8585 8953 8588
rect 8987 8585 8999 8619
rect 8941 8579 8999 8585
rect 2958 8548 2964 8560
rect 1872 8520 2964 8548
rect 1673 8511 1731 8517
rect 2958 8508 2964 8520
rect 3016 8508 3022 8560
rect 5445 8551 5503 8557
rect 5445 8517 5457 8551
rect 5491 8548 5503 8551
rect 5552 8548 5580 8576
rect 6730 8548 6736 8560
rect 5491 8520 5580 8548
rect 6380 8520 6736 8548
rect 5491 8517 5503 8520
rect 5445 8511 5503 8517
rect 1302 8440 1308 8492
rect 1360 8480 1366 8492
rect 1397 8483 1455 8489
rect 1397 8480 1409 8483
rect 1360 8452 1409 8480
rect 1360 8440 1366 8452
rect 1397 8449 1409 8452
rect 1443 8480 1455 8483
rect 1857 8483 1915 8489
rect 1857 8480 1869 8483
rect 1443 8452 1869 8480
rect 1443 8449 1455 8452
rect 1397 8443 1455 8449
rect 1857 8449 1869 8452
rect 1903 8449 1915 8483
rect 1857 8443 1915 8449
rect 3326 8440 3332 8492
rect 3384 8480 3390 8492
rect 5215 8483 5273 8489
rect 5215 8480 5227 8483
rect 3384 8452 5227 8480
rect 3384 8440 3390 8452
rect 5215 8449 5227 8452
rect 5261 8449 5273 8483
rect 5215 8443 5273 8449
rect 5350 8440 5356 8492
rect 5408 8440 5414 8492
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8480 5595 8483
rect 5718 8480 5724 8492
rect 5583 8452 5724 8480
rect 5583 8449 5595 8452
rect 5537 8443 5595 8449
rect 5718 8440 5724 8452
rect 5776 8440 5782 8492
rect 6380 8489 6408 8520
rect 6730 8508 6736 8520
rect 6788 8508 6794 8560
rect 7650 8508 7656 8560
rect 7708 8508 7714 8560
rect 9306 8548 9312 8560
rect 8496 8520 9312 8548
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 7926 8440 7932 8492
rect 7984 8480 7990 8492
rect 8496 8489 8524 8520
rect 9306 8508 9312 8520
rect 9364 8508 9370 8560
rect 8205 8483 8263 8489
rect 8205 8480 8217 8483
rect 7984 8452 8217 8480
rect 7984 8440 7990 8452
rect 8205 8449 8217 8452
rect 8251 8449 8263 8483
rect 8205 8443 8263 8449
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8449 8539 8483
rect 8481 8443 8539 8449
rect 8662 8440 8668 8492
rect 8720 8480 8726 8492
rect 8757 8483 8815 8489
rect 8757 8480 8769 8483
rect 8720 8452 8769 8480
rect 8720 8440 8726 8452
rect 8757 8449 8769 8452
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 2866 8372 2872 8424
rect 2924 8372 2930 8424
rect 2961 8415 3019 8421
rect 2961 8381 2973 8415
rect 3007 8381 3019 8415
rect 2961 8375 3019 8381
rect 2590 8236 2596 8288
rect 2648 8276 2654 8288
rect 2976 8276 3004 8375
rect 3142 8372 3148 8424
rect 3200 8412 3206 8424
rect 5077 8415 5135 8421
rect 5077 8412 5089 8415
rect 3200 8384 5089 8412
rect 3200 8372 3206 8384
rect 5077 8381 5089 8384
rect 5123 8412 5135 8415
rect 5626 8412 5632 8424
rect 5123 8384 5632 8412
rect 5123 8381 5135 8384
rect 5077 8375 5135 8381
rect 5626 8372 5632 8384
rect 5684 8412 5690 8424
rect 6178 8412 6184 8424
rect 5684 8384 6184 8412
rect 5684 8372 5690 8384
rect 6178 8372 6184 8384
rect 6236 8372 6242 8424
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 6730 8412 6736 8424
rect 6687 8384 6736 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 6730 8372 6736 8384
rect 6788 8372 6794 8424
rect 7834 8304 7840 8356
rect 7892 8344 7898 8356
rect 8202 8344 8208 8356
rect 7892 8316 8208 8344
rect 7892 8304 7898 8316
rect 8202 8304 8208 8316
rect 8260 8344 8266 8356
rect 8665 8347 8723 8353
rect 8665 8344 8677 8347
rect 8260 8316 8677 8344
rect 8260 8304 8266 8316
rect 8665 8313 8677 8316
rect 8711 8313 8723 8347
rect 8665 8307 8723 8313
rect 4706 8276 4712 8288
rect 2648 8248 4712 8276
rect 2648 8236 2654 8248
rect 4706 8236 4712 8248
rect 4764 8276 4770 8288
rect 5258 8276 5264 8288
rect 4764 8248 5264 8276
rect 4764 8236 4770 8248
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 5721 8279 5779 8285
rect 5721 8245 5733 8279
rect 5767 8276 5779 8279
rect 6362 8276 6368 8288
rect 5767 8248 6368 8276
rect 5767 8245 5779 8248
rect 5721 8239 5779 8245
rect 6362 8236 6368 8248
rect 6420 8236 6426 8288
rect 1104 8186 11316 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 11316 8186
rect 1104 8112 11316 8134
rect 2501 8075 2559 8081
rect 2501 8041 2513 8075
rect 2547 8072 2559 8075
rect 2866 8072 2872 8084
rect 2547 8044 2872 8072
rect 2547 8041 2559 8044
rect 2501 8035 2559 8041
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 6730 8032 6736 8084
rect 6788 8072 6794 8084
rect 6825 8075 6883 8081
rect 6825 8072 6837 8075
rect 6788 8044 6837 8072
rect 6788 8032 6794 8044
rect 6825 8041 6837 8044
rect 6871 8041 6883 8075
rect 6825 8035 6883 8041
rect 2774 7964 2780 8016
rect 2832 7964 2838 8016
rect 6638 8004 6644 8016
rect 5368 7976 6644 8004
rect 1302 7828 1308 7880
rect 1360 7868 1366 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 1360 7840 1409 7868
rect 1360 7828 1366 7840
rect 1397 7837 1409 7840
rect 1443 7868 1455 7871
rect 1765 7871 1823 7877
rect 1765 7868 1777 7871
rect 1443 7840 1777 7868
rect 1443 7837 1455 7840
rect 1397 7831 1455 7837
rect 1765 7837 1777 7840
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 2682 7828 2688 7880
rect 2740 7828 2746 7880
rect 2792 7877 2820 7964
rect 4062 7896 4068 7948
rect 4120 7936 4126 7948
rect 5368 7936 5396 7976
rect 6638 7964 6644 7976
rect 6696 7964 6702 8016
rect 4120 7908 5396 7936
rect 4120 7896 4126 7908
rect 6270 7896 6276 7948
rect 6328 7896 6334 7948
rect 6362 7896 6368 7948
rect 6420 7896 6426 7948
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7837 2835 7871
rect 2777 7831 2835 7837
rect 3142 7828 3148 7880
rect 3200 7828 3206 7880
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7868 6515 7871
rect 6546 7868 6552 7880
rect 6503 7840 6552 7868
rect 6503 7837 6515 7840
rect 6457 7831 6515 7837
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 2869 7803 2927 7809
rect 2869 7769 2881 7803
rect 2915 7769 2927 7803
rect 2869 7763 2927 7769
rect 1578 7692 1584 7744
rect 1636 7692 1642 7744
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 2884 7732 2912 7763
rect 2958 7760 2964 7812
rect 3016 7809 3022 7812
rect 3016 7803 3045 7809
rect 3033 7769 3045 7803
rect 3016 7763 3045 7769
rect 3016 7760 3022 7763
rect 4338 7760 4344 7812
rect 4396 7760 4402 7812
rect 4448 7772 4830 7800
rect 2832 7704 2912 7732
rect 2832 7692 2838 7704
rect 3878 7692 3884 7744
rect 3936 7732 3942 7744
rect 4448 7732 4476 7772
rect 3936 7704 4476 7732
rect 3936 7692 3942 7704
rect 5350 7692 5356 7744
rect 5408 7732 5414 7744
rect 5813 7735 5871 7741
rect 5813 7732 5825 7735
rect 5408 7704 5825 7732
rect 5408 7692 5414 7704
rect 5813 7701 5825 7704
rect 5859 7701 5871 7735
rect 5813 7695 5871 7701
rect 1104 7642 11316 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 11316 7642
rect 1104 7568 11316 7590
rect 1578 7488 1584 7540
rect 1636 7528 1642 7540
rect 1636 7500 4292 7528
rect 1636 7488 1642 7500
rect 1670 7460 1676 7472
rect 1412 7432 1676 7460
rect 1412 7401 1440 7432
rect 1670 7420 1676 7432
rect 1728 7420 1734 7472
rect 3878 7460 3884 7472
rect 2898 7432 3884 7460
rect 3878 7420 3884 7432
rect 3936 7420 3942 7472
rect 4264 7460 4292 7500
rect 4338 7488 4344 7540
rect 4396 7528 4402 7540
rect 4709 7531 4767 7537
rect 4709 7528 4721 7531
rect 4396 7500 4721 7528
rect 4396 7488 4402 7500
rect 4709 7497 4721 7500
rect 4755 7497 4767 7531
rect 4709 7491 4767 7497
rect 5077 7531 5135 7537
rect 5077 7497 5089 7531
rect 5123 7528 5135 7531
rect 5350 7528 5356 7540
rect 5123 7500 5356 7528
rect 5123 7497 5135 7500
rect 5077 7491 5135 7497
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 6023 7463 6081 7469
rect 6023 7460 6035 7463
rect 4264 7432 6035 7460
rect 6023 7429 6035 7432
rect 6069 7429 6081 7463
rect 6023 7423 6081 7429
rect 8110 7420 8116 7472
rect 8168 7460 8174 7472
rect 9493 7463 9551 7469
rect 9493 7460 9505 7463
rect 8168 7432 9505 7460
rect 8168 7420 8174 7432
rect 9493 7429 9505 7432
rect 9539 7429 9551 7463
rect 9493 7423 9551 7429
rect 9950 7420 9956 7472
rect 10008 7420 10014 7472
rect 1397 7395 1455 7401
rect 1397 7361 1409 7395
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 3421 7395 3479 7401
rect 3421 7361 3433 7395
rect 3467 7361 3479 7395
rect 3421 7355 3479 7361
rect 1670 7284 1676 7336
rect 1728 7284 1734 7336
rect 3436 7268 3464 7355
rect 3510 7352 3516 7404
rect 3568 7352 3574 7404
rect 3602 7352 3608 7404
rect 3660 7352 3666 7404
rect 3694 7352 3700 7404
rect 3752 7401 3758 7404
rect 3752 7395 3781 7401
rect 3769 7361 3781 7395
rect 3752 7355 3781 7361
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7392 5227 7395
rect 5537 7395 5595 7401
rect 5537 7392 5549 7395
rect 5215 7364 5549 7392
rect 5215 7361 5227 7364
rect 5169 7355 5227 7361
rect 5537 7361 5549 7364
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 3752 7352 3758 7355
rect 3878 7284 3884 7336
rect 3936 7284 3942 7336
rect 5258 7284 5264 7336
rect 5316 7284 5322 7336
rect 2958 7216 2964 7268
rect 3016 7256 3022 7268
rect 3237 7259 3295 7265
rect 3237 7256 3249 7259
rect 3016 7228 3249 7256
rect 3016 7216 3022 7228
rect 3237 7225 3249 7228
rect 3283 7225 3295 7259
rect 3237 7219 3295 7225
rect 3418 7216 3424 7268
rect 3476 7256 3482 7268
rect 5736 7256 5764 7355
rect 3476 7228 5764 7256
rect 3476 7216 3482 7228
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 3050 7188 3056 7200
rect 2832 7160 3056 7188
rect 2832 7148 2838 7160
rect 3050 7148 3056 7160
rect 3108 7188 3114 7200
rect 3145 7191 3203 7197
rect 3145 7188 3157 7191
rect 3108 7160 3157 7188
rect 3108 7148 3114 7160
rect 3145 7157 3157 7160
rect 3191 7157 3203 7191
rect 3145 7151 3203 7157
rect 3510 7148 3516 7200
rect 3568 7188 3574 7200
rect 4062 7188 4068 7200
rect 3568 7160 4068 7188
rect 3568 7148 3574 7160
rect 4062 7148 4068 7160
rect 4120 7188 4126 7200
rect 5828 7188 5856 7355
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 6178 7352 6184 7404
rect 6236 7352 6242 7404
rect 8754 7352 8760 7404
rect 8812 7392 8818 7404
rect 9217 7395 9275 7401
rect 9217 7392 9229 7395
rect 8812 7364 9229 7392
rect 8812 7352 8818 7364
rect 9217 7361 9229 7364
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 4120 7160 5856 7188
rect 4120 7148 4126 7160
rect 10962 7148 10968 7200
rect 11020 7148 11026 7200
rect 1104 7098 11316 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 11316 7098
rect 1104 7024 11316 7046
rect 1670 6944 1676 6996
rect 1728 6984 1734 6996
rect 2225 6987 2283 6993
rect 2225 6984 2237 6987
rect 1728 6956 2237 6984
rect 1728 6944 1734 6956
rect 2225 6953 2237 6956
rect 2271 6953 2283 6987
rect 2225 6947 2283 6953
rect 3237 6987 3295 6993
rect 3237 6953 3249 6987
rect 3283 6984 3295 6987
rect 3418 6984 3424 6996
rect 3283 6956 3424 6984
rect 3283 6953 3295 6956
rect 3237 6947 3295 6953
rect 3418 6944 3424 6956
rect 3476 6944 3482 6996
rect 1581 6919 1639 6925
rect 1581 6885 1593 6919
rect 1627 6914 1639 6919
rect 3694 6916 3700 6928
rect 1627 6886 1661 6914
rect 2608 6888 3700 6916
rect 1627 6885 1639 6886
rect 1581 6879 1639 6885
rect 1596 6848 1624 6879
rect 2608 6848 2636 6888
rect 3694 6876 3700 6888
rect 3752 6876 3758 6928
rect 2777 6851 2835 6857
rect 2777 6848 2789 6851
rect 1596 6820 2636 6848
rect 2700 6820 2789 6848
rect 2700 6792 2728 6820
rect 2777 6817 2789 6820
rect 2823 6817 2835 6851
rect 2777 6811 2835 6817
rect 6638 6808 6644 6860
rect 6696 6808 6702 6860
rect 10778 6808 10784 6860
rect 10836 6808 10842 6860
rect 1210 6740 1216 6792
rect 1268 6780 1274 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 1268 6752 1409 6780
rect 1268 6740 1274 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6749 1731 6783
rect 1673 6743 1731 6749
rect 1302 6672 1308 6724
rect 1360 6712 1366 6724
rect 1688 6712 1716 6743
rect 2682 6740 2688 6792
rect 2740 6740 2746 6792
rect 2866 6740 2872 6792
rect 2924 6780 2930 6792
rect 3145 6783 3203 6789
rect 3145 6780 3157 6783
rect 2924 6752 3157 6780
rect 2924 6740 2930 6752
rect 3145 6749 3157 6752
rect 3191 6780 3203 6783
rect 5718 6780 5724 6792
rect 3191 6752 5724 6780
rect 3191 6749 3203 6752
rect 3145 6743 3203 6749
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 10962 6740 10968 6792
rect 11020 6740 11026 6792
rect 1949 6715 2007 6721
rect 1949 6712 1961 6715
rect 1360 6684 1961 6712
rect 1360 6672 1366 6684
rect 1949 6681 1961 6684
rect 1995 6681 2007 6715
rect 1949 6675 2007 6681
rect 2593 6715 2651 6721
rect 2593 6681 2605 6715
rect 2639 6712 2651 6715
rect 3050 6712 3056 6724
rect 2639 6684 3056 6712
rect 2639 6681 2651 6684
rect 2593 6675 2651 6681
rect 3050 6672 3056 6684
rect 3108 6672 3114 6724
rect 4801 6715 4859 6721
rect 4801 6681 4813 6715
rect 4847 6681 4859 6715
rect 4801 6675 4859 6681
rect 1854 6604 1860 6656
rect 1912 6604 1918 6656
rect 2685 6647 2743 6653
rect 2685 6613 2697 6647
rect 2731 6644 2743 6647
rect 2958 6644 2964 6656
rect 2731 6616 2964 6644
rect 2731 6613 2743 6616
rect 2685 6607 2743 6613
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 4614 6604 4620 6656
rect 4672 6644 4678 6656
rect 4816 6644 4844 6675
rect 6914 6672 6920 6724
rect 6972 6672 6978 6724
rect 7650 6672 7656 6724
rect 7708 6672 7714 6724
rect 4672 6616 4844 6644
rect 4672 6604 4678 6616
rect 5442 6604 5448 6656
rect 5500 6644 5506 6656
rect 6089 6647 6147 6653
rect 6089 6644 6101 6647
rect 5500 6616 6101 6644
rect 5500 6604 5506 6616
rect 6089 6613 6101 6616
rect 6135 6613 6147 6647
rect 6089 6607 6147 6613
rect 7926 6604 7932 6656
rect 7984 6644 7990 6656
rect 8389 6647 8447 6653
rect 8389 6644 8401 6647
rect 7984 6616 8401 6644
rect 7984 6604 7990 6616
rect 8389 6613 8401 6616
rect 8435 6613 8447 6647
rect 8389 6607 8447 6613
rect 1104 6554 11316 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 11316 6554
rect 1104 6480 11316 6502
rect 1210 6400 1216 6452
rect 1268 6400 1274 6452
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 2774 6440 2780 6452
rect 1627 6412 2780 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 2774 6400 2780 6412
rect 2832 6400 2838 6452
rect 3878 6400 3884 6452
rect 3936 6440 3942 6452
rect 3936 6412 6684 6440
rect 3936 6400 3942 6412
rect 1228 6372 1256 6400
rect 1673 6375 1731 6381
rect 1673 6372 1685 6375
rect 1228 6344 1685 6372
rect 1673 6341 1685 6344
rect 1719 6341 1731 6375
rect 1673 6335 1731 6341
rect 3142 6332 3148 6384
rect 3200 6332 3206 6384
rect 3970 6332 3976 6384
rect 4028 6372 4034 6384
rect 4028 6344 5198 6372
rect 4028 6332 4034 6344
rect 1210 6264 1216 6316
rect 1268 6304 1274 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 1268 6276 1409 6304
rect 1268 6264 1274 6276
rect 1397 6273 1409 6276
rect 1443 6304 1455 6307
rect 1857 6307 1915 6313
rect 1857 6304 1869 6307
rect 1443 6276 1869 6304
rect 1443 6273 1455 6276
rect 1397 6267 1455 6273
rect 1857 6273 1869 6276
rect 1903 6273 1915 6307
rect 1857 6267 1915 6273
rect 5994 6264 6000 6316
rect 6052 6304 6058 6316
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 6052 6276 6377 6304
rect 6052 6264 6058 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 6454 6264 6460 6316
rect 6512 6304 6518 6316
rect 6656 6313 6684 6412
rect 6914 6400 6920 6452
rect 6972 6440 6978 6452
rect 7377 6443 7435 6449
rect 7377 6440 7389 6443
rect 6972 6412 7389 6440
rect 6972 6400 6978 6412
rect 7377 6409 7389 6412
rect 7423 6409 7435 6443
rect 7377 6403 7435 6409
rect 8018 6400 8024 6452
rect 8076 6440 8082 6452
rect 8076 6412 8984 6440
rect 8076 6400 8082 6412
rect 8757 6375 8815 6381
rect 8757 6372 8769 6375
rect 8036 6344 8769 6372
rect 6641 6307 6699 6313
rect 6641 6304 6653 6307
rect 6512 6276 6653 6304
rect 6512 6264 6518 6276
rect 6641 6273 6653 6276
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6304 7619 6307
rect 7742 6304 7748 6316
rect 7607 6276 7748 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 2133 6239 2191 6245
rect 2133 6205 2145 6239
rect 2179 6205 2191 6239
rect 2133 6199 2191 6205
rect 1394 6128 1400 6180
rect 1452 6168 1458 6180
rect 2148 6168 2176 6199
rect 2406 6196 2412 6248
rect 2464 6196 2470 6248
rect 4433 6239 4491 6245
rect 4433 6205 4445 6239
rect 4479 6205 4491 6239
rect 4433 6199 4491 6205
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6236 4767 6239
rect 4798 6236 4804 6248
rect 4755 6208 4804 6236
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 1452 6140 2176 6168
rect 1452 6128 1458 6140
rect 2958 6060 2964 6112
rect 3016 6100 3022 6112
rect 3602 6100 3608 6112
rect 3016 6072 3608 6100
rect 3016 6060 3022 6072
rect 3602 6060 3608 6072
rect 3660 6100 3666 6112
rect 3881 6103 3939 6109
rect 3881 6100 3893 6103
rect 3660 6072 3893 6100
rect 3660 6060 3666 6072
rect 3881 6069 3893 6072
rect 3927 6069 3939 6103
rect 4448 6100 4476 6199
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 4706 6100 4712 6112
rect 4448 6072 4712 6100
rect 3881 6063 3939 6069
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 5902 6060 5908 6112
rect 5960 6100 5966 6112
rect 6181 6103 6239 6109
rect 6181 6100 6193 6103
rect 5960 6072 6193 6100
rect 5960 6060 5966 6072
rect 6181 6069 6193 6072
rect 6227 6069 6239 6103
rect 7576 6100 7604 6267
rect 7742 6264 7748 6276
rect 7800 6264 7806 6316
rect 7834 6264 7840 6316
rect 7892 6264 7898 6316
rect 7926 6264 7932 6316
rect 7984 6304 7990 6316
rect 8036 6313 8064 6344
rect 8757 6341 8769 6344
rect 8803 6341 8815 6375
rect 8757 6335 8815 6341
rect 8021 6307 8079 6313
rect 8021 6304 8033 6307
rect 7984 6276 8033 6304
rect 7984 6264 7990 6276
rect 8021 6273 8033 6276
rect 8067 6273 8079 6307
rect 8021 6267 8079 6273
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 8481 6307 8539 6313
rect 8251 6276 8432 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 7653 6239 7711 6245
rect 7653 6205 7665 6239
rect 7699 6236 7711 6239
rect 8113 6239 8171 6245
rect 8113 6236 8125 6239
rect 7699 6208 8125 6236
rect 7699 6205 7711 6208
rect 7653 6199 7711 6205
rect 8113 6205 8125 6208
rect 8159 6236 8171 6239
rect 8294 6236 8300 6248
rect 8159 6208 8300 6236
rect 8159 6205 8171 6208
rect 8113 6199 8171 6205
rect 8294 6196 8300 6208
rect 8352 6196 8358 6248
rect 8404 6236 8432 6276
rect 8481 6273 8493 6307
rect 8527 6304 8539 6307
rect 8846 6304 8852 6316
rect 8527 6276 8852 6304
rect 8527 6273 8539 6276
rect 8481 6267 8539 6273
rect 8846 6264 8852 6276
rect 8904 6264 8910 6316
rect 8956 6313 8984 6412
rect 9309 6375 9367 6381
rect 9309 6341 9321 6375
rect 9355 6372 9367 6375
rect 10962 6372 10968 6384
rect 9355 6344 10968 6372
rect 9355 6341 9367 6344
rect 9309 6335 9367 6341
rect 8941 6307 8999 6313
rect 8941 6273 8953 6307
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 8570 6236 8576 6248
rect 8404 6208 8576 6236
rect 8570 6196 8576 6208
rect 8628 6196 8634 6248
rect 9324 6236 9352 6335
rect 10962 6332 10968 6344
rect 11020 6332 11026 6384
rect 8772 6208 9352 6236
rect 7742 6128 7748 6180
rect 7800 6128 7806 6180
rect 8110 6100 8116 6112
rect 7576 6072 8116 6100
rect 6181 6063 6239 6069
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 8297 6103 8355 6109
rect 8297 6069 8309 6103
rect 8343 6100 8355 6103
rect 8386 6100 8392 6112
rect 8343 6072 8392 6100
rect 8343 6069 8355 6072
rect 8297 6063 8355 6069
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 8662 6060 8668 6112
rect 8720 6100 8726 6112
rect 8772 6109 8800 6208
rect 8757 6103 8815 6109
rect 8757 6100 8769 6103
rect 8720 6072 8769 6100
rect 8720 6060 8726 6072
rect 8757 6069 8769 6072
rect 8803 6069 8815 6103
rect 8757 6063 8815 6069
rect 9306 6060 9312 6112
rect 9364 6060 9370 6112
rect 9490 6060 9496 6112
rect 9548 6060 9554 6112
rect 1104 6010 11316 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 11316 6010
rect 1104 5936 11316 5958
rect 2406 5856 2412 5908
rect 2464 5896 2470 5908
rect 2593 5899 2651 5905
rect 2593 5896 2605 5899
rect 2464 5868 2605 5896
rect 2464 5856 2470 5868
rect 2593 5865 2605 5868
rect 2639 5865 2651 5899
rect 2593 5859 2651 5865
rect 4798 5856 4804 5908
rect 4856 5896 4862 5908
rect 4985 5899 5043 5905
rect 4985 5896 4997 5899
rect 4856 5868 4997 5896
rect 4856 5856 4862 5868
rect 4985 5865 4997 5868
rect 5031 5865 5043 5899
rect 8846 5896 8852 5908
rect 4985 5859 5043 5865
rect 7852 5868 8852 5896
rect 1581 5831 1639 5837
rect 1581 5797 1593 5831
rect 1627 5828 1639 5831
rect 6638 5828 6644 5840
rect 1627 5800 6644 5828
rect 1627 5797 1639 5800
rect 1581 5791 1639 5797
rect 6638 5788 6644 5800
rect 6696 5788 6702 5840
rect 2866 5720 2872 5772
rect 2924 5760 2930 5772
rect 3234 5760 3240 5772
rect 2924 5732 3240 5760
rect 2924 5720 2930 5732
rect 3234 5720 3240 5732
rect 3292 5760 3298 5772
rect 5258 5760 5264 5772
rect 3292 5732 5264 5760
rect 3292 5720 3298 5732
rect 5258 5720 5264 5732
rect 5316 5760 5322 5772
rect 5537 5763 5595 5769
rect 5537 5760 5549 5763
rect 5316 5732 5549 5760
rect 5316 5720 5322 5732
rect 5537 5729 5549 5732
rect 5583 5729 5595 5763
rect 5537 5723 5595 5729
rect 5718 5720 5724 5772
rect 5776 5760 5782 5772
rect 5776 5732 6040 5760
rect 5776 5720 5782 5732
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 1397 5695 1455 5701
rect 1397 5692 1409 5695
rect 1360 5664 1409 5692
rect 1360 5652 1366 5664
rect 1397 5661 1409 5664
rect 1443 5692 1455 5695
rect 1673 5695 1731 5701
rect 1673 5692 1685 5695
rect 1443 5664 1685 5692
rect 1443 5661 1455 5664
rect 1397 5655 1455 5661
rect 1673 5661 1685 5664
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 2958 5652 2964 5704
rect 3016 5652 3022 5704
rect 5353 5695 5411 5701
rect 5353 5661 5365 5695
rect 5399 5692 5411 5695
rect 5902 5692 5908 5704
rect 5399 5664 5908 5692
rect 5399 5661 5411 5664
rect 5353 5655 5411 5661
rect 5902 5652 5908 5664
rect 5960 5652 5966 5704
rect 6012 5701 6040 5732
rect 6454 5720 6460 5772
rect 6512 5720 6518 5772
rect 5997 5695 6055 5701
rect 5997 5661 6009 5695
rect 6043 5661 6055 5695
rect 5997 5655 6055 5661
rect 7561 5695 7619 5701
rect 7561 5661 7573 5695
rect 7607 5692 7619 5695
rect 7852 5692 7880 5868
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 9030 5856 9036 5908
rect 9088 5896 9094 5908
rect 9306 5896 9312 5908
rect 9088 5868 9312 5896
rect 9088 5856 9094 5868
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 7929 5831 7987 5837
rect 7929 5797 7941 5831
rect 7975 5828 7987 5831
rect 8294 5828 8300 5840
rect 7975 5800 8300 5828
rect 7975 5797 7987 5800
rect 7929 5791 7987 5797
rect 8294 5788 8300 5800
rect 8352 5828 8358 5840
rect 8478 5828 8484 5840
rect 8352 5800 8484 5828
rect 8352 5788 8358 5800
rect 8478 5788 8484 5800
rect 8536 5788 8542 5840
rect 8662 5828 8668 5840
rect 8588 5800 8668 5828
rect 8018 5720 8024 5772
rect 8076 5720 8082 5772
rect 8588 5760 8616 5800
rect 8662 5788 8668 5800
rect 8720 5788 8726 5840
rect 9048 5828 9076 5856
rect 8864 5800 9076 5828
rect 8404 5732 8616 5760
rect 7607 5664 7880 5692
rect 7607 5661 7619 5664
rect 7561 5655 7619 5661
rect 1854 5584 1860 5636
rect 1912 5624 1918 5636
rect 1912 5596 5948 5624
rect 1912 5584 1918 5596
rect 3050 5516 3056 5568
rect 3108 5516 3114 5568
rect 5445 5559 5503 5565
rect 5445 5525 5457 5559
rect 5491 5556 5503 5559
rect 5813 5559 5871 5565
rect 5813 5556 5825 5559
rect 5491 5528 5825 5556
rect 5491 5525 5503 5528
rect 5445 5519 5503 5525
rect 5813 5525 5825 5528
rect 5859 5525 5871 5559
rect 5920 5556 5948 5596
rect 6086 5584 6092 5636
rect 6144 5584 6150 5636
rect 6178 5584 6184 5636
rect 6236 5584 6242 5636
rect 6299 5627 6357 5633
rect 6299 5624 6311 5627
rect 6288 5593 6311 5624
rect 6345 5593 6357 5627
rect 8036 5624 8064 5720
rect 8110 5652 8116 5704
rect 8168 5652 8174 5704
rect 8205 5695 8263 5701
rect 8205 5661 8217 5695
rect 8251 5692 8263 5695
rect 8294 5692 8300 5704
rect 8251 5664 8300 5692
rect 8251 5661 8263 5664
rect 8205 5655 8263 5661
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 8404 5701 8432 5732
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5661 8447 5695
rect 8389 5655 8447 5661
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5692 8631 5695
rect 8864 5692 8892 5800
rect 8941 5763 8999 5769
rect 8941 5729 8953 5763
rect 8987 5760 8999 5763
rect 9214 5760 9220 5772
rect 8987 5732 9220 5760
rect 8987 5729 8999 5732
rect 8941 5723 8999 5729
rect 9214 5720 9220 5732
rect 9272 5720 9278 5772
rect 8619 5664 8892 5692
rect 8619 5661 8631 5664
rect 8573 5655 8631 5661
rect 8481 5627 8539 5633
rect 8481 5624 8493 5627
rect 8036 5596 8493 5624
rect 6288 5587 6357 5593
rect 8481 5593 8493 5596
rect 8527 5593 8539 5627
rect 8481 5587 8539 5593
rect 6288 5556 6316 5587
rect 5920 5528 6316 5556
rect 8588 5556 8616 5655
rect 9217 5627 9275 5633
rect 9217 5593 9229 5627
rect 9263 5593 9275 5627
rect 9217 5587 9275 5593
rect 8662 5556 8668 5568
rect 8588 5528 8668 5556
rect 5813 5519 5871 5525
rect 8662 5516 8668 5528
rect 8720 5516 8726 5568
rect 8757 5559 8815 5565
rect 8757 5525 8769 5559
rect 8803 5556 8815 5559
rect 9232 5556 9260 5587
rect 9674 5584 9680 5636
rect 9732 5584 9738 5636
rect 8803 5528 9260 5556
rect 8803 5525 8815 5528
rect 8757 5519 8815 5525
rect 9306 5516 9312 5568
rect 9364 5556 9370 5568
rect 10689 5559 10747 5565
rect 10689 5556 10701 5559
rect 9364 5528 10701 5556
rect 9364 5516 9370 5528
rect 10689 5525 10701 5528
rect 10735 5525 10747 5559
rect 10689 5519 10747 5525
rect 1104 5466 11316 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 11316 5466
rect 1104 5392 11316 5414
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3237 5355 3295 5361
rect 3237 5352 3249 5355
rect 3108 5324 3249 5352
rect 3108 5312 3114 5324
rect 3237 5321 3249 5324
rect 3283 5321 3295 5355
rect 3237 5315 3295 5321
rect 3418 5312 3424 5364
rect 3476 5352 3482 5364
rect 3476 5324 6040 5352
rect 3476 5312 3482 5324
rect 2774 5293 2780 5296
rect 2751 5287 2780 5293
rect 2751 5253 2763 5287
rect 2751 5247 2780 5253
rect 2774 5244 2780 5247
rect 2832 5244 2838 5296
rect 2961 5287 3019 5293
rect 2961 5253 2973 5287
rect 3007 5284 3019 5287
rect 3326 5284 3332 5296
rect 3007 5256 3332 5284
rect 3007 5253 3019 5256
rect 2961 5247 3019 5253
rect 3326 5244 3332 5256
rect 3384 5284 3390 5296
rect 4062 5284 4068 5296
rect 3384 5256 4068 5284
rect 3384 5244 3390 5256
rect 4062 5244 4068 5256
rect 4120 5284 4126 5296
rect 4982 5284 4988 5296
rect 4120 5256 4988 5284
rect 4120 5244 4126 5256
rect 4982 5244 4988 5256
rect 5040 5244 5046 5296
rect 5718 5244 5724 5296
rect 5776 5244 5782 5296
rect 1210 5176 1216 5228
rect 1268 5216 1274 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 1268 5188 1409 5216
rect 1268 5176 1274 5188
rect 1397 5185 1409 5188
rect 1443 5216 1455 5219
rect 1673 5219 1731 5225
rect 1673 5216 1685 5219
rect 1443 5188 1685 5216
rect 1443 5185 1455 5188
rect 1397 5179 1455 5185
rect 1673 5185 1685 5188
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 2866 5176 2872 5228
rect 2924 5176 2930 5228
rect 3050 5176 3056 5228
rect 3108 5216 3114 5228
rect 3418 5216 3424 5228
rect 3108 5188 3424 5216
rect 3108 5176 3114 5188
rect 3418 5176 3424 5188
rect 3476 5176 3482 5228
rect 6012 5216 6040 5324
rect 6638 5312 6644 5364
rect 6696 5352 6702 5364
rect 6696 5324 6868 5352
rect 6696 5312 6702 5324
rect 6270 5244 6276 5296
rect 6328 5284 6334 5296
rect 6840 5293 6868 5324
rect 7742 5312 7748 5364
rect 7800 5312 7806 5364
rect 8294 5312 8300 5364
rect 8352 5352 8358 5364
rect 8389 5355 8447 5361
rect 8389 5352 8401 5355
rect 8352 5324 8401 5352
rect 8352 5312 8358 5324
rect 8389 5321 8401 5324
rect 8435 5321 8447 5355
rect 8389 5315 8447 5321
rect 8573 5355 8631 5361
rect 8573 5321 8585 5355
rect 8619 5352 8631 5355
rect 8846 5352 8852 5364
rect 8619 5324 8852 5352
rect 8619 5321 8631 5324
rect 8573 5315 8631 5321
rect 8846 5312 8852 5324
rect 8904 5352 8910 5364
rect 9306 5352 9312 5364
rect 8904 5324 9312 5352
rect 8904 5312 8910 5324
rect 9306 5312 9312 5324
rect 9364 5312 9370 5364
rect 9674 5312 9680 5364
rect 9732 5312 9738 5364
rect 10962 5312 10968 5364
rect 11020 5312 11026 5364
rect 6733 5287 6791 5293
rect 6733 5284 6745 5287
rect 6328 5256 6745 5284
rect 6328 5244 6334 5256
rect 6733 5253 6745 5256
rect 6779 5253 6791 5287
rect 6840 5287 6909 5293
rect 6840 5256 6863 5287
rect 6733 5247 6791 5253
rect 6851 5253 6863 5256
rect 6897 5253 6909 5287
rect 6851 5247 6909 5253
rect 7484 5256 8432 5284
rect 7484 5225 7512 5256
rect 8404 5228 8432 5256
rect 9490 5244 9496 5296
rect 9548 5244 9554 5296
rect 9692 5284 9720 5312
rect 9692 5256 9982 5284
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 6012 5188 6561 5216
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 2593 5151 2651 5157
rect 2593 5117 2605 5151
rect 2639 5148 2651 5151
rect 3878 5148 3884 5160
rect 2639 5120 3884 5148
rect 2639 5117 2651 5120
rect 2593 5111 2651 5117
rect 3878 5108 3884 5120
rect 3936 5108 3942 5160
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5148 4491 5151
rect 4709 5151 4767 5157
rect 4479 5120 4568 5148
rect 4479 5117 4491 5120
rect 4433 5111 4491 5117
rect 1394 5040 1400 5092
rect 1452 5080 1458 5092
rect 4540 5080 4568 5120
rect 4709 5117 4721 5151
rect 4755 5148 4767 5151
rect 4798 5148 4804 5160
rect 4755 5120 4804 5148
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 4798 5108 4804 5120
rect 4856 5108 4862 5160
rect 5074 5108 5080 5160
rect 5132 5148 5138 5160
rect 6656 5148 6684 5179
rect 7926 5176 7932 5228
rect 7984 5176 7990 5228
rect 8386 5176 8392 5228
rect 8444 5176 8450 5228
rect 8478 5176 8484 5228
rect 8536 5216 8542 5228
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8536 5188 8953 5216
rect 8536 5176 8542 5188
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 5132 5120 6684 5148
rect 7009 5151 7067 5157
rect 5132 5108 5138 5120
rect 7009 5117 7021 5151
rect 7055 5117 7067 5151
rect 7009 5111 7067 5117
rect 8113 5151 8171 5157
rect 8113 5117 8125 5151
rect 8159 5148 8171 5151
rect 8570 5148 8576 5160
rect 8159 5120 8576 5148
rect 8159 5117 8171 5120
rect 8113 5111 8171 5117
rect 1452 5052 4568 5080
rect 1452 5040 1458 5052
rect 1578 4972 1584 5024
rect 1636 4972 1642 5024
rect 4540 5012 4568 5052
rect 6454 5040 6460 5092
rect 6512 5080 6518 5092
rect 7024 5080 7052 5111
rect 8570 5108 8576 5120
rect 8628 5108 8634 5160
rect 9214 5108 9220 5160
rect 9272 5108 9278 5160
rect 6512 5052 7052 5080
rect 7653 5083 7711 5089
rect 6512 5040 6518 5052
rect 7653 5049 7665 5083
rect 7699 5080 7711 5083
rect 8478 5080 8484 5092
rect 7699 5052 8484 5080
rect 7699 5049 7711 5052
rect 7653 5043 7711 5049
rect 8478 5040 8484 5052
rect 8536 5080 8542 5092
rect 8754 5080 8760 5092
rect 8536 5052 8760 5080
rect 8536 5040 8542 5052
rect 8754 5040 8760 5052
rect 8812 5040 8818 5092
rect 4706 5012 4712 5024
rect 4540 4984 4712 5012
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 6178 4972 6184 5024
rect 6236 4972 6242 5024
rect 6362 4972 6368 5024
rect 6420 4972 6426 5024
rect 7374 4972 7380 5024
rect 7432 5012 7438 5024
rect 8573 5015 8631 5021
rect 8573 5012 8585 5015
rect 7432 4984 8585 5012
rect 7432 4972 7438 4984
rect 8573 4981 8585 4984
rect 8619 5012 8631 5015
rect 8662 5012 8668 5024
rect 8619 4984 8668 5012
rect 8619 4981 8631 4984
rect 8573 4975 8631 4981
rect 8662 4972 8668 4984
rect 8720 4972 8726 5024
rect 1104 4922 11316 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 11316 4922
rect 1104 4848 11316 4870
rect 2866 4768 2872 4820
rect 2924 4808 2930 4820
rect 3145 4811 3203 4817
rect 3145 4808 3157 4811
rect 2924 4780 3157 4808
rect 2924 4768 2930 4780
rect 3145 4777 3157 4780
rect 3191 4777 3203 4811
rect 3145 4771 3203 4777
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 8113 4811 8171 4817
rect 8113 4808 8125 4811
rect 7708 4780 8125 4808
rect 7708 4768 7714 4780
rect 8113 4777 8125 4780
rect 8159 4808 8171 4811
rect 9674 4808 9680 4820
rect 8159 4780 9680 4808
rect 8159 4777 8171 4780
rect 8113 4771 8171 4777
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 4062 4700 4068 4752
rect 4120 4740 4126 4752
rect 4157 4743 4215 4749
rect 4157 4740 4169 4743
rect 4120 4712 4169 4740
rect 4120 4700 4126 4712
rect 4157 4709 4169 4712
rect 4203 4709 4215 4743
rect 8297 4743 8355 4749
rect 8297 4740 8309 4743
rect 4157 4703 4215 4709
rect 7484 4712 8309 4740
rect 4706 4672 4712 4684
rect 4632 4644 4712 4672
rect 1394 4564 1400 4616
rect 1452 4564 1458 4616
rect 4632 4613 4660 4644
rect 4706 4632 4712 4644
rect 4764 4672 4770 4684
rect 4764 4644 6776 4672
rect 4764 4632 4770 4644
rect 6748 4616 6776 4644
rect 7374 4632 7380 4684
rect 7432 4632 7438 4684
rect 4617 4607 4675 4613
rect 4617 4573 4629 4607
rect 4663 4573 4675 4607
rect 4617 4567 4675 4573
rect 5077 4607 5135 4613
rect 5077 4573 5089 4607
rect 5123 4604 5135 4607
rect 5442 4604 5448 4616
rect 5123 4576 5448 4604
rect 5123 4573 5135 4576
rect 5077 4567 5135 4573
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 6730 4564 6736 4616
rect 6788 4564 6794 4616
rect 7484 4613 7512 4712
rect 8297 4709 8309 4712
rect 8343 4709 8355 4743
rect 8297 4703 8355 4709
rect 7561 4675 7619 4681
rect 7561 4641 7573 4675
rect 7607 4672 7619 4675
rect 8665 4675 8723 4681
rect 8665 4672 8677 4675
rect 7607 4644 8677 4672
rect 7607 4641 7619 4644
rect 7561 4635 7619 4641
rect 8665 4641 8677 4644
rect 8711 4641 8723 4675
rect 8665 4635 8723 4641
rect 7469 4607 7527 4613
rect 7469 4573 7481 4607
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 7653 4607 7711 4613
rect 7653 4573 7665 4607
rect 7699 4604 7711 4607
rect 8110 4604 8116 4616
rect 7699 4576 8116 4604
rect 7699 4573 7711 4576
rect 7653 4567 7711 4573
rect 1670 4496 1676 4548
rect 1728 4496 1734 4548
rect 3142 4536 3148 4548
rect 2898 4508 3148 4536
rect 3142 4496 3148 4508
rect 3200 4496 3206 4548
rect 4341 4539 4399 4545
rect 4341 4505 4353 4539
rect 4387 4536 4399 4539
rect 6086 4536 6092 4548
rect 4387 4508 6092 4536
rect 4387 4505 4399 4508
rect 4341 4499 4399 4505
rect 6086 4496 6092 4508
rect 6144 4536 6150 4548
rect 7484 4536 7512 4567
rect 6144 4508 7512 4536
rect 6144 4496 6150 4508
rect 7558 4496 7564 4548
rect 7616 4536 7622 4548
rect 7668 4536 7696 4567
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 8478 4564 8484 4616
rect 8536 4564 8542 4616
rect 8570 4564 8576 4616
rect 8628 4564 8634 4616
rect 7616 4508 7696 4536
rect 8021 4539 8079 4545
rect 7616 4496 7622 4508
rect 8021 4505 8033 4539
rect 8067 4505 8079 4539
rect 8021 4499 8079 4505
rect 7006 4428 7012 4480
rect 7064 4468 7070 4480
rect 7193 4471 7251 4477
rect 7193 4468 7205 4471
rect 7064 4440 7205 4468
rect 7064 4428 7070 4440
rect 7193 4437 7205 4440
rect 7239 4437 7251 4471
rect 7193 4431 7251 4437
rect 7466 4428 7472 4480
rect 7524 4468 7530 4480
rect 8036 4468 8064 4499
rect 7524 4440 8064 4468
rect 7524 4428 7530 4440
rect 1104 4378 11316 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 11316 4378
rect 1104 4304 11316 4326
rect 1670 4224 1676 4276
rect 1728 4264 1734 4276
rect 2133 4267 2191 4273
rect 2133 4264 2145 4267
rect 1728 4236 2145 4264
rect 1728 4224 1734 4236
rect 2133 4233 2145 4236
rect 2179 4233 2191 4267
rect 2133 4227 2191 4233
rect 2501 4267 2559 4273
rect 2501 4233 2513 4267
rect 2547 4264 2559 4267
rect 2866 4264 2872 4276
rect 2547 4236 2872 4264
rect 2547 4233 2559 4236
rect 2501 4227 2559 4233
rect 2866 4224 2872 4236
rect 2924 4224 2930 4276
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 3108 4236 4568 4264
rect 3108 4224 3114 4236
rect 1578 4156 1584 4208
rect 1636 4196 1642 4208
rect 3447 4199 3505 4205
rect 3447 4196 3459 4199
rect 1636 4168 3459 4196
rect 1636 4156 1642 4168
rect 3447 4165 3459 4168
rect 3493 4165 3505 4199
rect 3447 4159 3505 4165
rect 4062 4156 4068 4208
rect 4120 4196 4126 4208
rect 4433 4199 4491 4205
rect 4433 4196 4445 4199
rect 4120 4168 4445 4196
rect 4120 4156 4126 4168
rect 4433 4165 4445 4168
rect 4479 4165 4491 4199
rect 4433 4159 4491 4165
rect 1210 4088 1216 4140
rect 1268 4128 1274 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 1268 4100 1409 4128
rect 1268 4088 1274 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 2961 4131 3019 4137
rect 2961 4128 2973 4131
rect 2639 4100 2973 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 2961 4097 2973 4100
rect 3007 4097 3019 4131
rect 2961 4091 3019 4097
rect 1302 4020 1308 4072
rect 1360 4060 1366 4072
rect 1688 4060 1716 4091
rect 3050 4088 3056 4140
rect 3108 4128 3114 4140
rect 3145 4131 3203 4137
rect 3145 4128 3157 4131
rect 3108 4100 3157 4128
rect 3108 4088 3114 4100
rect 3145 4097 3157 4100
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 3234 4088 3240 4140
rect 3292 4088 3298 4140
rect 3326 4088 3332 4140
rect 3384 4088 3390 4140
rect 4540 4137 4568 4236
rect 4798 4224 4804 4276
rect 4856 4264 4862 4276
rect 5077 4267 5135 4273
rect 5077 4264 5089 4267
rect 4856 4236 5089 4264
rect 4856 4224 4862 4236
rect 5077 4233 5089 4236
rect 5123 4233 5135 4267
rect 5077 4227 5135 4233
rect 5537 4267 5595 4273
rect 5537 4233 5549 4267
rect 5583 4264 5595 4267
rect 6362 4264 6368 4276
rect 5583 4236 6368 4264
rect 5583 4233 5595 4236
rect 5537 4227 5595 4233
rect 6362 4224 6368 4236
rect 6420 4224 6426 4276
rect 6730 4224 6736 4276
rect 6788 4264 6794 4276
rect 8481 4267 8539 4273
rect 6788 4236 8340 4264
rect 6788 4224 6794 4236
rect 5445 4199 5503 4205
rect 5445 4165 5457 4199
rect 5491 4196 5503 4199
rect 6178 4196 6184 4208
rect 5491 4168 6184 4196
rect 5491 4165 5503 4168
rect 5445 4159 5503 4165
rect 6178 4156 6184 4168
rect 6236 4156 6242 4208
rect 6748 4137 6776 4224
rect 7006 4156 7012 4208
rect 7064 4156 7070 4208
rect 7650 4156 7656 4208
rect 7708 4156 7714 4208
rect 8312 4196 8340 4236
rect 8481 4233 8493 4267
rect 8527 4264 8539 4267
rect 8570 4264 8576 4276
rect 8527 4236 8576 4264
rect 8527 4233 8539 4236
rect 8481 4227 8539 4233
rect 8570 4224 8576 4236
rect 8628 4224 8634 4276
rect 9214 4196 9220 4208
rect 8312 4168 9220 4196
rect 9214 4156 9220 4168
rect 9272 4156 9278 4208
rect 4203 4131 4261 4137
rect 4203 4128 4215 4131
rect 3436 4100 4215 4128
rect 1949 4063 2007 4069
rect 1949 4060 1961 4063
rect 1360 4032 1961 4060
rect 1360 4020 1366 4032
rect 1949 4029 1961 4032
rect 1995 4029 2007 4063
rect 1949 4023 2007 4029
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4060 2743 4063
rect 2866 4060 2872 4072
rect 2731 4032 2872 4060
rect 2731 4029 2743 4032
rect 2685 4023 2743 4029
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 3436 3992 3464 4100
rect 4203 4097 4215 4100
rect 4249 4097 4261 4131
rect 4203 4091 4261 4097
rect 4341 4131 4399 4137
rect 4341 4097 4353 4131
rect 4387 4097 4399 4131
rect 4341 4091 4399 4097
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 6733 4131 6791 4137
rect 6733 4097 6745 4131
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 3605 4063 3663 4069
rect 3605 4029 3617 4063
rect 3651 4060 3663 4063
rect 3878 4060 3884 4072
rect 3651 4032 3884 4060
rect 3651 4029 3663 4032
rect 3605 4023 3663 4029
rect 3878 4020 3884 4032
rect 3936 4060 3942 4072
rect 4065 4063 4123 4069
rect 4065 4060 4077 4063
rect 3936 4032 4077 4060
rect 3936 4020 3942 4032
rect 4065 4029 4077 4032
rect 4111 4029 4123 4063
rect 4356 4060 4384 4091
rect 4798 4060 4804 4072
rect 4356 4032 4804 4060
rect 4065 4023 4123 4029
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 5258 4020 5264 4072
rect 5316 4060 5322 4072
rect 5629 4063 5687 4069
rect 5629 4060 5641 4063
rect 5316 4032 5641 4060
rect 5316 4020 5322 4032
rect 5629 4029 5641 4032
rect 5675 4029 5687 4063
rect 7558 4060 7564 4072
rect 5629 4023 5687 4029
rect 6840 4032 7564 4060
rect 6840 3992 6868 4032
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 1627 3964 3464 3992
rect 4632 3964 6868 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 1854 3884 1860 3936
rect 1912 3884 1918 3936
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 4632 3924 4660 3964
rect 2832 3896 4660 3924
rect 4709 3927 4767 3933
rect 2832 3884 2838 3896
rect 4709 3893 4721 3927
rect 4755 3924 4767 3927
rect 5258 3924 5264 3936
rect 4755 3896 5264 3924
rect 4755 3893 4767 3896
rect 4709 3887 4767 3893
rect 5258 3884 5264 3896
rect 5316 3884 5322 3936
rect 1104 3834 11316 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 11316 3834
rect 1104 3760 11316 3782
rect 1210 3680 1216 3732
rect 1268 3720 1274 3732
rect 1673 3723 1731 3729
rect 1673 3720 1685 3723
rect 1268 3692 1685 3720
rect 1268 3680 1274 3692
rect 1673 3689 1685 3692
rect 1719 3689 1731 3723
rect 1673 3683 1731 3689
rect 2038 3680 2044 3732
rect 2096 3720 2102 3732
rect 3881 3723 3939 3729
rect 2096 3692 2912 3720
rect 2096 3680 2102 3692
rect 1581 3655 1639 3661
rect 1581 3621 1593 3655
rect 1627 3652 1639 3655
rect 2774 3652 2780 3664
rect 1627 3624 2544 3652
rect 1627 3621 1639 3624
rect 1581 3615 1639 3621
rect 1854 3544 1860 3596
rect 1912 3584 1918 3596
rect 1912 3556 2452 3584
rect 1912 3544 1918 3556
rect 1118 3476 1124 3528
rect 1176 3516 1182 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 1176 3488 1409 3516
rect 1176 3476 1182 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 2038 3476 2044 3528
rect 2096 3476 2102 3528
rect 2424 3525 2452 3556
rect 2516 3525 2544 3624
rect 2700 3624 2780 3652
rect 2700 3525 2728 3624
rect 2774 3612 2780 3624
rect 2832 3612 2838 3664
rect 2884 3525 2912 3692
rect 3881 3689 3893 3723
rect 3927 3720 3939 3723
rect 3970 3720 3976 3732
rect 3927 3692 3976 3720
rect 3927 3689 3939 3692
rect 3881 3683 3939 3689
rect 3970 3680 3976 3692
rect 4028 3680 4034 3732
rect 3142 3612 3148 3664
rect 3200 3652 3206 3664
rect 4157 3655 4215 3661
rect 4157 3652 4169 3655
rect 3200 3624 4169 3652
rect 3200 3612 3206 3624
rect 4157 3621 4169 3624
rect 4203 3652 4215 3655
rect 5718 3652 5724 3664
rect 4203 3624 5724 3652
rect 4203 3621 4215 3624
rect 4157 3615 4215 3621
rect 5718 3612 5724 3624
rect 5776 3612 5782 3664
rect 5258 3544 5264 3596
rect 5316 3544 5322 3596
rect 5350 3544 5356 3596
rect 5408 3544 5414 3596
rect 2409 3519 2467 3525
rect 2409 3485 2421 3519
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 2501 3519 2559 3525
rect 2501 3485 2513 3519
rect 2547 3485 2559 3519
rect 2501 3479 2559 3485
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3485 2743 3519
rect 2685 3479 2743 3485
rect 2869 3519 2927 3525
rect 2869 3485 2881 3519
rect 2915 3485 2927 3519
rect 4798 3516 4804 3528
rect 2869 3479 2927 3485
rect 3160 3488 4804 3516
rect 2133 3451 2191 3457
rect 2133 3417 2145 3451
rect 2179 3417 2191 3451
rect 2133 3411 2191 3417
rect 2225 3451 2283 3457
rect 2225 3417 2237 3451
rect 2271 3448 2283 3451
rect 2700 3448 2728 3479
rect 2271 3420 2728 3448
rect 2777 3451 2835 3457
rect 2271 3417 2283 3420
rect 2225 3411 2283 3417
rect 2777 3417 2789 3451
rect 2823 3448 2835 3451
rect 3160 3448 3188 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3516 5227 3519
rect 6270 3516 6276 3528
rect 5215 3488 6276 3516
rect 5215 3485 5227 3488
rect 5169 3479 5227 3485
rect 6270 3476 6276 3488
rect 6328 3476 6334 3528
rect 2823 3420 3188 3448
rect 2823 3417 2835 3420
rect 2777 3411 2835 3417
rect 1762 3340 1768 3392
rect 1820 3380 1826 3392
rect 1857 3383 1915 3389
rect 1857 3380 1869 3383
rect 1820 3352 1869 3380
rect 1820 3340 1826 3352
rect 1857 3349 1869 3352
rect 1903 3349 1915 3383
rect 2148 3380 2176 3411
rect 3234 3408 3240 3460
rect 3292 3408 3298 3460
rect 3973 3451 4031 3457
rect 3973 3417 3985 3451
rect 4019 3417 4031 3451
rect 3973 3411 4031 3417
rect 2682 3380 2688 3392
rect 2148 3352 2688 3380
rect 1857 3343 1915 3349
rect 2682 3340 2688 3352
rect 2740 3340 2746 3392
rect 2866 3340 2872 3392
rect 2924 3380 2930 3392
rect 3053 3383 3111 3389
rect 3053 3380 3065 3383
rect 2924 3352 3065 3380
rect 2924 3340 2930 3352
rect 3053 3349 3065 3352
rect 3099 3349 3111 3383
rect 3053 3343 3111 3349
rect 3329 3383 3387 3389
rect 3329 3349 3341 3383
rect 3375 3380 3387 3383
rect 3988 3380 4016 3411
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 4341 3451 4399 3457
rect 4341 3448 4353 3451
rect 4120 3420 4353 3448
rect 4120 3408 4126 3420
rect 4341 3417 4353 3420
rect 4387 3417 4399 3451
rect 7466 3448 7472 3460
rect 4341 3411 4399 3417
rect 4632 3420 7472 3448
rect 4632 3380 4660 3420
rect 7466 3408 7472 3420
rect 7524 3408 7530 3460
rect 3375 3352 4660 3380
rect 3375 3349 3387 3352
rect 3329 3343 3387 3349
rect 4706 3340 4712 3392
rect 4764 3380 4770 3392
rect 4801 3383 4859 3389
rect 4801 3380 4813 3383
rect 4764 3352 4813 3380
rect 4764 3340 4770 3352
rect 4801 3349 4813 3352
rect 4847 3349 4859 3383
rect 4801 3343 4859 3349
rect 1104 3290 11316 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 11316 3290
rect 1104 3216 11316 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3176 1639 3179
rect 3234 3176 3240 3188
rect 1627 3148 3240 3176
rect 1627 3145 1639 3148
rect 1581 3139 1639 3145
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 4341 3179 4399 3185
rect 4341 3145 4353 3179
rect 4387 3176 4399 3179
rect 4798 3176 4804 3188
rect 4387 3148 4804 3176
rect 4387 3145 4399 3148
rect 4341 3139 4399 3145
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 6181 3179 6239 3185
rect 6181 3145 6193 3179
rect 6227 3176 6239 3179
rect 6270 3176 6276 3188
rect 6227 3148 6276 3176
rect 6227 3145 6239 3148
rect 6181 3139 6239 3145
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 9674 3136 9680 3188
rect 9732 3136 9738 3188
rect 1118 3068 1124 3120
rect 1176 3108 1182 3120
rect 1673 3111 1731 3117
rect 1673 3108 1685 3111
rect 1176 3080 1685 3108
rect 1176 3068 1182 3080
rect 1673 3077 1685 3080
rect 1719 3077 1731 3111
rect 1673 3071 1731 3077
rect 2866 3068 2872 3120
rect 2924 3068 2930 3120
rect 3142 3068 3148 3120
rect 3200 3108 3206 3120
rect 3200 3080 3358 3108
rect 3200 3068 3206 3080
rect 4706 3068 4712 3120
rect 4764 3068 4770 3120
rect 5718 3068 5724 3120
rect 5776 3068 5782 3120
rect 9398 3068 9404 3120
rect 9456 3108 9462 3120
rect 9493 3111 9551 3117
rect 9493 3108 9505 3111
rect 9456 3080 9505 3108
rect 9456 3068 9462 3080
rect 9493 3077 9505 3080
rect 9539 3077 9551 3111
rect 9692 3108 9720 3136
rect 9692 3080 9982 3108
rect 9493 3071 9551 3077
rect 1302 3000 1308 3052
rect 1360 3040 1366 3052
rect 1397 3043 1455 3049
rect 1397 3040 1409 3043
rect 1360 3012 1409 3040
rect 1360 3000 1366 3012
rect 1397 3009 1409 3012
rect 1443 3040 1455 3043
rect 1857 3043 1915 3049
rect 1857 3040 1869 3043
rect 1443 3012 1869 3040
rect 1443 3009 1455 3012
rect 1397 3003 1455 3009
rect 1857 3009 1869 3012
rect 1903 3009 1915 3043
rect 1857 3003 1915 3009
rect 9214 3000 9220 3052
rect 9272 3000 9278 3052
rect 2406 2932 2412 2984
rect 2464 2972 2470 2984
rect 2593 2975 2651 2981
rect 2593 2972 2605 2975
rect 2464 2944 2605 2972
rect 2464 2932 2470 2944
rect 2593 2941 2605 2944
rect 2639 2972 2651 2975
rect 4433 2975 4491 2981
rect 4433 2972 4445 2975
rect 2639 2944 4445 2972
rect 2639 2941 2651 2944
rect 2593 2935 2651 2941
rect 4433 2941 4445 2944
rect 4479 2941 4491 2975
rect 4433 2935 4491 2941
rect 3234 2796 3240 2848
rect 3292 2836 3298 2848
rect 3510 2836 3516 2848
rect 3292 2808 3516 2836
rect 3292 2796 3298 2808
rect 3510 2796 3516 2808
rect 3568 2796 3574 2848
rect 10962 2796 10968 2848
rect 11020 2796 11026 2848
rect 1104 2746 11316 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 11316 2746
rect 1104 2672 11316 2694
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 3145 2635 3203 2641
rect 3145 2632 3157 2635
rect 2832 2604 3157 2632
rect 2832 2592 2838 2604
rect 3145 2601 3157 2604
rect 3191 2632 3203 2635
rect 3326 2632 3332 2644
rect 3191 2604 3332 2632
rect 3191 2601 3203 2604
rect 3145 2595 3203 2601
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 1394 2456 1400 2508
rect 1452 2496 1458 2508
rect 2406 2496 2412 2508
rect 1452 2468 2412 2496
rect 1452 2456 1458 2468
rect 2406 2456 2412 2468
rect 2464 2456 2470 2508
rect 10962 2388 10968 2440
rect 11020 2388 11026 2440
rect 1673 2363 1731 2369
rect 1673 2329 1685 2363
rect 1719 2360 1731 2363
rect 1762 2360 1768 2372
rect 1719 2332 1768 2360
rect 1719 2329 1731 2332
rect 1673 2323 1731 2329
rect 1762 2320 1768 2332
rect 1820 2320 1826 2372
rect 3510 2360 3516 2372
rect 2898 2332 3516 2360
rect 3510 2320 3516 2332
rect 3568 2320 3574 2372
rect 10686 2320 10692 2372
rect 10744 2320 10750 2372
rect 1104 2202 11316 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 11316 2202
rect 1104 2128 11316 2150
<< via1 >>
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 4804 11840 4856 11892
rect 1308 11772 1360 11824
rect 1124 11704 1176 11756
rect 1860 11747 1912 11756
rect 1860 11713 1869 11747
rect 1869 11713 1903 11747
rect 1903 11713 1912 11747
rect 1860 11704 1912 11713
rect 2412 11704 2464 11756
rect 2504 11747 2556 11756
rect 2504 11713 2513 11747
rect 2513 11713 2547 11747
rect 2547 11713 2556 11747
rect 2504 11704 2556 11713
rect 10692 11815 10744 11824
rect 10692 11781 10701 11815
rect 10701 11781 10735 11815
rect 10735 11781 10744 11815
rect 10692 11772 10744 11781
rect 1216 11636 1268 11688
rect 10968 11747 11020 11756
rect 10968 11713 10977 11747
rect 10977 11713 11011 11747
rect 11011 11713 11020 11747
rect 10968 11704 11020 11713
rect 5724 11568 5776 11620
rect 2412 11543 2464 11552
rect 2412 11509 2421 11543
rect 2421 11509 2455 11543
rect 2455 11509 2464 11543
rect 2412 11500 2464 11509
rect 3056 11500 3108 11552
rect 3148 11543 3200 11552
rect 3148 11509 3157 11543
rect 3157 11509 3191 11543
rect 3191 11509 3200 11543
rect 3148 11500 3200 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 2780 11296 2832 11348
rect 3332 11160 3384 11212
rect 5448 11160 5500 11212
rect 10968 11339 11020 11348
rect 10968 11305 10977 11339
rect 10977 11305 11011 11339
rect 11011 11305 11020 11339
rect 10968 11296 11020 11305
rect 6460 11271 6512 11280
rect 6460 11237 6469 11271
rect 6469 11237 6503 11271
rect 6503 11237 6512 11271
rect 6460 11228 6512 11237
rect 3240 11135 3292 11144
rect 3240 11101 3249 11135
rect 3249 11101 3283 11135
rect 3283 11101 3292 11135
rect 3240 11092 3292 11101
rect 7472 11160 7524 11212
rect 2780 11024 2832 11076
rect 6644 11135 6696 11144
rect 6644 11101 6653 11135
rect 6653 11101 6687 11135
rect 6687 11101 6696 11135
rect 6644 11092 6696 11101
rect 8760 11092 8812 11144
rect 4804 11024 4856 11076
rect 1860 10956 1912 11008
rect 7748 11024 7800 11076
rect 8668 11024 8720 11076
rect 9496 11067 9548 11076
rect 9496 11033 9505 11067
rect 9505 11033 9539 11067
rect 9539 11033 9548 11067
rect 9496 11024 9548 11033
rect 9956 11024 10008 11076
rect 5264 10956 5316 11008
rect 6368 10999 6420 11008
rect 6368 10965 6377 10999
rect 6377 10965 6411 10999
rect 6411 10965 6420 10999
rect 6368 10956 6420 10965
rect 8116 10956 8168 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 3608 10727 3660 10736
rect 3608 10693 3617 10727
rect 3617 10693 3651 10727
rect 3651 10693 3660 10727
rect 3608 10684 3660 10693
rect 3884 10684 3936 10736
rect 4896 10684 4948 10736
rect 5264 10752 5316 10804
rect 5816 10752 5868 10804
rect 6368 10752 6420 10804
rect 9496 10752 9548 10804
rect 6644 10684 6696 10736
rect 8024 10684 8076 10736
rect 1308 10616 1360 10668
rect 1860 10659 1912 10668
rect 1860 10625 1869 10659
rect 1869 10625 1903 10659
rect 1903 10625 1912 10659
rect 1860 10616 1912 10625
rect 2688 10591 2740 10600
rect 2688 10557 2697 10591
rect 2697 10557 2731 10591
rect 2731 10557 2740 10591
rect 2688 10548 2740 10557
rect 3332 10659 3384 10668
rect 3332 10625 3341 10659
rect 3341 10625 3375 10659
rect 3375 10625 3384 10659
rect 3332 10616 3384 10625
rect 2964 10523 3016 10532
rect 2964 10489 2973 10523
rect 2973 10489 3007 10523
rect 3007 10489 3016 10523
rect 2964 10480 3016 10489
rect 1860 10412 1912 10464
rect 2044 10455 2096 10464
rect 2044 10421 2053 10455
rect 2053 10421 2087 10455
rect 2087 10421 2096 10455
rect 2044 10412 2096 10421
rect 2504 10412 2556 10464
rect 4068 10412 4120 10464
rect 4896 10412 4948 10464
rect 5264 10548 5316 10600
rect 9220 10659 9272 10668
rect 9220 10625 9229 10659
rect 9229 10625 9263 10659
rect 9263 10625 9272 10659
rect 9220 10616 9272 10625
rect 9312 10616 9364 10668
rect 5540 10480 5592 10532
rect 7288 10548 7340 10600
rect 7932 10548 7984 10600
rect 8576 10548 8628 10600
rect 6276 10412 6328 10464
rect 6736 10412 6788 10464
rect 8392 10412 8444 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 2504 10251 2556 10260
rect 2504 10217 2513 10251
rect 2513 10217 2547 10251
rect 2547 10217 2556 10251
rect 2504 10208 2556 10217
rect 3608 10208 3660 10260
rect 5264 10251 5316 10260
rect 5264 10217 5273 10251
rect 5273 10217 5307 10251
rect 5307 10217 5316 10251
rect 5264 10208 5316 10217
rect 7288 10251 7340 10260
rect 7288 10217 7297 10251
rect 7297 10217 7331 10251
rect 7331 10217 7340 10251
rect 7288 10208 7340 10217
rect 1124 10072 1176 10124
rect 1216 10004 1268 10056
rect 4436 10115 4488 10124
rect 4436 10081 4445 10115
rect 4445 10081 4479 10115
rect 4479 10081 4488 10115
rect 4436 10072 4488 10081
rect 1860 10004 1912 10056
rect 2688 9979 2740 9988
rect 2688 9945 2697 9979
rect 2697 9945 2731 9979
rect 2731 9945 2740 9979
rect 2688 9936 2740 9945
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 2964 9936 3016 9988
rect 4620 10047 4672 10056
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 4620 10004 4672 10013
rect 4896 10047 4948 10056
rect 4896 10013 4905 10047
rect 4905 10013 4939 10047
rect 4939 10013 4948 10047
rect 4896 10004 4948 10013
rect 5264 10004 5316 10056
rect 4160 9868 4212 9920
rect 4252 9911 4304 9920
rect 4252 9877 4261 9911
rect 4261 9877 4295 9911
rect 4295 9877 4304 9911
rect 4252 9868 4304 9877
rect 4528 9868 4580 9920
rect 5448 9979 5500 9988
rect 5448 9945 5457 9979
rect 5457 9945 5491 9979
rect 5491 9945 5500 9979
rect 5448 9936 5500 9945
rect 6644 10140 6696 10192
rect 7748 10140 7800 10192
rect 6276 10072 6328 10124
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 9036 10004 9088 10056
rect 5540 9868 5592 9920
rect 6644 9868 6696 9920
rect 6736 9911 6788 9920
rect 6736 9877 6745 9911
rect 6745 9877 6779 9911
rect 6779 9877 6788 9911
rect 6736 9868 6788 9877
rect 7748 9911 7800 9920
rect 7748 9877 7757 9911
rect 7757 9877 7791 9911
rect 7791 9877 7800 9911
rect 7748 9868 7800 9877
rect 7840 9868 7892 9920
rect 8116 9868 8168 9920
rect 9404 9868 9456 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 1584 9664 1636 9716
rect 1308 9528 1360 9580
rect 2780 9596 2832 9648
rect 3516 9596 3568 9648
rect 4252 9596 4304 9648
rect 5724 9639 5776 9648
rect 5724 9605 5741 9639
rect 5741 9605 5776 9639
rect 5724 9596 5776 9605
rect 5816 9639 5868 9648
rect 5816 9605 5825 9639
rect 5825 9605 5859 9639
rect 5859 9605 5868 9639
rect 5816 9596 5868 9605
rect 5908 9639 5960 9648
rect 5908 9605 5916 9639
rect 5916 9605 5950 9639
rect 5950 9605 5960 9639
rect 5908 9596 5960 9605
rect 6644 9664 6696 9716
rect 6736 9664 6788 9716
rect 7748 9664 7800 9716
rect 3792 9528 3844 9580
rect 4068 9571 4120 9580
rect 4068 9537 4077 9571
rect 4077 9537 4111 9571
rect 4111 9537 4120 9571
rect 4068 9528 4120 9537
rect 4160 9528 4212 9580
rect 4896 9571 4948 9580
rect 4896 9537 4905 9571
rect 4905 9537 4939 9571
rect 4939 9537 4948 9571
rect 4896 9528 4948 9537
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 6644 9571 6696 9580
rect 6644 9537 6653 9571
rect 6653 9537 6687 9571
rect 6687 9537 6696 9571
rect 6644 9528 6696 9537
rect 8760 9596 8812 9648
rect 6920 9528 6972 9580
rect 7932 9528 7984 9580
rect 3148 9392 3200 9444
rect 3424 9392 3476 9444
rect 3516 9392 3568 9444
rect 5264 9460 5316 9512
rect 5632 9460 5684 9512
rect 5724 9460 5776 9512
rect 6184 9460 6236 9512
rect 6460 9460 6512 9512
rect 9312 9460 9364 9512
rect 3792 9367 3844 9376
rect 3792 9333 3801 9367
rect 3801 9333 3835 9367
rect 3835 9333 3844 9367
rect 3792 9324 3844 9333
rect 5908 9392 5960 9444
rect 8300 9392 8352 9444
rect 9220 9392 9272 9444
rect 4528 9324 4580 9376
rect 4620 9324 4672 9376
rect 5632 9324 5684 9376
rect 8116 9324 8168 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 5264 9120 5316 9172
rect 6920 9120 6972 9172
rect 3792 9052 3844 9104
rect 1676 9027 1728 9036
rect 1676 8993 1685 9027
rect 1685 8993 1719 9027
rect 1719 8993 1728 9027
rect 1676 8984 1728 8993
rect 4068 8984 4120 9036
rect 4896 9052 4948 9104
rect 5724 8984 5776 9036
rect 7472 8984 7524 9036
rect 1032 8916 1084 8968
rect 5356 8916 5408 8968
rect 6000 8916 6052 8968
rect 8760 8959 8812 8968
rect 8760 8925 8769 8959
rect 8769 8925 8803 8959
rect 8803 8925 8812 8959
rect 8760 8916 8812 8925
rect 1952 8891 2004 8900
rect 1952 8857 1961 8891
rect 1961 8857 1995 8891
rect 1995 8857 2004 8891
rect 1952 8848 2004 8857
rect 3884 8848 3936 8900
rect 8024 8848 8076 8900
rect 3332 8780 3384 8832
rect 3424 8823 3476 8832
rect 3424 8789 3433 8823
rect 3433 8789 3467 8823
rect 3467 8789 3476 8823
rect 3424 8780 3476 8789
rect 8208 8848 8260 8900
rect 9956 8916 10008 8968
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 1032 8508 1084 8560
rect 1952 8576 2004 8628
rect 3424 8576 3476 8628
rect 5540 8576 5592 8628
rect 6644 8576 6696 8628
rect 8300 8619 8352 8628
rect 8300 8585 8309 8619
rect 8309 8585 8343 8619
rect 8343 8585 8352 8619
rect 8300 8576 8352 8585
rect 2964 8508 3016 8560
rect 1308 8440 1360 8492
rect 3332 8440 3384 8492
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 5724 8440 5776 8492
rect 6736 8508 6788 8560
rect 7656 8508 7708 8560
rect 7932 8440 7984 8492
rect 9312 8508 9364 8560
rect 8668 8440 8720 8492
rect 2872 8415 2924 8424
rect 2872 8381 2881 8415
rect 2881 8381 2915 8415
rect 2915 8381 2924 8415
rect 2872 8372 2924 8381
rect 2596 8236 2648 8288
rect 3148 8372 3200 8424
rect 5632 8372 5684 8424
rect 6184 8372 6236 8424
rect 6736 8372 6788 8424
rect 7840 8304 7892 8356
rect 8208 8304 8260 8356
rect 4712 8236 4764 8288
rect 5264 8236 5316 8288
rect 6368 8236 6420 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 2872 8032 2924 8084
rect 6736 8032 6788 8084
rect 2780 7964 2832 8016
rect 1308 7828 1360 7880
rect 2688 7871 2740 7880
rect 2688 7837 2697 7871
rect 2697 7837 2731 7871
rect 2731 7837 2740 7871
rect 2688 7828 2740 7837
rect 4068 7939 4120 7948
rect 4068 7905 4077 7939
rect 4077 7905 4111 7939
rect 4111 7905 4120 7939
rect 6644 7964 6696 8016
rect 4068 7896 4120 7905
rect 6276 7939 6328 7948
rect 6276 7905 6285 7939
rect 6285 7905 6319 7939
rect 6319 7905 6328 7939
rect 6276 7896 6328 7905
rect 6368 7939 6420 7948
rect 6368 7905 6377 7939
rect 6377 7905 6411 7939
rect 6411 7905 6420 7939
rect 6368 7896 6420 7905
rect 3148 7871 3200 7880
rect 3148 7837 3157 7871
rect 3157 7837 3191 7871
rect 3191 7837 3200 7871
rect 3148 7828 3200 7837
rect 6552 7828 6604 7880
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 2780 7692 2832 7744
rect 2964 7803 3016 7812
rect 2964 7769 2999 7803
rect 2999 7769 3016 7803
rect 2964 7760 3016 7769
rect 4344 7803 4396 7812
rect 4344 7769 4353 7803
rect 4353 7769 4387 7803
rect 4387 7769 4396 7803
rect 4344 7760 4396 7769
rect 3884 7692 3936 7744
rect 5356 7692 5408 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 1584 7488 1636 7540
rect 1676 7420 1728 7472
rect 3884 7420 3936 7472
rect 4344 7488 4396 7540
rect 5356 7488 5408 7540
rect 8116 7420 8168 7472
rect 9956 7420 10008 7472
rect 1676 7327 1728 7336
rect 1676 7293 1685 7327
rect 1685 7293 1719 7327
rect 1719 7293 1728 7327
rect 1676 7284 1728 7293
rect 3516 7395 3568 7404
rect 3516 7361 3525 7395
rect 3525 7361 3559 7395
rect 3559 7361 3568 7395
rect 3516 7352 3568 7361
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 3700 7395 3752 7404
rect 3700 7361 3735 7395
rect 3735 7361 3752 7395
rect 3700 7352 3752 7361
rect 3884 7327 3936 7336
rect 3884 7293 3893 7327
rect 3893 7293 3927 7327
rect 3927 7293 3936 7327
rect 3884 7284 3936 7293
rect 5264 7327 5316 7336
rect 5264 7293 5273 7327
rect 5273 7293 5307 7327
rect 5307 7293 5316 7327
rect 5264 7284 5316 7293
rect 2964 7216 3016 7268
rect 3424 7216 3476 7268
rect 2780 7148 2832 7200
rect 3056 7148 3108 7200
rect 3516 7148 3568 7200
rect 4068 7148 4120 7200
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 8760 7352 8812 7404
rect 10968 7191 11020 7200
rect 10968 7157 10977 7191
rect 10977 7157 11011 7191
rect 11011 7157 11020 7191
rect 10968 7148 11020 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 1676 6944 1728 6996
rect 3424 6944 3476 6996
rect 3700 6876 3752 6928
rect 6644 6851 6696 6860
rect 6644 6817 6653 6851
rect 6653 6817 6687 6851
rect 6687 6817 6696 6851
rect 6644 6808 6696 6817
rect 10784 6851 10836 6860
rect 10784 6817 10793 6851
rect 10793 6817 10827 6851
rect 10827 6817 10836 6851
rect 10784 6808 10836 6817
rect 1216 6740 1268 6792
rect 1308 6672 1360 6724
rect 2688 6740 2740 6792
rect 2872 6740 2924 6792
rect 5724 6740 5776 6792
rect 10968 6783 11020 6792
rect 10968 6749 10977 6783
rect 10977 6749 11011 6783
rect 11011 6749 11020 6783
rect 10968 6740 11020 6749
rect 3056 6672 3108 6724
rect 1860 6647 1912 6656
rect 1860 6613 1869 6647
rect 1869 6613 1903 6647
rect 1903 6613 1912 6647
rect 1860 6604 1912 6613
rect 2964 6604 3016 6656
rect 4620 6647 4672 6656
rect 4620 6613 4629 6647
rect 4629 6613 4663 6647
rect 4663 6613 4672 6647
rect 6920 6715 6972 6724
rect 6920 6681 6929 6715
rect 6929 6681 6963 6715
rect 6963 6681 6972 6715
rect 6920 6672 6972 6681
rect 7656 6672 7708 6724
rect 4620 6604 4672 6613
rect 5448 6604 5500 6656
rect 7932 6604 7984 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 1216 6400 1268 6452
rect 2780 6400 2832 6452
rect 3884 6400 3936 6452
rect 3148 6332 3200 6384
rect 3976 6332 4028 6384
rect 1216 6264 1268 6316
rect 6000 6264 6052 6316
rect 6460 6264 6512 6316
rect 6920 6400 6972 6452
rect 8024 6400 8076 6452
rect 1400 6128 1452 6180
rect 2412 6239 2464 6248
rect 2412 6205 2421 6239
rect 2421 6205 2455 6239
rect 2455 6205 2464 6239
rect 2412 6196 2464 6205
rect 2964 6060 3016 6112
rect 3608 6060 3660 6112
rect 4804 6196 4856 6248
rect 4712 6060 4764 6112
rect 5908 6060 5960 6112
rect 7748 6264 7800 6316
rect 7840 6307 7892 6316
rect 7840 6273 7849 6307
rect 7849 6273 7883 6307
rect 7883 6273 7892 6307
rect 7840 6264 7892 6273
rect 7932 6264 7984 6316
rect 8300 6196 8352 6248
rect 8852 6264 8904 6316
rect 8576 6239 8628 6248
rect 8576 6205 8585 6239
rect 8585 6205 8619 6239
rect 8619 6205 8628 6239
rect 8576 6196 8628 6205
rect 10968 6332 11020 6384
rect 7748 6171 7800 6180
rect 7748 6137 7757 6171
rect 7757 6137 7791 6171
rect 7791 6137 7800 6171
rect 7748 6128 7800 6137
rect 8116 6060 8168 6112
rect 8392 6060 8444 6112
rect 8668 6060 8720 6112
rect 9312 6103 9364 6112
rect 9312 6069 9321 6103
rect 9321 6069 9355 6103
rect 9355 6069 9364 6103
rect 9312 6060 9364 6069
rect 9496 6103 9548 6112
rect 9496 6069 9505 6103
rect 9505 6069 9539 6103
rect 9539 6069 9548 6103
rect 9496 6060 9548 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 2412 5856 2464 5908
rect 4804 5856 4856 5908
rect 6644 5788 6696 5840
rect 2872 5720 2924 5772
rect 3240 5763 3292 5772
rect 3240 5729 3249 5763
rect 3249 5729 3283 5763
rect 3283 5729 3292 5763
rect 3240 5720 3292 5729
rect 5264 5720 5316 5772
rect 5724 5720 5776 5772
rect 1308 5652 1360 5704
rect 2964 5695 3016 5704
rect 2964 5661 2973 5695
rect 2973 5661 3007 5695
rect 3007 5661 3016 5695
rect 2964 5652 3016 5661
rect 5908 5652 5960 5704
rect 6460 5763 6512 5772
rect 6460 5729 6469 5763
rect 6469 5729 6503 5763
rect 6503 5729 6512 5763
rect 6460 5720 6512 5729
rect 8852 5856 8904 5908
rect 9036 5856 9088 5908
rect 9312 5856 9364 5908
rect 8300 5788 8352 5840
rect 8484 5788 8536 5840
rect 8024 5763 8076 5772
rect 8024 5729 8033 5763
rect 8033 5729 8067 5763
rect 8067 5729 8076 5763
rect 8024 5720 8076 5729
rect 8668 5788 8720 5840
rect 1860 5584 1912 5636
rect 3056 5559 3108 5568
rect 3056 5525 3065 5559
rect 3065 5525 3099 5559
rect 3099 5525 3108 5559
rect 3056 5516 3108 5525
rect 6092 5627 6144 5636
rect 6092 5593 6101 5627
rect 6101 5593 6135 5627
rect 6135 5593 6144 5627
rect 6092 5584 6144 5593
rect 6184 5627 6236 5636
rect 6184 5593 6193 5627
rect 6193 5593 6227 5627
rect 6227 5593 6236 5627
rect 6184 5584 6236 5593
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 8300 5652 8352 5704
rect 9220 5720 9272 5772
rect 8668 5516 8720 5568
rect 9680 5584 9732 5636
rect 9312 5516 9364 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 3056 5312 3108 5364
rect 3424 5312 3476 5364
rect 2780 5287 2832 5296
rect 2780 5253 2797 5287
rect 2797 5253 2832 5287
rect 2780 5244 2832 5253
rect 3332 5244 3384 5296
rect 4068 5244 4120 5296
rect 4988 5244 5040 5296
rect 5724 5244 5776 5296
rect 1216 5176 1268 5228
rect 2872 5219 2924 5228
rect 2872 5185 2881 5219
rect 2881 5185 2915 5219
rect 2915 5185 2924 5219
rect 2872 5176 2924 5185
rect 3056 5219 3108 5228
rect 3056 5185 3065 5219
rect 3065 5185 3099 5219
rect 3099 5185 3108 5219
rect 3056 5176 3108 5185
rect 3424 5176 3476 5228
rect 6644 5312 6696 5364
rect 6276 5244 6328 5296
rect 7748 5355 7800 5364
rect 7748 5321 7757 5355
rect 7757 5321 7791 5355
rect 7791 5321 7800 5355
rect 7748 5312 7800 5321
rect 8300 5312 8352 5364
rect 8852 5312 8904 5364
rect 9312 5312 9364 5364
rect 9680 5312 9732 5364
rect 10968 5355 11020 5364
rect 10968 5321 10977 5355
rect 10977 5321 11011 5355
rect 11011 5321 11020 5355
rect 10968 5312 11020 5321
rect 9496 5287 9548 5296
rect 9496 5253 9505 5287
rect 9505 5253 9539 5287
rect 9539 5253 9548 5287
rect 9496 5244 9548 5253
rect 3884 5108 3936 5160
rect 1400 5040 1452 5092
rect 4804 5108 4856 5160
rect 5080 5108 5132 5160
rect 7932 5219 7984 5228
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 8392 5176 8444 5228
rect 8484 5176 8536 5228
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 6460 5040 6512 5092
rect 8576 5108 8628 5160
rect 9220 5151 9272 5160
rect 9220 5117 9229 5151
rect 9229 5117 9263 5151
rect 9263 5117 9272 5151
rect 9220 5108 9272 5117
rect 8484 5040 8536 5092
rect 8760 5040 8812 5092
rect 4712 4972 4764 5024
rect 6184 5015 6236 5024
rect 6184 4981 6193 5015
rect 6193 4981 6227 5015
rect 6227 4981 6236 5015
rect 6184 4972 6236 4981
rect 6368 5015 6420 5024
rect 6368 4981 6377 5015
rect 6377 4981 6411 5015
rect 6411 4981 6420 5015
rect 6368 4972 6420 4981
rect 7380 4972 7432 5024
rect 8668 4972 8720 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 2872 4768 2924 4820
rect 7656 4768 7708 4820
rect 9680 4768 9732 4820
rect 4068 4700 4120 4752
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 4712 4632 4764 4684
rect 7380 4675 7432 4684
rect 7380 4641 7389 4675
rect 7389 4641 7423 4675
rect 7423 4641 7432 4675
rect 7380 4632 7432 4641
rect 5448 4564 5500 4616
rect 6736 4607 6788 4616
rect 6736 4573 6745 4607
rect 6745 4573 6779 4607
rect 6779 4573 6788 4607
rect 6736 4564 6788 4573
rect 1676 4539 1728 4548
rect 1676 4505 1685 4539
rect 1685 4505 1719 4539
rect 1719 4505 1728 4539
rect 1676 4496 1728 4505
rect 3148 4496 3200 4548
rect 6092 4496 6144 4548
rect 7564 4496 7616 4548
rect 8116 4564 8168 4616
rect 8484 4607 8536 4616
rect 8484 4573 8493 4607
rect 8493 4573 8527 4607
rect 8527 4573 8536 4607
rect 8484 4564 8536 4573
rect 8576 4607 8628 4616
rect 8576 4573 8585 4607
rect 8585 4573 8619 4607
rect 8619 4573 8628 4607
rect 8576 4564 8628 4573
rect 7012 4428 7064 4480
rect 7472 4428 7524 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 1676 4224 1728 4276
rect 2872 4224 2924 4276
rect 3056 4224 3108 4276
rect 1584 4156 1636 4208
rect 4068 4156 4120 4208
rect 1216 4088 1268 4140
rect 1308 4020 1360 4072
rect 3056 4088 3108 4140
rect 3240 4131 3292 4140
rect 3240 4097 3249 4131
rect 3249 4097 3283 4131
rect 3283 4097 3292 4131
rect 3240 4088 3292 4097
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 4804 4224 4856 4276
rect 6368 4224 6420 4276
rect 6736 4224 6788 4276
rect 6184 4156 6236 4208
rect 7012 4199 7064 4208
rect 7012 4165 7021 4199
rect 7021 4165 7055 4199
rect 7055 4165 7064 4199
rect 7012 4156 7064 4165
rect 7656 4156 7708 4208
rect 8576 4224 8628 4276
rect 9220 4156 9272 4208
rect 2872 4020 2924 4072
rect 3884 4020 3936 4072
rect 4804 4020 4856 4072
rect 5264 4020 5316 4072
rect 7564 4020 7616 4072
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 2780 3884 2832 3936
rect 5264 3884 5316 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 1216 3680 1268 3732
rect 2044 3680 2096 3732
rect 1860 3544 1912 3596
rect 1124 3476 1176 3528
rect 2044 3519 2096 3528
rect 2044 3485 2053 3519
rect 2053 3485 2087 3519
rect 2087 3485 2096 3519
rect 2044 3476 2096 3485
rect 2780 3612 2832 3664
rect 3976 3680 4028 3732
rect 3148 3612 3200 3664
rect 5724 3612 5776 3664
rect 5264 3587 5316 3596
rect 5264 3553 5273 3587
rect 5273 3553 5307 3587
rect 5307 3553 5316 3587
rect 5264 3544 5316 3553
rect 5356 3587 5408 3596
rect 5356 3553 5365 3587
rect 5365 3553 5399 3587
rect 5399 3553 5408 3587
rect 5356 3544 5408 3553
rect 4804 3476 4856 3528
rect 6276 3476 6328 3528
rect 1768 3340 1820 3392
rect 3240 3451 3292 3460
rect 3240 3417 3249 3451
rect 3249 3417 3283 3451
rect 3283 3417 3292 3451
rect 3240 3408 3292 3417
rect 2688 3340 2740 3392
rect 2872 3340 2924 3392
rect 4068 3408 4120 3460
rect 7472 3408 7524 3460
rect 4712 3340 4764 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 3240 3136 3292 3188
rect 4804 3136 4856 3188
rect 6276 3136 6328 3188
rect 9680 3136 9732 3188
rect 1124 3068 1176 3120
rect 2872 3111 2924 3120
rect 2872 3077 2881 3111
rect 2881 3077 2915 3111
rect 2915 3077 2924 3111
rect 2872 3068 2924 3077
rect 3148 3068 3200 3120
rect 4712 3111 4764 3120
rect 4712 3077 4721 3111
rect 4721 3077 4755 3111
rect 4755 3077 4764 3111
rect 4712 3068 4764 3077
rect 5724 3068 5776 3120
rect 9404 3068 9456 3120
rect 1308 3000 1360 3052
rect 9220 3043 9272 3052
rect 9220 3009 9229 3043
rect 9229 3009 9263 3043
rect 9263 3009 9272 3043
rect 9220 3000 9272 3009
rect 2412 2932 2464 2984
rect 3240 2796 3292 2848
rect 3516 2796 3568 2848
rect 10968 2839 11020 2848
rect 10968 2805 10977 2839
rect 10977 2805 11011 2839
rect 11011 2805 11020 2839
rect 10968 2796 11020 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 2780 2592 2832 2644
rect 3332 2592 3384 2644
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 2412 2456 2464 2508
rect 10968 2431 11020 2440
rect 10968 2397 10977 2431
rect 10977 2397 11011 2431
rect 11011 2397 11020 2431
rect 10968 2388 11020 2397
rect 1768 2320 1820 2372
rect 3516 2320 3568 2372
rect 10692 2363 10744 2372
rect 10692 2329 10701 2363
rect 10701 2329 10735 2363
rect 10735 2329 10744 2363
rect 10692 2320 10744 2329
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 1306 12336 1362 12345
rect 1306 12271 1362 12280
rect 1320 11830 1348 12271
rect 10690 12064 10746 12073
rect 4874 11996 5182 12005
rect 10690 11999 10746 12008
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 1308 11824 1360 11830
rect 1214 11792 1270 11801
rect 1124 11756 1176 11762
rect 1308 11766 1360 11772
rect 1214 11727 1270 11736
rect 1860 11756 1912 11762
rect 1124 11698 1176 11704
rect 1136 11257 1164 11698
rect 1228 11694 1256 11727
rect 1860 11698 1912 11704
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 1216 11688 1268 11694
rect 1216 11630 1268 11636
rect 1122 11248 1178 11257
rect 1122 11183 1178 11192
rect 1872 11014 1900 11698
rect 2424 11558 2452 11698
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1122 10704 1178 10713
rect 1872 10674 1900 10950
rect 1122 10639 1178 10648
rect 1308 10668 1360 10674
rect 1136 10130 1164 10639
rect 1308 10610 1360 10616
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1320 10169 1348 10610
rect 2516 10470 2544 11698
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2792 11082 2820 11290
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 1860 10464 1912 10470
rect 1860 10406 1912 10412
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 1306 10160 1362 10169
rect 1124 10124 1176 10130
rect 1306 10095 1362 10104
rect 1124 10066 1176 10072
rect 1872 10062 1900 10406
rect 1216 10056 1268 10062
rect 1216 9998 1268 10004
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1228 9625 1256 9998
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1596 9722 1624 9862
rect 1584 9716 1636 9722
rect 1584 9658 1636 9664
rect 1214 9616 1270 9625
rect 1214 9551 1270 9560
rect 1308 9580 1360 9586
rect 1308 9522 1360 9528
rect 1320 9081 1348 9522
rect 1306 9072 1362 9081
rect 1306 9007 1362 9016
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1032 8968 1084 8974
rect 1032 8910 1084 8916
rect 1044 8566 1072 8910
rect 1032 8560 1084 8566
rect 1030 8528 1032 8537
rect 1084 8528 1086 8537
rect 1030 8463 1086 8472
rect 1308 8492 1360 8498
rect 1308 8434 1360 8440
rect 1320 7993 1348 8434
rect 1306 7984 1362 7993
rect 1306 7919 1362 7928
rect 1308 7880 1360 7886
rect 1308 7822 1360 7828
rect 1320 7449 1348 7822
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1596 7546 1624 7686
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1688 7478 1716 8978
rect 1952 8900 2004 8906
rect 1952 8842 2004 8848
rect 1964 8634 1992 8842
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1676 7472 1728 7478
rect 1306 7440 1362 7449
rect 1676 7414 1728 7420
rect 1306 7375 1362 7384
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1688 7002 1716 7278
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1214 6896 1270 6905
rect 1214 6831 1270 6840
rect 1228 6798 1256 6831
rect 1216 6792 1268 6798
rect 1216 6734 1268 6740
rect 1228 6458 1256 6734
rect 1308 6724 1360 6730
rect 1308 6666 1360 6672
rect 1216 6452 1268 6458
rect 1216 6394 1268 6400
rect 1320 6361 1348 6666
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1306 6352 1362 6361
rect 1216 6316 1268 6322
rect 1306 6287 1362 6296
rect 1216 6258 1268 6264
rect 1228 5817 1256 6258
rect 1400 6180 1452 6186
rect 1400 6122 1452 6128
rect 1214 5808 1270 5817
rect 1214 5743 1270 5752
rect 1308 5704 1360 5710
rect 1308 5646 1360 5652
rect 1320 5273 1348 5646
rect 1306 5264 1362 5273
rect 1216 5228 1268 5234
rect 1306 5199 1362 5208
rect 1216 5170 1268 5176
rect 1228 4729 1256 5170
rect 1412 5098 1440 6122
rect 1872 5642 1900 6598
rect 1860 5636 1912 5642
rect 1860 5578 1912 5584
rect 1400 5092 1452 5098
rect 1400 5034 1452 5040
rect 1214 4720 1270 4729
rect 1214 4655 1270 4664
rect 1412 4622 1440 5034
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1214 4176 1270 4185
rect 1214 4111 1216 4120
rect 1268 4111 1270 4120
rect 1216 4082 1268 4088
rect 1228 3738 1256 4082
rect 1308 4072 1360 4078
rect 1308 4014 1360 4020
rect 1216 3732 1268 3738
rect 1216 3674 1268 3680
rect 1320 3641 1348 4014
rect 1306 3632 1362 3641
rect 1306 3567 1362 3576
rect 1124 3528 1176 3534
rect 1124 3470 1176 3476
rect 1136 3126 1164 3470
rect 1124 3120 1176 3126
rect 1122 3088 1124 3097
rect 1176 3088 1178 3097
rect 1122 3023 1178 3032
rect 1308 3052 1360 3058
rect 1308 2994 1360 3000
rect 1320 2553 1348 2994
rect 1306 2544 1362 2553
rect 1412 2514 1440 4558
rect 1596 4214 1624 4966
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 1688 4282 1716 4490
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1584 4208 1636 4214
rect 1584 4150 1636 4156
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1872 3602 1900 3878
rect 2056 3738 2084 10406
rect 2516 10266 2544 10406
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2700 9994 2728 10542
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2976 9994 3004 10474
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 3068 9602 3096 11494
rect 3160 11234 3188 11494
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3160 11206 3280 11234
rect 3252 11150 3280 11206
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3344 10674 3372 11154
rect 4816 11082 4844 11834
rect 10704 11830 10732 11999
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5460 11098 5488 11154
rect 4804 11076 4856 11082
rect 5460 11070 5580 11098
rect 4804 11018 4856 11024
rect 3608 10736 3660 10742
rect 3608 10678 3660 10684
rect 3884 10736 3936 10742
rect 3884 10678 3936 10684
rect 4816 10690 4844 11018
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5276 10810 5304 10950
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 4896 10736 4948 10742
rect 4816 10684 4896 10690
rect 4816 10678 4948 10684
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3620 10266 3648 10678
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3516 9648 3568 9654
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2608 6914 2636 8230
rect 2792 8022 2820 9590
rect 3068 9574 3280 9602
rect 3516 9590 3568 9596
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 2964 8560 3016 8566
rect 2964 8502 3016 8508
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2884 8090 2912 8366
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 2688 7880 2740 7886
rect 2740 7840 2912 7868
rect 2688 7822 2740 7828
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2792 7206 2820 7686
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2608 6886 2728 6914
rect 2700 6798 2728 6886
rect 2884 6798 2912 7840
rect 2976 7818 3004 8502
rect 3160 8430 3188 9386
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3160 7886 3188 8366
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 2964 7812 3016 7818
rect 2964 7754 3016 7760
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2976 6662 3004 7210
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 3068 6730 3096 7142
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2424 5914 2452 6190
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2792 5302 2820 6394
rect 3148 6384 3200 6390
rect 3148 6326 3200 6332
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2884 5522 2912 5714
rect 2976 5710 3004 6054
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 3056 5568 3108 5574
rect 2884 5494 3004 5522
rect 3056 5510 3108 5516
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2884 4826 2912 5170
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2884 4282 2912 4762
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2976 4162 3004 5494
rect 3068 5370 3096 5510
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 3068 4282 3096 5170
rect 3160 4554 3188 6326
rect 3252 5778 3280 9574
rect 3528 9450 3556 9590
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3424 9444 3476 9450
rect 3424 9386 3476 9392
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3436 8838 3464 9386
rect 3804 9382 3832 9522
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3804 9110 3832 9318
rect 3792 9104 3844 9110
rect 3792 9046 3844 9052
rect 3896 8906 3924 10678
rect 4816 10662 4936 10678
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4080 9586 4108 10406
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4816 10146 4844 10662
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4448 10130 4844 10146
rect 4436 10124 4844 10130
rect 4488 10118 4844 10124
rect 4436 10066 4488 10072
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4172 9586 4200 9862
rect 4264 9654 4292 9862
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4540 9382 4568 9862
rect 4632 9382 4660 9998
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3344 8498 3372 8774
rect 3436 8634 3464 8774
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3896 7750 3924 8842
rect 4080 7954 4108 8978
rect 4724 8294 4752 10118
rect 4908 10062 4936 10406
rect 5276 10266 5304 10542
rect 5552 10538 5580 11070
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 4908 9110 4936 9522
rect 5276 9518 5304 9998
rect 5448 9988 5500 9994
rect 5448 9930 5500 9936
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5276 9178 5304 9454
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 4896 9104 4948 9110
rect 4896 9046 4948 9052
rect 5368 8974 5396 9522
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3896 7478 3924 7686
rect 4356 7546 4384 7754
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 3884 7472 3936 7478
rect 3936 7420 4016 7426
rect 3884 7414 4016 7420
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3700 7404 3752 7410
rect 3896 7398 4016 7414
rect 3700 7346 3752 7352
rect 3424 7268 3476 7274
rect 3424 7210 3476 7216
rect 3436 7002 3464 7210
rect 3528 7206 3556 7346
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3436 5370 3464 6938
rect 3620 6118 3648 7346
rect 3712 6934 3740 7346
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3700 6928 3752 6934
rect 3700 6870 3752 6876
rect 3896 6458 3924 7278
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3332 5296 3384 5302
rect 3252 5244 3332 5250
rect 3252 5238 3384 5244
rect 3252 5222 3372 5238
rect 3436 5234 3464 5306
rect 3424 5228 3476 5234
rect 3148 4548 3200 4554
rect 3148 4490 3200 4496
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 2884 4134 3004 4162
rect 3068 4146 3096 4218
rect 3056 4140 3108 4146
rect 2884 4078 2912 4134
rect 3056 4082 3108 4088
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 2056 3534 2084 3674
rect 2792 3670 2820 3878
rect 3160 3670 3188 4490
rect 3252 4146 3280 5222
rect 3424 5170 3476 5176
rect 3896 5166 3924 6394
rect 3988 6390 4016 7398
rect 5276 7342 5304 8230
rect 5368 7750 5396 8434
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5368 7546 5396 7686
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 2688 3392 2740 3398
rect 2872 3392 2924 3398
rect 2740 3340 2820 3346
rect 2688 3334 2820 3340
rect 2872 3334 2924 3340
rect 1306 2479 1362 2488
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1780 2378 1808 3334
rect 2700 3318 2820 3334
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 2424 2514 2452 2926
rect 2792 2650 2820 3318
rect 2884 3126 2912 3334
rect 3160 3126 3188 3606
rect 3240 3460 3292 3466
rect 3240 3402 3292 3408
rect 3252 3194 3280 3402
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 2872 3120 2924 3126
rect 2872 3062 2924 3068
rect 3148 3120 3200 3126
rect 3148 3062 3200 3068
rect 3160 2938 3188 3062
rect 3160 2910 3280 2938
rect 3252 2854 3280 2910
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 3344 2650 3372 4082
rect 3896 4078 3924 5102
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 3988 3738 4016 6326
rect 4080 5302 4108 7142
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 5460 6662 5488 9930
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5552 8634 5580 9862
rect 5736 9654 5764 11562
rect 10980 11354 11008 11698
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 6460 11280 6512 11286
rect 6460 11222 6512 11228
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 6380 10810 6408 10950
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 5828 9654 5856 10746
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6288 10130 6316 10406
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5632 9512 5684 9518
rect 5630 9480 5632 9489
rect 5724 9512 5776 9518
rect 5684 9480 5686 9489
rect 5724 9454 5776 9460
rect 5630 9415 5686 9424
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5644 8430 5672 9318
rect 5736 9042 5764 9454
rect 5920 9450 5948 9590
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5736 8498 5764 8978
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5736 6798 5764 8434
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 4080 4758 4108 5238
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 4080 4214 4108 4694
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3988 3482 4016 3674
rect 3988 3466 4108 3482
rect 3988 3460 4120 3466
rect 3988 3454 4068 3460
rect 4068 3402 4120 3408
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 2412 2508 2464 2514
rect 2412 2450 2464 2456
rect 3528 2378 3556 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 1768 2372 1820 2378
rect 1768 2314 1820 2320
rect 3516 2372 3568 2378
rect 3516 2314 3568 2320
rect 4632 2009 4660 6598
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4724 5030 4752 6054
rect 4816 5914 4844 6190
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4988 5296 5040 5302
rect 5040 5244 5120 5250
rect 4988 5238 5120 5244
rect 5000 5222 5120 5238
rect 5092 5166 5120 5222
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4724 4690 4752 4966
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 4816 4282 4844 5102
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 5276 4078 5304 5714
rect 5460 4622 5488 6598
rect 5736 5778 5764 6734
rect 5920 6118 5948 7346
rect 6012 6322 6040 8910
rect 6196 8430 6224 9454
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6196 7410 6224 8366
rect 6288 7954 6316 10066
rect 6472 9518 6500 11222
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6656 10742 6684 11086
rect 6644 10736 6696 10742
rect 6644 10678 6696 10684
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6644 10192 6696 10198
rect 6644 10134 6696 10140
rect 6656 9926 6684 10134
rect 6748 9926 6776 10406
rect 7300 10266 7328 10542
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6656 9722 6684 9862
rect 6748 9722 6776 9862
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6460 9512 6512 9518
rect 6458 9480 6460 9489
rect 6512 9480 6514 9489
rect 6458 9415 6514 9424
rect 6656 8650 6684 9522
rect 6564 8634 6684 8650
rect 6564 8628 6696 8634
rect 6564 8622 6644 8628
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6380 7954 6408 8230
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6564 7886 6592 8622
rect 6644 8570 6696 8576
rect 6748 8566 6776 9658
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6932 9178 6960 9522
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 7484 9042 7512 11154
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 7760 10198 7788 11018
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8024 10736 8076 10742
rect 8024 10678 8076 10684
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7760 9722 7788 9862
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 7852 9602 7880 9862
rect 7760 9574 7880 9602
rect 7944 9586 7972 10542
rect 7932 9580 7984 9586
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 6736 8560 6788 8566
rect 6656 8508 6736 8514
rect 6656 8502 6788 8508
rect 6656 8486 6776 8502
rect 6656 8022 6684 8486
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6748 8090 6776 8366
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6656 6866 6684 7958
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 6932 6458 6960 6666
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5920 5710 5948 6054
rect 6472 5778 6500 6258
rect 6644 5840 6696 5846
rect 6644 5782 6696 5788
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 5724 5296 5776 5302
rect 5724 5238 5776 5244
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 5264 4072 5316 4078
rect 5316 4020 5396 4026
rect 5264 4014 5396 4020
rect 4816 3534 4844 4014
rect 5276 3998 5396 4014
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5276 3602 5304 3878
rect 5368 3602 5396 3998
rect 5736 3670 5764 5238
rect 6104 4554 6132 5578
rect 6196 5030 6224 5578
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6092 4548 6144 4554
rect 6092 4490 6144 4496
rect 6196 4214 6224 4966
rect 6184 4208 6236 4214
rect 6184 4150 6236 4156
rect 5724 3664 5776 3670
rect 5724 3606 5776 3612
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4724 3126 4752 3334
rect 4816 3194 4844 3470
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 5736 3126 5764 3606
rect 6288 3534 6316 5238
rect 6472 5098 6500 5714
rect 6656 5370 6684 5782
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6460 5092 6512 5098
rect 6460 5034 6512 5040
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 6380 4282 6408 4966
rect 7392 4690 7420 4966
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6748 4282 6776 4558
rect 7484 4486 7512 8978
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7668 6730 7696 8502
rect 7656 6724 7708 6730
rect 7656 6666 7708 6672
rect 7668 4826 7696 6666
rect 7760 6322 7788 9574
rect 7932 9522 7984 9528
rect 7944 8498 7972 9522
rect 8036 8906 8064 10678
rect 8128 10062 8156 10950
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8404 10062 8432 10406
rect 8588 10062 8616 10542
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8128 9926 8156 9998
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 7852 6322 7880 8298
rect 8128 7478 8156 9318
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8220 8362 8248 8842
rect 8312 8634 8340 9386
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8680 8498 8708 11018
rect 8772 9654 8800 11086
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9508 10810 9536 11018
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8772 8974 8800 9590
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7944 6322 7972 6598
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 7760 5370 7788 6122
rect 7748 5364 7800 5370
rect 7748 5306 7800 5312
rect 7944 5234 7972 6258
rect 8036 5778 8064 6394
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8680 6202 8708 8434
rect 8772 7410 8800 8910
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 8128 5710 8156 6054
rect 8312 5846 8340 6190
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8300 5840 8352 5846
rect 8300 5782 8352 5788
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 7024 4214 7052 4422
rect 7012 4208 7064 4214
rect 7012 4150 7064 4156
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6288 3194 6316 3470
rect 7484 3466 7512 4422
rect 7576 4078 7604 4490
rect 7668 4214 7696 4762
rect 8128 4622 8156 5646
rect 8312 5370 8340 5646
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8404 5234 8432 6054
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8496 5234 8524 5782
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8588 5166 8616 6190
rect 8680 6174 8800 6202
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8680 5846 8708 6054
rect 8668 5840 8720 5846
rect 8668 5782 8720 5788
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8484 5092 8536 5098
rect 8484 5034 8536 5040
rect 8496 4622 8524 5034
rect 8588 4622 8616 5102
rect 8680 5030 8708 5510
rect 8772 5098 8800 6174
rect 8864 5914 8892 6258
rect 9048 5914 9076 9998
rect 9232 9450 9260 10610
rect 9324 9518 9352 10610
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9220 9444 9272 9450
rect 9220 9386 9272 9392
rect 9324 8566 9352 9454
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9324 5914 9352 6054
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 8864 5370 8892 5850
rect 9220 5772 9272 5778
rect 9220 5714 9272 5720
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 9232 5166 9260 5714
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9324 5370 9352 5510
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8588 4282 8616 4558
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 9232 4214 9260 5102
rect 7656 4208 7708 4214
rect 7656 4150 7708 4156
rect 9220 4208 9272 4214
rect 9220 4150 9272 4156
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7472 3460 7524 3466
rect 7472 3402 7524 3408
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 5724 3120 5776 3126
rect 5724 3062 5776 3068
rect 9232 3058 9260 4150
rect 9416 3126 9444 9862
rect 9968 8974 9996 11018
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9968 7478 9996 8910
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 10968 7200 11020 7206
rect 10782 7168 10838 7177
rect 10968 7142 11020 7148
rect 10782 7103 10838 7112
rect 10796 6866 10824 7103
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10980 6798 11008 7142
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9508 5302 9536 6054
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9692 5370 9720 5578
rect 10980 5370 11008 6326
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9692 4826 9720 5306
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9692 3194 9720 4762
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 10980 2446 11008 2790
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 10692 2372 10744 2378
rect 10692 2314 10744 2320
rect 10704 2281 10732 2314
rect 10690 2272 10746 2281
rect 4874 2204 5182 2213
rect 10690 2207 10746 2216
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 4618 2000 4674 2009
rect 4618 1935 4674 1944
<< via2 >>
rect 1306 12280 1362 12336
rect 10690 12008 10746 12064
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 1214 11736 1270 11792
rect 1122 11192 1178 11248
rect 1122 10648 1178 10704
rect 1306 10104 1362 10160
rect 1214 9560 1270 9616
rect 1306 9016 1362 9072
rect 1030 8508 1032 8528
rect 1032 8508 1084 8528
rect 1084 8508 1086 8528
rect 1030 8472 1086 8508
rect 1306 7928 1362 7984
rect 1306 7384 1362 7440
rect 1214 6840 1270 6896
rect 1306 6296 1362 6352
rect 1214 5752 1270 5808
rect 1306 5208 1362 5264
rect 1214 4664 1270 4720
rect 1214 4140 1270 4176
rect 1214 4120 1216 4140
rect 1216 4120 1268 4140
rect 1268 4120 1270 4140
rect 1306 3576 1362 3632
rect 1122 3068 1124 3088
rect 1124 3068 1176 3088
rect 1176 3068 1178 3088
rect 1122 3032 1178 3068
rect 1306 2488 1362 2544
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 5630 9460 5632 9480
rect 5632 9460 5684 9480
rect 5684 9460 5686 9480
rect 5630 9424 5686 9460
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 6458 9460 6460 9480
rect 6460 9460 6512 9480
rect 6512 9460 6514 9480
rect 6458 9424 6514 9460
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 10782 7112 10838 7168
rect 10690 2216 10746 2272
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 4618 1944 4674 2000
<< metal3 >>
rect 0 12338 800 12368
rect 1301 12338 1367 12341
rect 0 12336 1367 12338
rect 0 12280 1306 12336
rect 1362 12280 1367 12336
rect 0 12278 1367 12280
rect 0 12248 800 12278
rect 1301 12275 1367 12278
rect 10685 12066 10751 12069
rect 11702 12066 12502 12096
rect 10685 12064 12502 12066
rect 10685 12008 10690 12064
rect 10746 12008 12502 12064
rect 10685 12006 12502 12008
rect 10685 12003 10751 12006
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 11702 11976 12502 12006
rect 4870 11935 5186 11936
rect 0 11794 800 11824
rect 1209 11794 1275 11797
rect 0 11792 1275 11794
rect 0 11736 1214 11792
rect 1270 11736 1275 11792
rect 0 11734 1275 11736
rect 0 11704 800 11734
rect 1209 11731 1275 11734
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 0 11250 800 11280
rect 1117 11250 1183 11253
rect 0 11248 1183 11250
rect 0 11192 1122 11248
rect 1178 11192 1183 11248
rect 0 11190 1183 11192
rect 0 11160 800 11190
rect 1117 11187 1183 11190
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 0 10706 800 10736
rect 1117 10706 1183 10709
rect 0 10704 1183 10706
rect 0 10648 1122 10704
rect 1178 10648 1183 10704
rect 0 10646 1183 10648
rect 0 10616 800 10646
rect 1117 10643 1183 10646
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 0 10162 800 10192
rect 1301 10162 1367 10165
rect 0 10160 1367 10162
rect 0 10104 1306 10160
rect 1362 10104 1367 10160
rect 0 10102 1367 10104
rect 0 10072 800 10102
rect 1301 10099 1367 10102
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 0 9618 800 9648
rect 1209 9618 1275 9621
rect 0 9616 1275 9618
rect 0 9560 1214 9616
rect 1270 9560 1275 9616
rect 0 9558 1275 9560
rect 0 9528 800 9558
rect 1209 9555 1275 9558
rect 5625 9482 5691 9485
rect 6453 9482 6519 9485
rect 5625 9480 6519 9482
rect 5625 9424 5630 9480
rect 5686 9424 6458 9480
rect 6514 9424 6519 9480
rect 5625 9422 6519 9424
rect 5625 9419 5691 9422
rect 6453 9419 6519 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 0 9074 800 9104
rect 1301 9074 1367 9077
rect 0 9072 1367 9074
rect 0 9016 1306 9072
rect 1362 9016 1367 9072
rect 0 9014 1367 9016
rect 0 8984 800 9014
rect 1301 9011 1367 9014
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 0 8530 800 8560
rect 1025 8530 1091 8533
rect 0 8528 1091 8530
rect 0 8472 1030 8528
rect 1086 8472 1091 8528
rect 0 8470 1091 8472
rect 0 8440 800 8470
rect 1025 8467 1091 8470
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 0 7986 800 8016
rect 1301 7986 1367 7989
rect 0 7984 1367 7986
rect 0 7928 1306 7984
rect 1362 7928 1367 7984
rect 0 7926 1367 7928
rect 0 7896 800 7926
rect 1301 7923 1367 7926
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 0 7442 800 7472
rect 1301 7442 1367 7445
rect 0 7440 1367 7442
rect 0 7384 1306 7440
rect 1362 7384 1367 7440
rect 0 7382 1367 7384
rect 0 7352 800 7382
rect 1301 7379 1367 7382
rect 10777 7170 10843 7173
rect 11702 7170 12502 7200
rect 10777 7168 12502 7170
rect 10777 7112 10782 7168
rect 10838 7112 12502 7168
rect 10777 7110 12502 7112
rect 10777 7107 10843 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 11702 7080 12502 7110
rect 4210 7039 4526 7040
rect 0 6898 800 6928
rect 1209 6898 1275 6901
rect 0 6896 1275 6898
rect 0 6840 1214 6896
rect 1270 6840 1275 6896
rect 0 6838 1275 6840
rect 0 6808 800 6838
rect 1209 6835 1275 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 0 6354 800 6384
rect 1301 6354 1367 6357
rect 0 6352 1367 6354
rect 0 6296 1306 6352
rect 1362 6296 1367 6352
rect 0 6294 1367 6296
rect 0 6264 800 6294
rect 1301 6291 1367 6294
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 0 5810 800 5840
rect 1209 5810 1275 5813
rect 0 5808 1275 5810
rect 0 5752 1214 5808
rect 1270 5752 1275 5808
rect 0 5750 1275 5752
rect 0 5720 800 5750
rect 1209 5747 1275 5750
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 0 5266 800 5296
rect 1301 5266 1367 5269
rect 0 5264 1367 5266
rect 0 5208 1306 5264
rect 1362 5208 1367 5264
rect 0 5206 1367 5208
rect 0 5176 800 5206
rect 1301 5203 1367 5206
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 0 4722 800 4752
rect 1209 4722 1275 4725
rect 0 4720 1275 4722
rect 0 4664 1214 4720
rect 1270 4664 1275 4720
rect 0 4662 1275 4664
rect 0 4632 800 4662
rect 1209 4659 1275 4662
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 0 4178 800 4208
rect 1209 4178 1275 4181
rect 0 4176 1275 4178
rect 0 4120 1214 4176
rect 1270 4120 1275 4176
rect 0 4118 1275 4120
rect 0 4088 800 4118
rect 1209 4115 1275 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 0 3634 800 3664
rect 1301 3634 1367 3637
rect 0 3632 1367 3634
rect 0 3576 1306 3632
rect 1362 3576 1367 3632
rect 0 3574 1367 3576
rect 0 3544 800 3574
rect 1301 3571 1367 3574
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 0 3090 800 3120
rect 1117 3090 1183 3093
rect 0 3088 1183 3090
rect 0 3032 1122 3088
rect 1178 3032 1183 3088
rect 0 3030 1183 3032
rect 0 3000 800 3030
rect 1117 3027 1183 3030
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 0 2546 800 2576
rect 1301 2546 1367 2549
rect 0 2544 1367 2546
rect 0 2488 1306 2544
rect 1362 2488 1367 2544
rect 0 2486 1367 2488
rect 0 2456 800 2486
rect 1301 2483 1367 2486
rect 10685 2274 10751 2277
rect 11702 2274 12502 2304
rect 10685 2272 12502 2274
rect 10685 2216 10690 2272
rect 10746 2216 12502 2272
rect 10685 2214 12502 2216
rect 10685 2211 10751 2214
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 11702 2184 12502 2214
rect 4870 2143 5186 2144
rect 0 2002 800 2032
rect 4613 2002 4679 2005
rect 0 2000 4679 2002
rect 0 1944 4618 2000
rect 4674 1944 4679 2000
rect 0 1942 4679 1944
rect 0 1912 800 1942
rect 4613 1939 4679 1942
<< via3 >>
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 11456 4528 12016
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 12000 5188 12016
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _046_
timestamp -25199
transform 1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _047_
timestamp -25199
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _048_
timestamp -25199
transform -1 0 2116 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _049_
timestamp -25199
transform -1 0 2944 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _050_
timestamp -25199
transform -1 0 3496 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _051_
timestamp -25199
transform 1 0 2116 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _052_
timestamp -25199
transform 1 0 8004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _053_
timestamp -25199
transform 1 0 7544 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _054_
timestamp -25199
transform -1 0 8832 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _055_
timestamp -25199
transform 1 0 2668 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _056_
timestamp -25199
transform -1 0 8740 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _057_
timestamp -25199
transform 1 0 7176 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _058_
timestamp -25199
transform -1 0 8188 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _059_
timestamp -25199
transform 1 0 7360 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _060_
timestamp -25199
transform -1 0 9016 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _061_
timestamp -25199
transform -1 0 8832 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _062_
timestamp -25199
transform 1 0 8924 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _063_
timestamp -25199
transform -1 0 8832 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _064_
timestamp -25199
transform -1 0 6256 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _065_
timestamp -25199
transform 1 0 2484 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _066_
timestamp -25199
transform -1 0 2484 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _067_
timestamp -25199
transform -1 0 4784 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _068_
timestamp -25199
transform 1 0 4784 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _069_
timestamp -25199
transform 1 0 2944 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _070_
timestamp -25199
transform 1 0 2116 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _071_
timestamp -25199
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _072_
timestamp -25199
transform 1 0 5060 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _073_
timestamp -25199
transform -1 0 3312 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _074_
timestamp -25199
transform 1 0 2576 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _075_
timestamp -25199
transform 1 0 5796 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _076_
timestamp -25199
transform 1 0 4968 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _077_
timestamp -25199
transform 1 0 3220 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _078_
timestamp -25199
transform 1 0 2208 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _079_
timestamp -25199
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _080_
timestamp -25199
transform 1 0 4692 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _081_
timestamp -25199
transform 1 0 2484 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _082_
timestamp -25199
transform 1 0 2392 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _083_
timestamp -25199
transform -1 0 5796 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _084_
timestamp -25199
transform -1 0 6900 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _085_
timestamp -25199
transform -1 0 3680 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _086_
timestamp -25199
transform 1 0 3772 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _087_
timestamp -25199
transform -1 0 7084 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _088_
timestamp -25199
transform 1 0 7268 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _089_
timestamp -25199
transform -1 0 5336 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _090_
timestamp -25199
transform 1 0 5152 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _091_
timestamp -25199
transform -1 0 9660 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _092_
timestamp -25199
transform 1 0 2576 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _093_
timestamp -25199
transform 1 0 1380 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _094_
timestamp -25199
transform 1 0 4416 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _095_
timestamp -25199
transform 1 0 1380 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _096_
timestamp -25199
transform 1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _097_
timestamp -25199
transform 1 0 2116 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _098_
timestamp -25199
transform 1 0 4416 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _099_
timestamp -25199
transform 1 0 1380 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _100_
timestamp -25199
transform 1 0 4048 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _101_
timestamp -25199
transform 1 0 1656 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _102_
timestamp -25199
transform 1 0 6348 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _103_
timestamp -25199
transform 1 0 3312 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _104_
timestamp -25199
transform 1 0 6348 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _105_
timestamp -25199
transform 1 0 4600 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _106_
timestamp -25199
transform -1 0 3220 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _107_
timestamp -25199
transform 1 0 9200 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _108_
timestamp -25199
transform 1 0 9200 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _109_
timestamp -25199
transform 1 0 9200 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _110_
timestamp -25199
transform 1 0 6716 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _111_
timestamp -25199
transform 1 0 6624 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _112_
timestamp -25199
transform 1 0 8924 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _113_
timestamp -25199
transform 1 0 9200 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _114_
timestamp -25199
transform -1 0 8832 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp -25199
transform -1 0 4784 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp -25199
transform -1 0 1840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp -25199
transform -1 0 1840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp -25199
transform -1 0 1840 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp -25199
transform -1 0 2300 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp -25199
transform -1 0 1840 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp -25199
transform -1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp -25199
transform -1 0 3588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp -25199
transform -1 0 2116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp -25199
transform -1 0 1840 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp -25199
transform -1 0 1840 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp -25199
transform -1 0 1840 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp -25199
transform -1 0 2024 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp -25199
transform -1 0 2116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp -25199
transform -1 0 1840 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp -25199
transform -1 0 1840 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp -25199
transform -1 0 2024 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp -25199
transform -1 0 3404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp -25199
transform -1 0 2024 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -25199
transform 1 0 4784 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp -25199
transform 1 0 5060 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp -25199
transform 1 0 5428 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp -25199
transform 1 0 4508 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout23
timestamp -25199
transform 1 0 3036 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout24
timestamp -25199
transform -1 0 4048 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout25
timestamp -25199
transform 1 0 8188 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  fanout26
timestamp -25199
transform 1 0 4048 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout27
timestamp -25199
transform -1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout28
timestamp -25199
transform -1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout29
timestamp -25199
transform -1 0 8188 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout30
timestamp -25199
transform 1 0 8740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout31
timestamp -25199
transform 1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout32
timestamp -25199
transform 1 0 8188 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout33
timestamp -25199
transform -1 0 6716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout34
timestamp -25199
transform 1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout35
timestamp -25199
transform -1 0 2668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout36
timestamp -25199
transform 1 0 6348 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout37
timestamp -25199
transform -1 0 5520 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout38
timestamp -25199
transform -1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout39
timestamp -25199
transform -1 0 4140 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout40
timestamp -25199
transform 1 0 7912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout41
timestamp -25199
transform 1 0 8924 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout42
timestamp -25199
transform 1 0 3128 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp -25199
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -25199
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636943256
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636943256
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -25199
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636943256
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636943256
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -25199
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636943256
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp -25199
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101
timestamp -25199
transform 1 0 10396 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_10
timestamp -25199
transform 1 0 2024 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636943256
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636943256
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_81
timestamp -25199
transform 1 0 8556 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_87
timestamp -25199
transform 1 0 9108 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp -25199
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_37
timestamp -25199
transform 1 0 4508 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_49
timestamp 1636943256
transform 1 0 5612 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_61
timestamp 1636943256
transform 1 0 6716 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_73
timestamp -25199
transform 1 0 7820 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp -25199
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636943256
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_97
timestamp -25199
transform 1 0 10028 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_105
timestamp -25199
transform 1 0 10764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_28
timestamp -25199
transform 1 0 3680 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_40
timestamp -25199
transform 1 0 4784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp -25199
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp -25199
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636943256
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636943256
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_105
timestamp -25199
transform 1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp -25199
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -25199
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp -25199
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_63
timestamp -25199
transform 1 0 6900 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_73
timestamp -25199
transform 1 0 7820 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636943256
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_97
timestamp -25199
transform 1 0 10028 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_105
timestamp -25199
transform 1 0 10764 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_8
timestamp -25199
transform 1 0 1840 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_24
timestamp 1636943256
transform 1 0 3312 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_65
timestamp -25199
transform 1 0 7084 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_77
timestamp -25199
transform 1 0 8188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_86
timestamp -25199
transform 1 0 9016 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_8
timestamp -25199
transform 1 0 1840 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp -25199
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636943256
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_41
timestamp -25199
transform 1 0 4876 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_59
timestamp -25199
transform 1 0 6532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_67
timestamp -25199
transform 1 0 7268 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_105
timestamp -25199
transform 1 0 10764 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_10
timestamp -25199
transform 1 0 2024 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_31
timestamp -25199
transform 1 0 3956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_35
timestamp -25199
transform 1 0 4324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_67
timestamp -25199
transform 1 0 7268 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_84
timestamp -25199
transform 1 0 8832 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_92
timestamp 1636943256
transform 1 0 9568 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_104
timestamp -25199
transform 1 0 10672 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_11
timestamp -25199
transform 1 0 2116 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp -25199
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp -25199
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_37
timestamp -25199
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp -25199
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636943256
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_97
timestamp -25199
transform 1 0 10028 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_101
timestamp -25199
transform 1 0 10396 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_31
timestamp -25199
transform 1 0 3956 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636943256
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636943256
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_81
timestamp -25199
transform 1 0 8556 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_87
timestamp -25199
transform 1 0 9108 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_8
timestamp -25199
transform 1 0 1840 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_14
timestamp -25199
transform 1 0 2392 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp -25199
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -25199
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp -25199
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_52
timestamp -25199
transform 1 0 5888 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_63
timestamp 1636943256
transform 1 0 6900 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_75
timestamp -25199
transform 1 0 8004 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp -25199
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636943256
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp -25199
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_105
timestamp -25199
transform 1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_10
timestamp -25199
transform 1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_23
timestamp 1636943256
transform 1 0 3220 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_35
timestamp -25199
transform 1 0 4324 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp -25199
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp -25199
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_86
timestamp 1636943256
transform 1 0 9016 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_98
timestamp -25199
transform 1 0 10120 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_106
timestamp -25199
transform 1 0 10856 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp -25199
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636943256
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636943256
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_53
timestamp -25199
transform 1 0 5980 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_61
timestamp -25199
transform 1 0 6716 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_95
timestamp 1636943256
transform 1 0 9844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_107
timestamp -25199
transform 1 0 10948 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_8
timestamp 1636943256
transform 1 0 1840 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_35
timestamp -25199
transform 1 0 4324 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_65
timestamp 1636943256
transform 1 0 7084 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_77
timestamp 1636943256
transform 1 0 8188 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_89
timestamp 1636943256
transform 1 0 9292 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_101
timestamp -25199
transform 1 0 10396 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_107
timestamp -25199
transform 1 0 10948 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_13
timestamp -25199
transform 1 0 2300 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp -25199
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_46
timestamp -25199
transform 1 0 5336 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1636943256
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_97
timestamp -25199
transform 1 0 10028 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_105
timestamp -25199
transform 1 0 10764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_23
timestamp -25199
transform 1 0 3220 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp -25199
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1636943256
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_105
timestamp -25199
transform 1 0 10764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp -25199
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_29
timestamp -25199
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_37
timestamp -25199
transform 1 0 4508 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_61
timestamp 1636943256
transform 1 0 6716 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp -25199
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_85
timestamp -25199
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp -25199
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_29
timestamp 1636943256
transform 1 0 3772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_41
timestamp 1636943256
transform 1 0 4876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp -25199
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636943256
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1636943256
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_81
timestamp -25199
transform 1 0 8556 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_85
timestamp 1636943256
transform 1 0 8924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_97
timestamp -25199
transform 1 0 10028 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_101
timestamp -25199
transform 1 0 10396 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp -25199
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp -25199
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp -25199
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp -25199
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp -25199
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp -25199
transform -1 0 1932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp -25199
transform -1 0 2944 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp -25199
transform -1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp -25199
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp -25199
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp -25199
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp -25199
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp -25199
transform -1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp -25199
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp -25199
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp -25199
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp -25199
transform -1 0 3220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp -25199
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  output19
timestamp -25199
transform -1 0 11040 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output20
timestamp -25199
transform -1 0 11040 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output21
timestamp -25199
transform -1 0 1932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output22
timestamp -25199
transform -1 0 11040 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_18
timestamp -25199
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -25199
transform -1 0 11316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_19
timestamp -25199
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -25199
transform -1 0 11316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_20
timestamp -25199
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -25199
transform -1 0 11316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_21
timestamp -25199
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -25199
transform -1 0 11316 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_22
timestamp -25199
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -25199
transform -1 0 11316 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_23
timestamp -25199
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -25199
transform -1 0 11316 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_24
timestamp -25199
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -25199
transform -1 0 11316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_25
timestamp -25199
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -25199
transform -1 0 11316 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_26
timestamp -25199
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -25199
transform -1 0 11316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_27
timestamp -25199
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -25199
transform -1 0 11316 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_28
timestamp -25199
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -25199
transform -1 0 11316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_29
timestamp -25199
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -25199
transform -1 0 11316 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_30
timestamp -25199
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -25199
transform -1 0 11316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_31
timestamp -25199
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -25199
transform -1 0 11316 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_32
timestamp -25199
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -25199
transform -1 0 11316 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_33
timestamp -25199
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -25199
transform -1 0 11316 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_34
timestamp -25199
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -25199
transform -1 0 11316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_35
timestamp -25199
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -25199
transform -1 0 11316 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -25199
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -25199
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_38
timestamp -25199
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp -25199
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_40
timestamp -25199
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_41
timestamp -25199
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_42
timestamp -25199
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_43
timestamp -25199
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_44
timestamp -25199
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_45
timestamp -25199
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_46
timestamp -25199
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_47
timestamp -25199
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_48
timestamp -25199
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_49
timestamp -25199
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_50
timestamp -25199
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_51
timestamp -25199
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_52
timestamp -25199
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_53
timestamp -25199
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_54
timestamp -25199
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_55
timestamp -25199
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_56
timestamp -25199
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_57
timestamp -25199
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_58
timestamp -25199
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_59
timestamp -25199
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_60
timestamp -25199
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_61
timestamp -25199
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_62
timestamp -25199
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_63
timestamp -25199
transform 1 0 3680 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_64
timestamp -25199
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_65
timestamp -25199
transform 1 0 8832 0 -1 11968
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 11702 2184 12502 2304 0 FreeSans 480 0 0 0 data_serial_o[0]
port 1 nsew signal output
flabel metal3 s 11702 7080 12502 7200 0 FreeSans 480 0 0 0 data_serial_o[1]
port 2 nsew signal output
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 fifo_data_i[0]
port 3 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 fifo_data_i[10]
port 4 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 fifo_data_i[11]
port 5 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 fifo_data_i[12]
port 6 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 fifo_data_i[13]
port 7 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 fifo_data_i[14]
port 8 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 fifo_data_i[15]
port 9 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 fifo_data_i[1]
port 10 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 fifo_data_i[2]
port 11 nsew signal input
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 fifo_data_i[3]
port 12 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 fifo_data_i[4]
port 13 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 fifo_data_i[5]
port 14 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 fifo_data_i[6]
port 15 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 fifo_data_i[7]
port 16 nsew signal input
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 fifo_data_i[8]
port 17 nsew signal input
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 fifo_data_i[9]
port 18 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 fifo_empty_i
port 19 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 fifo_rd_en_o
port 20 nsew signal output
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 rst_n
port 21 nsew signal input
flabel metal3 s 11702 11976 12502 12096 0 FreeSans 480 0 0 0 valid_serial_o
port 22 nsew signal output
flabel metal4 s 4208 2128 4528 12016 0 FreeSans 1920 90 0 0 vccd1
port 23 nsew power bidirectional
flabel metal4 s 4868 2128 5188 12016 0 FreeSans 1920 90 0 0 vssd1
port 24 nsew ground bidirectional
rlabel metal1 6210 11424 6210 11424 0 vccd1
rlabel metal1 6210 11968 6210 11968 0 vssd1
rlabel metal2 2898 3230 2898 3230 0 _000_
rlabel metal1 1748 2346 1748 2346 0 _001_
rlabel metal2 4738 3230 4738 3230 0 _002_
rlabel metal1 1932 4250 1932 4250 0 _003_
rlabel metal1 4968 4250 4968 4250 0 _004_
rlabel metal1 2530 5882 2530 5882 0 _005_
rlabel metal1 4922 5882 4922 5882 0 _006_
rlabel metal1 1978 6970 1978 6970 0 _007_
rlabel metal1 4554 7514 4554 7514 0 _008_
rlabel metal1 2208 8602 2208 8602 0 _009_
rlabel metal1 6808 8058 6808 8058 0 _010_
rlabel metal1 3726 10234 3726 10234 0 _011_
rlabel metal2 7314 10404 7314 10404 0 _012_
rlabel metal1 5244 10778 5244 10778 0 _013_
rlabel metal1 3956 9622 3956 9622 0 _014_
rlabel metal1 7406 9690 7406 9690 0 _015_
rlabel metal2 5290 10404 5290 10404 0 _016_
rlabel metal2 5382 9248 5382 9248 0 _017_
rlabel metal1 8142 4658 8142 4658 0 _018_
rlabel metal2 2070 6970 2070 6970 0 _019_
rlabel metal2 2530 10982 2530 10982 0 _020_
rlabel metal2 6670 10914 6670 10914 0 _021_
rlabel metal1 8234 5814 8234 5814 0 _022_
rlabel metal2 8050 6086 8050 6086 0 _023_
rlabel metal1 7498 5236 7498 5236 0 _024_
rlabel metal2 4094 9996 4094 9996 0 _025_
rlabel metal2 7774 5746 7774 5746 0 _026_
rlabel metal1 8372 5338 8372 5338 0 _027_
rlabel metal2 5290 3740 5290 3740 0 _028_
rlabel metal1 2806 4114 2806 4114 0 _029_
rlabel metal1 5980 4250 5980 4250 0 _030_
rlabel metal1 3174 5338 3174 5338 0 _031_
rlabel metal1 5658 5542 5658 5542 0 _032_
rlabel metal2 2990 6936 2990 6936 0 _033_
rlabel metal1 5382 7378 5382 7378 0 _034_
rlabel metal2 2898 8228 2898 8228 0 _035_
rlabel metal2 6394 8092 6394 8092 0 _036_
rlabel metal1 3128 11050 3128 11050 0 _037_
rlabel metal1 8280 8330 8280 8330 0 _038_
rlabel metal2 7038 4318 7038 4318 0 _039_
rlabel metal1 7176 6426 7176 6426 0 _040_
rlabel metal1 9246 5576 9246 5576 0 _041_
rlabel metal2 9522 5678 9522 5678 0 _042_
rlabel metal1 9476 3094 9476 3094 0 _043_
rlabel metal1 8832 7446 8832 7446 0 _044_
rlabel metal1 9568 10778 9568 10778 0 _045_
rlabel metal3 2660 1972 2660 1972 0 clk
rlabel metal1 5796 6630 5796 6630 0 clknet_0_clk
rlabel metal1 2530 2958 2530 2958 0 clknet_1_0__leaf_clk
rlabel metal1 9016 11118 9016 11118 0 clknet_1_1__leaf_clk
rlabel metal2 8602 4420 8602 4420 0 count\[0\]
rlabel metal1 8004 6290 8004 6290 0 count\[1\]
rlabel metal1 8970 5338 8970 5338 0 count\[2\]
rlabel metal1 10166 6358 10166 6358 0 count\[3\]
rlabel metal2 10718 2295 10718 2295 0 data_serial_o[0]
rlabel metal2 10810 6987 10810 6987 0 data_serial_o[1]
rlabel metal1 1426 3094 1426 3094 0 fifo_data_i[0]
rlabel metal1 1380 8534 1380 8534 0 fifo_data_i[10]
rlabel metal1 1380 9554 1380 9554 0 fifo_data_i[11]
rlabel metal1 1334 10030 1334 10030 0 fifo_data_i[12]
rlabel metal1 1380 10642 1380 10642 0 fifo_data_i[13]
rlabel metal1 1702 10064 1702 10064 0 fifo_data_i[14]
rlabel metal1 2714 11764 2714 11764 0 fifo_data_i[15]
rlabel metal1 1702 4080 1702 4080 0 fifo_data_i[1]
rlabel metal1 1334 4114 1334 4114 0 fifo_data_i[2]
rlabel metal1 1334 5202 1334 5202 0 fifo_data_i[3]
rlabel metal1 1380 5678 1380 5678 0 fifo_data_i[4]
rlabel metal1 1334 6290 1334 6290 0 fifo_data_i[5]
rlabel metal1 1702 6732 1702 6732 0 fifo_data_i[6]
rlabel metal1 1334 6766 1334 6766 0 fifo_data_i[7]
rlabel metal1 1380 7854 1380 7854 0 fifo_data_i[8]
rlabel metal1 1380 8466 1380 8466 0 fifo_data_i[9]
rlabel metal2 1242 11713 1242 11713 0 fifo_empty_i
rlabel metal1 1472 11798 1472 11798 0 fifo_rd_en_o
rlabel metal1 2530 3570 2530 3570 0 net1
rlabel metal2 1610 4590 1610 4590 0 net10
rlabel viali 6867 5270 6867 5270 0 net11
rlabel metal2 2806 5848 2806 5848 0 net12
rlabel metal2 1886 6120 1886 6120 0 net13
rlabel metal1 2116 6834 2116 6834 0 net14
rlabel metal2 1610 7616 1610 7616 0 net15
rlabel via1 3003 7786 3003 7786 0 net16
rlabel metal2 3266 11169 3266 11169 0 net17
rlabel metal2 3266 3298 3266 3298 0 net18
rlabel metal2 10994 2618 10994 2618 0 net19
rlabel metal2 3358 8636 3358 8636 0 net2
rlabel metal2 10994 6970 10994 6970 0 net20
rlabel metal2 1886 10812 1886 10812 0 net21
rlabel metal2 10994 11526 10994 11526 0 net22
rlabel metal1 3450 7310 3450 7310 0 net23
rlabel metal1 5658 8466 5658 8466 0 net24
rlabel metal1 8004 4998 8004 4998 0 net25
rlabel metal1 8096 10574 8096 10574 0 net26
rlabel metal2 3542 7276 3542 7276 0 net27
rlabel metal2 6118 5066 6118 5066 0 net28
rlabel metal1 3082 9622 3082 9622 0 net29
rlabel metal1 1610 9486 1610 9486 0 net3
rlabel metal2 8326 9010 8326 9010 0 net30
rlabel metal1 8740 8466 8740 8466 0 net31
rlabel metal1 2714 3570 2714 3570 0 net32
rlabel metal1 9384 10642 9384 10642 0 net33
rlabel metal1 2714 6800 2714 6800 0 net34
rlabel metal1 2254 11730 2254 11730 0 net35
rlabel metal1 4002 4046 4002 4046 0 net36
rlabel via1 5658 8398 5658 8398 0 net37
rlabel metal1 3227 2346 3227 2346 0 net38
rlabel metal1 3549 8874 3549 8874 0 net39
rlabel metal2 1610 9792 1610 9792 0 net4
rlabel metal2 7682 7616 7682 7616 0 net40
rlabel metal1 9614 8942 9614 8942 0 net41
rlabel metal1 6026 11227 6026 11227 0 net42
rlabel metal2 1886 10234 1886 10234 0 net5
rlabel metal1 5566 10064 5566 10064 0 net6
rlabel via1 5737 9622 5737 9622 0 net7
rlabel metal1 2438 3536 2438 3536 0 net8
rlabel metal1 3450 4046 3450 4046 0 net9
rlabel metal1 1380 3026 1380 3026 0 rst_n
rlabel metal1 5612 7718 5612 7718 0 shift_reg\[10\]
rlabel metal2 3450 8704 3450 8704 0 shift_reg\[11\]
rlabel metal1 6532 7854 6532 7854 0 shift_reg\[12\]
rlabel metal2 4922 10234 4922 10234 0 shift_reg\[13\]
rlabel metal2 8418 10234 8418 10234 0 shift_reg\[14\]
rlabel metal1 5980 10778 5980 10778 0 shift_reg\[15\]
rlabel metal1 4600 3162 4600 3162 0 shift_reg\[2\]
rlabel metal1 3266 2618 3266 2618 0 shift_reg\[3\]
rlabel metal1 6256 3162 6256 3162 0 shift_reg\[4\]
rlabel metal1 3036 4794 3036 4794 0 shift_reg\[5\]
rlabel metal2 6210 4590 6210 4590 0 shift_reg\[6\]
rlabel metal1 3450 6086 3450 6086 0 shift_reg\[7\]
rlabel metal1 6072 6086 6072 6086 0 shift_reg\[8\]
rlabel metal1 3128 7174 3128 7174 0 shift_reg\[9\]
rlabel metal1 2116 10642 2116 10642 0 state\[1\]
rlabel metal2 10718 11917 10718 11917 0 valid_serial_o
<< properties >>
string FIXED_BBOX 0 0 12502 14646
<< end >>
